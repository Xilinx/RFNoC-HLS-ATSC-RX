shortreal in[16384] =
'{0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1.55128708908113e-20,
2.71657093985046e-18,
1.05870672892733e-17,
3.24532699719380e-17,
7.61605836405662e-17,
1.60771591479415e-16,
3.01779151442308e-16,
5.17871179390951e-16,
8.17885061231622e-16,
1.18562293297442e-15,
1.58563201885378e-15,
1.89793888985795e-15,
1.97049742618565e-15,
1.46331495555610e-15,
-9.11947434749502e-18,
-3.18499126540899e-15,
-8.87777264896306e-15,
-1.82260687119941e-14,
-3.23757405433500e-14,
-5.28958489151837e-14,
-8.12892979383355e-14,
-1.19557982221005e-13,
-1.69257091523801e-13,
-2.32477502960099e-13,
-3.11355487832982e-13,
-4.08807102753039e-13,
-5.27515531256739e-13,
-6.70210740204291e-13,
-8.39825171211617e-13,
-1.03759557369687e-12,
-1.26547654733661e-12,
-1.52133904432472e-12,
-1.80394349631741e-12,
-2.10851626956943e-12,
-2.43075980350949e-12,
-2.76105570698459e-12,
-3.08908649528095e-12,
-3.39701379005464e-12,
-3.66376200211516e-12,
-3.85296265378865e-12,
-3.92384562342141e-12,
-3.94662861419315e-12,
-3.97893913997582e-12,
-3.98548164956547e-12,
-3.90327874189023e-12,
-3.67370413603685e-12,
-3.30098925624411e-12,
-2.84357823746029e-12,
-2.54764091767168e-12,
-2.79160527159872e-12,
-3.91323952408929e-12,
-6.26440435982922e-12,
-1.02095224635557e-11,
-1.60789472014589e-11,
-2.41682958368461e-11,
-3.45954445646335e-11,
-4.74964373387010e-11,
-6.32347160745006e-11,
-8.20315620986278e-11,
-1.04066463779695e-10,
-1.29554561523193e-10,
-1.58734109190206e-10,
-1.91875959565380e-10,
-2.29215174618602e-10,
-2.71115574435044e-10,
-3.17858961373929e-10,
-3.69827807267242e-10,
-4.27465174368535e-10,
-4.91043483652476e-10,
-5.60795576642903e-10,
-6.36930674868808e-10,
-7.19619475120226e-10,
-8.08861200241040e-10,
-9.04818331370905e-10,
-1.00777952649622e-09,
-1.11793241330815e-09,
-1.23562227116736e-09,
-1.36132038974779e-09,
-1.49543188943113e-09,
-1.63818247855829e-09,
-1.78978776244065e-09,
-1.95041494066572e-09,
-2.12019379830508e-09,
-2.29939911555732e-09,
-2.48816500736382e-09,
-2.68653255197648e-09,
-2.89457613433797e-09,
-3.11225867299925e-09,
-3.33954153219906e-09,
-3.57646801063538e-09,
-3.82300946455416e-09,
-4.07915345945753e-09,
-4.34507940738627e-09,
-4.62105642640154e-09,
-4.90751439485848e-09,
-5.20507414947247e-09,
-5.51456791342275e-09,
-5.83696069256234e-09,
-6.17313622441884e-09,
-6.52393428168807e-09,
-6.89022972011344e-09,
-7.27296622926588e-09,
-7.67315722072226e-09,
-8.09206213148173e-09,
-8.53090842412030e-09,
-8.99095731199395e-09,
-9.47367784220887e-09,
-9.98034010990523e-09,
-1.05122666127500e-08,
-1.10708926470693e-08,
-1.16577734132761e-08,
-1.22745227315590e-08,
-1.29226966905094e-08,
-1.36040396725434e-08,
-1.43202489866212e-08,
-1.50728602932304e-08,
-1.58633834956845e-08,
-1.66933507017575e-08,
-1.75644974120814e-08,
-1.84785982071389e-08,
-1.94372820061517e-08,
-2.04423002969634e-08,
-2.14954667399070e-08,
-2.25984955193326e-08,
-2.37531097013743e-08,
-2.49611620262158e-08,
-2.62246100390939e-08,
-2.75453473363996e-08,
-2.89253918595023e-08,
-3.03667384571327e-08,
-3.18713091473910e-08,
-3.34412106894888e-08,
-3.50784610247956e-08,
-3.67852024396598e-08,
-3.85636766964126e-08,
-4.04159976596930e-08,
-4.23443218267039e-08,
-4.43506813496697e-08,
-4.64370941699599e-08,
-4.86058304716153e-08,
-5.08591675441039e-08,
-5.31994146513171e-08,
-5.56289734277016e-08,
-5.81501140572982e-08,
-6.07651813311350e-08,
-6.34766408325049e-08,
-6.62870576206842e-08,
-6.91991175472140e-08,
-7.22154709364986e-08,
-7.53388036400793e-08,
-7.85717872986425e-08,
-8.19171788180029e-08,
-8.53778843179498e-08,
-8.89566535988706e-08,
-9.26563785696999e-08,
-9.64800861424919e-08,
-1.00430732175028e-07,
-1.04511464371626e-07,
-1.08725330960624e-07,
-1.13075344643221e-07,
-1.17564574964035e-07,
-1.22195928042856e-07,
-1.26972267366909e-07,
-1.31896740640514e-07,
-1.36972516884271e-07,
-1.42202637221089e-07,
-1.47590426990973e-07,
-1.53139183112216e-07,
-1.58852344611660e-07,
-1.64733378937854e-07,
-1.70785710906785e-07,
-1.77012950075550e-07,
-1.83418890742360e-07,
-1.90007298783712e-07,
-1.96781925865253e-07,
-2.03746623128609e-07,
-2.10905071185152e-07,
-2.18260851170271e-07,
-2.25817586851917e-07,
-2.33579029895736e-07,
-2.41548974599937e-07,
-2.49731300527856e-07,
-2.58129858821121e-07,
-2.66748543253925e-07,
-2.75591276022169e-07,
-2.84661894056626e-07,
-2.93964291131488e-07,
-3.03502304177528e-07,
-3.13279713282100e-07,
-3.23300326954268e-07,
-3.33568038968224e-07,
-3.44086885206707e-07,
-3.54860929974166e-07,
-3.65894408105305e-07,
-3.77191554434830e-07,
-3.88756575375737e-07,
-4.00593961558116e-07,
-4.12708203612056e-07,
-4.25103706902519e-07,
-4.37784848372758e-07,
-4.50755976544315e-07,
-4.64021695734118e-07,
-4.77586638680805e-07,
-4.91455580231559e-07,
-5.05633408920403e-07,
-5.20125070124777e-07,
-5.34935225005029e-07,
-5.50068705251761e-07,
-5.65530342555576e-07,
-5.81324911763659e-07,
-5.97457358253450e-07,
-6.13932684245810e-07,
-6.30755891961599e-07,
-6.47931926778256e-07,
-6.65465790916642e-07,
-6.83362543441035e-07,
-7.01627300259133e-07,
-7.20265290965472e-07,
-7.39281858841423e-07,
-7.58682460855198e-07,
-7.78472553975007e-07,
-7.98657708855899e-07,
-8.19243439309503e-07,
-8.40235202304029e-07,
-8.61638852711621e-07,
-8.83460131717584e-07,
-9.05704837350640e-07,
-9.28378653952677e-07,
-9.51487436395837e-07,
-9.75036982708843e-07,
-9.99032977233583e-07,
-1.02348110431194e-06,
-1.04838716197264e-06,
-1.07375717561808e-06,
-1.09959705696383e-06,
-1.12591283141228e-06,
-1.15271018330532e-06,
-1.17999513804534e-06,
-1.20777360734792e-06,
-1.23605161661544e-06,
-1.26483519125031e-06,
-1.29413047034177e-06,
-1.32394382035272e-06,
-1.35428115299874e-06,
-1.38514872105588e-06,
-1.41655266361340e-06,
-1.44849923344736e-06,
-1.48099491070752e-06,
-1.51404594816995e-06,
-1.54765882598440e-06,
-1.58183991061378e-06,
-1.61659568220784e-06,
-1.65193239354267e-06,
-1.68785641108116e-06,
-1.72437432865991e-06,
-1.76149274011550e-06,
-1.79921812559769e-06,
-1.83755696525623e-06,
-1.87651596661453e-06,
-1.91610183719604e-06,
-1.95632128452417e-06,
-1.99718101612234e-06,
-2.03868739845348e-06,
-2.08084748010151e-06,
-2.12366740015568e-06,
-2.16715397982625e-06,
-2.21131358557614e-06,
-2.25615303861559e-06,
-2.30167893278122e-06,
-2.34789808928326e-06,
-2.39481755670568e-06,
-2.44244415625872e-06,
-2.49078470915265e-06,
-2.53984626397141e-06,
-2.58963609667262e-06,
-2.64016125584021e-06,
-2.69142879005813e-06,
-2.74344574791030e-06,
-2.79621963272803e-06,
-2.84975726572156e-06,
-2.90406615022221e-06,
-2.95915333481389e-06,
-3.01502609545423e-06,
-3.07169193547452e-06,
-3.12915767608502e-06,
-3.18743059324333e-06,
-3.24651773553342e-06,
-3.30642569679185e-06,
-3.36716175297624e-06,
-3.42873272529687e-06,
-3.49114566233766e-06,
-3.55440738530888e-06,
-3.61852471542079e-06,
-3.68350447388366e-06,
-3.74935348190775e-06,
-3.81607878807699e-06,
-3.88368744097534e-06,
-3.95218694393407e-06,
-4.02158366341610e-06,
-4.09188533012639e-06,
-4.16309876527521e-06,
-4.23523124482017e-06,
-4.30829004471889e-06,
-4.38228244092898e-06,
-4.45721570940805e-06,
-4.53309758086107e-06,
-4.60993487649830e-06,
-4.68773441753001e-06,
-4.76650393466116e-06,
-4.84625070384936e-06,
-4.92698200105224e-06,
-5.00870510222740e-06,
-5.09142819282715e-06,
-5.17515854880912e-06,
-5.25990390087827e-06,
-5.34567197973956e-06,
-5.43247006135061e-06,
-5.52030633116374e-06,
-5.60918851988390e-06,
-5.69912435821607e-06,
-5.79012248635991e-06,
-5.88219063502038e-06,
-5.97533698964980e-06,
-6.06956973570050e-06,
-6.16489751337213e-06,
-6.26132850811700e-06,
-6.35887136013480e-06,
-6.45753425487783e-06,
-6.55732537779841e-06,
-6.65825336909620e-06,
-6.76032595947618e-06,
-6.86355178913800e-06,
-6.96793904353399e-06,
-7.07349636286381e-06,
-7.18023147783242e-06,
-7.28815302863950e-06,
-7.39726965548471e-06,
-7.50758908907301e-06,
-7.61911996960407e-06,
-7.73187093727756e-06,
-7.84584972279845e-06,
-7.96106542111374e-06,
-8.07752712717047e-06,
-8.19524302642094e-06,
-8.31422221381217e-06,
-8.43447378429119e-06,
-8.55600592331030e-06,
-8.67882772581652e-06,
-8.80294737726217e-06,
-8.92837488208897e-06,
-9.05511842574924e-06,
-9.18318710318999e-06,
-9.31259000935825e-06,
-9.44333532970632e-06,
-9.57543215918122e-06,
-9.70888959272998e-06,
-9.84371581580490e-06,
-9.97991992335301e-06,
-1.01175101008266e-05,
-1.02564954431728e-05,
-1.03968841358437e-05,
-1.05386843642918e-05,
-1.06819052234641e-05,
-1.08265558083076e-05,
-1.09726443042746e-05,
-1.11201798063121e-05,
-1.12691714093671e-05,
-1.14196272988920e-05,
-1.15715574793285e-05,
-1.17249701361288e-05,
-1.18798734547454e-05,
-1.20362774396199e-05,
-1.21941911856993e-05,
-1.23536237879307e-05,
-1.25145843412611e-05,
-1.26770810311427e-05,
-1.28411238620174e-05,
-1.30067219288321e-05,
-1.31738843265339e-05,
-1.33426210595644e-05,
-1.35129412228707e-05,
-1.36848539113998e-05,
-1.38583682200988e-05,
-1.40334941534093e-05,
-1.42102408062783e-05,
-1.43886181831476e-05,
-1.45686344694695e-05,
-1.47502996696858e-05,
-1.49336228787433e-05,
-1.51186131915892e-05,
-1.53052806126652e-05,
-1.54936333274236e-05,
-1.56836813403061e-05,
-1.58754337462597e-05,
-1.60688996402314e-05,
-1.62640899361577e-05,
-1.64610119099962e-05,
-1.66596764756832e-05,
-1.68600909091765e-05,
-1.70622661244124e-05,
-1.72662112163380e-05,
-1.74719352799002e-05,
-1.76794474100461e-05,
-1.78887585207121e-05,
-1.80998777068453e-05,
-1.83128140633926e-05,
-1.85275785042904e-05,
-1.87441801244859e-05,
-1.89626298379153e-05,
-1.91829367395258e-05,
-1.94051117432537e-05,
-1.96291639440460e-05,
-1.98551042558393e-05,
-2.00829417735804e-05,
-2.03126874112058e-05,
-2.05443484446732e-05,
-2.07779376069084e-05,
-2.10134621738689e-05,
-2.12509330594912e-05,
-2.14903593587223e-05,
-2.17317501665093e-05,
-2.19751163967885e-05,
-2.22204671445070e-05,
-2.24678115046117e-05,
-2.27171603910392e-05,
-2.29685228987364e-05,
-2.32219099416398e-05,
-2.34773324336857e-05,
-2.37347976508318e-05,
-2.39943183260039e-05,
-2.42559035541490e-05,
-2.45195660681929e-05,
-2.47853149630828e-05,
-2.50531593337655e-05,
-2.53231119131669e-05,
-2.55951817962341e-05,
-2.58693798969034e-05,
-2.61457171291113e-05,
-2.64242025878048e-05,
-2.67048471869202e-05,
-2.69876618403941e-05,
-2.72726574621629e-05,
-2.75598449661629e-05,
-2.78492352663307e-05,
-2.81408392766025e-05,
-2.84346660919255e-05,
-2.87307266262360e-05,
-2.90290336124599e-05,
-2.93295961455442e-05,
-2.96324269584147e-05,
-2.99375351460185e-05,
-3.02449316222919e-05,
-3.05546273011714e-05,
-3.08666349155828e-05,
-3.11809635604732e-05,
-3.14976241497789e-05,
-3.18166275974363e-05,
-3.21379848173820e-05,
-3.24617067235522e-05,
-3.27878078678623e-05,
-3.31162955262698e-05,
-3.34471842506900e-05,
-3.37804813170806e-05,
-3.41162012773566e-05,
-3.44543514074758e-05,
-3.47949462593533e-05,
-3.51379967469256e-05,
-3.54835137841292e-05,
-3.58315082849003e-05,
-3.61819948011544e-05,
-3.65349806088489e-05,
-3.68904766219202e-05,
-3.72484973922838e-05,
-3.76090538338758e-05,
-3.79721568606328e-05,
-3.83378173864912e-05,
-3.87060499633662e-05,
-3.90768618672155e-05,
-3.94502676499542e-05,
-3.98262782255188e-05,
-4.02049045078456e-05,
-4.05861574108712e-05,
-4.09700478485320e-05,
-4.13565903727431e-05,
-4.17457922594622e-05,
-4.21376680606045e-05,
-4.25322286901064e-05,
-4.29294850619044e-05,
-4.33294517279137e-05,
-4.37321359640919e-05,
-4.41375523223542e-05,
-4.45457080786582e-05,
-4.49566177849192e-05,
-4.53702923550736e-05,
-4.57867427030578e-05,
-4.62059833807871e-05,
-4.66280216642190e-05,
-4.70528721052688e-05,
-4.74805456178729e-05,
-4.79110567539465e-05,
-4.83444127894472e-05,
-4.87806282762904e-05,
-4.92197141284123e-05,
-4.96616848977283e-05,
-5.01065514981747e-05,
-5.05543248436879e-05,
-5.10050158482045e-05,
-5.14586390636396e-05,
-5.19152017659508e-05,
-5.23747185070533e-05,
-5.28372038388625e-05,
-5.33026650373358e-05,
-5.37711166543886e-05,
-5.42425696039572e-05,
-5.47170384379569e-05,
-5.51945340703242e-05,
-5.56750674149953e-05,
-5.61586493859068e-05,
-5.66452945349738e-05,
-5.71350137761328e-05,
-5.76278180233203e-05,
-5.81237181904726e-05,
-5.86227288295049e-05,
-5.91248644923326e-05,
-5.96301360928919e-05,
-6.01385545451194e-05,
-6.06501307629515e-05,
-6.11648792983033e-05,
-6.16828110651113e-05,
-6.22039442532696e-05,
-6.27282861387357e-05,
-6.32558512734249e-05,
-6.37866469332948e-05,
-6.43206949462183e-05,
-6.48580025881529e-05,
-6.53985844110139e-05,
-6.59424476907589e-05,
-6.64896069793031e-05,
-6.70400768285617e-05,
-6.75938717904501e-05,
-6.81509991409257e-05,
-6.87114734319039e-05,
-6.92753092152998e-05,
-6.98425210430287e-05,
-7.04131161910482e-05,
-7.09871092112735e-05,
-7.15645073796623e-05,
-7.21453325240873e-05,
-7.27295919205062e-05,
-7.33173001208343e-05,
-7.39084716769867e-05,
-7.45031211408787e-05,
-7.51012557884678e-05,
-7.57028901716694e-05,
-7.63080388423987e-05,
-7.69167163525708e-05,
-7.75289372541010e-05,
-7.81447160989046e-05,
-7.87640601629391e-05,
-7.93869839981198e-05,
-8.00135021563619e-05,
-8.06436219136231e-05,
-8.12773650977761e-05,
-8.19147389847785e-05,
-8.25557508505881e-05,
-8.32004225230776e-05,
-8.38487612782046e-05,
-8.45007889438421e-05,
-8.51565127959475e-05,
-8.58159401104786e-05,
-8.64790927153081e-05,
-8.71459778863937e-05,
-8.78166174516082e-05,
-8.84910186869092e-05,
-8.91691961442120e-05,
-8.98511643754318e-05,
-9.05369379324839e-05,
-9.12265240913257e-05,
-9.19199446798302e-05,
-9.26172142499127e-05,
-9.33183400775306e-05,
-9.40233367145993e-05,
-9.47322259889916e-05,
-9.54450151766650e-05,
-9.61617188295350e-05,
-9.68823514995165e-05,
-9.76069277385250e-05,
-9.83354620984756e-05,
-9.90679691312835e-05,
-9.98044561129063e-05,
-0.000100544944871217,
-0.000101289442682173,
-0.000102037971373647,
-0.000102790538221598,
-0.000103547157777939,
-0.000104307844594587,
-0.000105072613223456,
-0.000105841478216462,
-0.000106614446849562,
-0.000107391540950630,
-0.000108172775071580,
-0.000108958156488370,
-0.000109747707028873,
-0.000110541433969047,
-0.000111339351860806,
-0.000112141482532024,
-0.000112947833258659,
-0.000113758418592624,
-0.000114573253085837,
-0.000115392351290211,
-0.000116215727757663,
-0.000117043404316064,
-0.000117875388241373,
-0.000118711694085505,
-0.000119552336400375,
-0.000120397329737898,
-0.000121246688649990,
-0.000122100420412608,
-0.000122958546853624,
-0.000123821082524955,
-0.000124688056530431,
-0.000125559468870051,
-0.000126435334095731,
-0.000127315666759387,
-0.000128200481412932,
-0.000129089792608283,
-0.000129983629449271,
-0.000130881991935894,
-0.000131784894620068,
-0.000132692366605625,
-0.000133604407892562,
-0.000134521047584713,
-0.000135442285682075,
-0.000136368151288480,
-0.000137298658955842,
-0.000138233808684163,
-0.000139173629577272,
-0.000140118136187084,
-0.000141067343065515,
-0.000142021264764480,
-0.000142979915835895,
-0.000143943310831673,
-0.000144911464303732,
-0.000145884390803985,
-0.000146862104884349,
-0.000147844635648653,
-0.000148831983096898,
-0.000149824176332913,
-0.000150821215356700,
-0.000151823129272088,
-0.000152829918079078,
-0.000153841610881500,
-0.000154858222231269,
-0.000155879766680300,
-0.000156906258780509,
-0.000157937713083811,
-0.000158974144142121,
-0.000160015566507354,
-0.000161062009283341,
-0.000162113472470082,
-0.000163169985171407,
-0.000164231547387317,
-0.000165298188221641,
-0.000166369907674380,
-0.000167446734849364,
-0.000168528684298508,
-0.000169615770573728,
-0.000170708008226939,
-0.000171805411810055,
-0.000172907995874994,
-0.000174015774973668,
-0.000175128763657995,
-0.000176246991031803,
-0.000177370457095094,
-0.000178499176399782,
-0.000179633178049698,
-0.000180772462044843,
-0.000181917057489045,
-0.000183066978934221,
-0.000184222240932286,
-0.000185382858035155,
-0.000186548830242828,
-0.000187720201211050,
-0.000188896970939823,
-0.000190079153981060,
-0.000191266764886677,
-0.000192459832760505,
-0.000193658357602544,
-0.000194862368516624,
-0.000196071880054660,
-0.000197286892216653,
-0.000198507434106432,
-0.000199733520275913,
-0.000200965165277012,
-0.000202202398213558,
-0.000203445219085552,
-0.000204693656996824,
-0.000205947711947374,
-0.000207207413041033,
-0.000208472774829716,
-0.000209743811865337,
-0.000211020538699813,
-0.000212302969885059,
-0.000213591119972989,
-0.000214885018067434,
-0.000216184678720310,
-0.000217490101931617,
-0.000218801316805184,
-0.000220118337892927,
-0.000221441194298677,
-0.000222769886022434,
-0.000224104427616112,
-0.000225444848183543,
-0.000226791162276641,
-0.000228143384447321,
-0.000229501529247500,
-0.000230865611229092,
-0.000232235659495927,
-0.000233611674048007,
-0.000234993683989160,
-0.000236381703871302,
-0.000237775748246349,
-0.000239175831666216,
-0.000240581983234733,
-0.000241994202951901,
-0.000243412519921549,
-0.000244836963247508,
-0.000246267532929778,
-0.000247704243520275,
-0.000249147124122828,
-0.000250596174737439,
-0.000252051424467936,
-0.000253512902418152,
-0.000254980608588085,
-0.000256454572081566,
-0.000257934792898595,
-0.000259421300143003,
-0.000260914122918621,
-0.000262413261225447,
-0.000263918744167313,
-0.000265430571744218,
-0.000266948773059994,
-0.000268473348114640,
-0.000270004326011986,
-0.000271541735855863,
-0.000273085577646270,
-0.000274635851383209,
-0.000276192615274340,
-0.000277755869319662,
-0.000279325613519177,
-0.000280901876976714,
-0.000282484688796103,
-0.000284074048977345,
-0.000285669986624271,
-0.000287272501736879,
-0.000288881623419002,
-0.000290497380774468,
-0.000292119773803279,
-0.000293748831609264,
-0.000295384554192424,
-0.000297026970656589,
-0.000298676081001759,
-0.000300331943435594,
-0.000301994528854266,
-0.000303663895465434,
-0.000305340043269098,
-0.000307022972265258,
-0.000308712740661576,
-0.000310409348458052,
-0.000312112795654684,
-0.000313823111355305,
-0.000315540324663743,
-0.000317264435580000,
-0.000318995473207906,
-0.000320733466651291,
-0.000322478415910155,
-0.000324230350088328,
-0.000325989269185811,
-0.000327755202306435,
-0.000329528178554028,
-0.000331308197928593,
-0.000333095289533958,
-0.000334889482473955,
-0.000336690776748583,
-0.000338499201461673,
-0.000340314756613225,
-0.000342137471307069,
-0.000343967374647036,
-0.000345804495736957,
-0.000347648805473000,
-0.000349500362062827,
-0.000351359165506437,
-0.000353225244907662,
-0.000355098629370332,
-0.000356979318894446,
-0.000358867342583835,
-0.000360762729542330,
-0.000362665479769930,
-0.000364575622370467,
-0.000366493157343939,
-0.000368418113794178,
-0.000370350520825014,
-0.000372290407540277,
-0.000374237773939967,
-0.000376192649127916,
-0.000378155033104122,
-0.000380124984076247,
-0.000382102502044290,
-0.000384087587008253,
-0.000386080268071964,
-0.000388080574339256,
-0.000390088534913957,
-0.000392104149796069,
-0.000394127448089421,
-0.000396158429794014,
-0.000398197153117508,
-0.000400243588956073,
-0.000402297795517370,
-0.000404359772801399,
-0.000406429549911991,
-0.000408507155952975,
-0.000410592590924352,
-0.000412685883929953,
-0.000414787064073607,
-0.000416896131355315,
-0.000419013114878908,
-0.000421138043748215,
-0.000423270947067067,
-0.000425411824835464,
-0.000427560706157237,
-0.000429717620136216,
-0.000431882566772401,
-0.000434055575169623,
-0.000436236674431711,
-0.000438425893662497,
-0.000440623232861981,
-0.000442828721133992,
-0.000445042387582362,
-0.000447264232207090,
-0.000449494284112006,
-0.000451732572400942,
-0.000453979126177728,
-0.000456233945442364,
-0.000458497059298679,
-0.000460768496850505,
-0.000463048287201673,
-0.000465336430352181,
-0.000467632955405861,
-0.000469937891466543,
-0.000472251238534227,
-0.000474573025712743,
-0.000476903282105923,
-0.000479242036817595,
-0.000481589289847761,
-0.000483945099404082,
-0.000486309465486556,
-0.000488682417199016,
-0.000491063925437629,
-0.000493454048410058,
-0.000495852844323963,
-0.000498260313179344,
-0.000500676454976201,
-0.000503101327922195,
-0.000505534932017326,
-0.000507977267261595,
-0.000510428391862661,
-0.000512888305820525,
-0.000515357067342848,
-0.000517834618221968,
-0.000520321074873209,
-0.000522816379088908,
-0.000525320589076728,
-0.000527833763044328,
-0.000530355900991708,
-0.000532887002918869,
-0.000535427068825811,
-0.000537976156920195,
-0.000540534325409681,
-0.000543101516086608,
-0.000545677845366299,
-0.000548263255041093,
-0.000550857803318650,
-0.000553461490198970,
-0.000556074373889715,
-0.000558696454390883,
-0.000561327789910138,
-0.000563968380447477,
-0.000566618226002902,
-0.000569277384784073,
-0.000571945856790990,
-0.000574623642023653,
-0.000577310798689723,
-0.000580007326789200,
-0.000582713284529746,
-0.000585428671911359,
-0.000588153547141701,
-0.000590887910220772,
-0.000593631761148572,
-0.000596385158132762,
-0.000599148101173341,
-0.000601920648477972,
-0.000604702800046653,
-0.000607494555879384,
-0.000610295974183828,
-0.000613107054959983,
-0.000615927856415510,
-0.000618758378550410,
-0.000621598679572344,
-0.000624448759481311,
-0.000627308618277311,
-0.000630178314168006,
-0.000633057847153395,
-0.000635947275441140,
-0.000638846599031240,
-0.000641755817923695,
-0.000644674990326166,
-0.000647604116238654,
-0.000650543253868818,
-0.000653492403216660,
-0.000656451622489840,
-0.000659420911688358,
-0.000662400329019874,
-0.000665389816276729,
-0.000668389489874244,
-0.000671399349812418,
-0.000674419396091253,
-0.000677449628710747,
-0.000680490164086223,
-0.000683540944010019,
-0.000686602026689798,
-0.000689673470333219,
-0.000692755216732621,
-0.000695847382303327,
-0.000698949967045337,
-0.000702062970958650,
-0.000705186394043267,
-0.000708320294506848,
-0.000711464730557054,
-0.000714619702193886,
-0.000717785209417343,
-0.000720961310435087,
-0.000724148063454777,
-0.000727345468476415,
-0.000730553525500000,
-0.000733772234525532,
-0.000737001711968333,
-0.000740241899620742,
-0.000743492855690420,
-0.000746754638385028,
-0.000750027247704566,
-0.000753310683649033,
-0.000756605004426092,
-0.000759910268243402,
-0.000763226416893303,
-0.000766553566791117,
-0.000769891717936844,
-0.000773240870330483,
-0.000776601082179695,
-0.000779972353484482,
-0.000783354684244841,
-0.000786748132668436,
-0.000790152756962925,
-0.000793568557128310,
-0.000796995591372252,
-0.000800433801487088,
-0.000803883303888142,
-0.000807344098575413,
-0.000810816185548902,
-0.000814299623016268,
-0.000817794410977513,
-0.000821300607640296,
-0.000824818213004619,
-0.000828347285278142,
-0.000831887824460864,
-0.000835439888760448,
-0.000839003478176892,
-0.000842578650917858,
-0.000846165406983346,
-0.000849763746373355,
-0.000853373727295548,
-0.000856995407957584,
-0.000860628788359463,
-0.000864273926708847,
-0.000867930823005736,
-0.000871599477250129,
-0.000875279947649688,
-0.000878972292412072,
-0.000882676511537284,
-0.000886392605025321,
-0.000890120631083846,
-0.000893860647920519,
-0.000897612655535340,
-0.000901376653928310,
-0.000905152701307088,
-0.000908940855879337,
-0.000912741117645055,
-0.000916553486604244,
-0.000920378020964563,
-0.000924214778933674,
-0.000928063760511577,
-0.000931924965698272,
-0.000935798452701420,
-0.000939684221521020,
-0.000943582330364734,
-0.000947492837440223,
-0.000951415742747486,
-0.000955351046286523,
-0.000959298806264997,
-0.000963259080890566,
-0.000967231870163232,
-0.000971217174082995,
-0.000975215050857514,
-0.000979225500486791,
-0.000983248581178486,
-0.000987284351140261,
-0.000991332810372114,
-0.000995393958874047,
-0.000999467913061380,
-0.00100355455651879,
-0.00100765400566161,
-0.00101176637690514,
-0.00101589155383408,
-0.00102002965286374,
-0.00102418067399412,
-0.00102834461722523,
-0.00103252159897238,
-0.00103671161923558,
-0.00104091467801481,
-0.00104513077531010,
-0.00104936002753675,
-0.00105360243469477,
-0.00105785799678415,
-0.00106212683022022,
-0.00106640881858766,
-0.00107070407830179,
-0.00107501260936260,
-0.00107933452818543,
-0.00108366983477026,
-0.00108801852911711,
-0.00109238061122596,
-0.00109675608109683,
-0.00110114505514503,
-0.00110554753337055,
-0.00110996363218874,
-0.00111439323518425,
-0.00111883645877242,
-0.00112329330295324,
-0.00112776388414204,
-0.00113224808592349,
-0.00113674602471292,
-0.00114125781692564,
-0.00114578334614635,
-0.00115032272879034,
-0.00115487596485764,
-0.00115944305434823,
-0.00116402399726212,
-0.00116861891001463,
-0.00117322779260576,
-0.00117785076145083,
-0.00118248770013452,
-0.00118713872507215,
-0.00119180383626372,
-0.00119648315012455,
-0.00120117655023932,
-0.00120588415302336,
-0.00121060607489198,
-0.00121534219942987,
-0.00122009264305234,
-0.00122485740575939,
-0.00122963648755103,
-0.00123443000484258,
-0.00123923795763403,
-0.00124406034592539,
-0.00124889716971666,
-0.00125374854542315,
-0.00125861447304487,
-0.00126349495258182,
-0.00126839010044932,
-0.00127329980023205,
-0.00127822416834533,
-0.00128316332120448,
-0.00128811714239419,
-0.00129308574832976,
-0.00129806913901120,
-0.00130306731443852,
-0.00130808039102703,
-0.00131310836877674,
-0.00131815124768764,
-0.00132320914417505,
-0.00132828194182366,
-0.00133336975704879,
-0.00133847270626575,
-0.00134359067305923,
-0.00134872377384454,
-0.00135387200862169,
-0.00135903537739068,
-0.00136421399656683,
-0.00136940786615014,
-0.00137461698614061,
-0.00137984147295356,
-0.00138508121017367,
-0.00139033631421626,
-0.00139560690149665,
-0.00140089285559952,
-0.00140619429294020,
-0.00141151121351868,
-0.00141684361733496,
-0.00142219162080437,
-0.00142755522392690,
-0.00143293442670256,
-0.00143832934554666,
-0.00144373986404389,
-0.00144916609860957,
-0.00145460816565901,
-0.00146006594877690,
-0.00146553956437856,
-0.00147102901246399,
-0.00147653440944850,
-0.00148205563891679,
-0.00148759281728417,
-0.00149314594455063,
-0.00149871513713151,
-0.00150430039502680,
-0.00150990171823651,
-0.00151551910676062,
-0.00152115267701447,
-0.00152680242899805,
-0.00153246836271137,
-0.00153815047815442,
-0.00154384889174253,
-0.00154956360347569,
-0.00155529461335391,
-0.00156104203779250,
-0.00156680587679148,
-0.00157258613035083,
-0.00157838279847056,
-0.00158419599756598,
-0.00159002572763711,
-0.00159587198868394,
-0.00160173478070647,
-0.00160761422012001,
-0.00161351030692458,
-0.00161942304112017,
-0.00162535253912210,
-0.00163129880093038,
-0.00163726182654500,
-0.00164324161596596,
-0.00164923828560859,
-0.00165525183547288,
-0.00166128226555884,
-0.00166732969228178,
-0.00167339411564171,
-0.00167947553563863,
-0.00168557395227253,
-0.00169168948195875,
-0.00169782200828195,
-0.00170397176407278,
-0.00171013863291591,
-0.00171632273122668,
-0.00172252405900508,
-0.00172874261625111,
-0.00173497851938009,
-0.00174123165197670,
-0.00174750224687159,
-0.00175379018764943,
-0.00176009559072554,
-0.00176641845609993,
-0.00177275878377259,
-0.00177911657374352,
-0.00178549194242805,
-0.00179188488982618,
-0.00179829541593790,
-0.00180472363717854,
-0.00181116943713278,
-0.00181763304863125,
-0.00182411435525864,
-0.00183061347343028,
-0.00183713028673083,
-0.00184366502799094,
-0.00185021758079529,
-0.00185678806155920,
-0.00186337647028267,
-0.00186998280696571,
-0.00187660707160831,
-0.00188324938062578,
-0.00188990973401815,
-0.00189658813178539,
-0.00190328469034284,
-0.00190999940969050,
-0.00191673228982836,
-0.00192348333075643,
-0.00193025264889002,
-0.00193704024422914,
-0.00194384611677378,
-0.00195067038293928,
-0.00195751292631030,
-0.00196437397971749,
-0.00197125342674553,
-0.00197815126739442,
-0.00198506750166416,
-0.00199200236238539,
-0.00199895584955812,
-0.00200592773035169,
-0.00201291823759675,
-0.00201992760412395,
-0.00202695559710264,
-0.00203400221653283,
-0.00204106769524515,
-0.00204815180040896,
-0.00205525476485491,
-0.00206237658858299,
-0.00206951727159321,
-0.00207667681388557,
-0.00208385521546006,
-0.00209105270914733,
-0.00209826906211674,
-0.00210550450719893,
-0.00211275904439390,
-0.00212003267370164,
-0.00212732539512217,
-0.00213463720865548,
-0.00214196834713221,
-0.00214931857772172,
-0.00215668813325465,
-0.00216407701373100,
-0.00217148521915078,
-0.00217891274951398,
-0.00218635960482061,
-0.00219382578507066,
-0.00220131152309477,
-0.00220881658606231,
-0.00221634120680392,
-0.00222388538531959,
-0.00223144912160933,
-0.00223903241567314,
-0.00224663526751101,
-0.00225425790995359,
-0.00226190034300089,
-0.00226956233382225,
-0.00227724411524832,
-0.00228494568727911,
-0.00229266704991460,
-0.00230040843598545,
-0.00230816961266100,
-0.00231595081277192,
-0.00232375180348754,
-0.00233157281763852,
-0.00233941385522485,
-0.00234727491624653,
-0.00235515623353422,
-0.00236305757425725,
-0.00237097917124629,
-0.00237892079167068,
-0.00238688266836107,
-0.00239486480131745,
-0.00240286719053984,
-0.00241089006885886,
-0.00241893320344389,
-0.00242699682712555,
-0.00243508070707321,
-0.00244318507611752,
-0.00245130993425846,
-0.00245945528149605,
-0.00246762111783028,
-0.00247580767609179,
-0.00248401472344995,
-0.00249224249273539,
-0.00250049098394811,
-0.00250876019708812,
-0.00251705013215542,
-0.00252536078915000,
-0.00253369240090251,
-0.00254204473458231,
-0.00255041802302003,
-0.00255881226621568,
-0.00256722746416926,
-0.00257566361688077,
-0.00258412072435021,
-0.00259259901940823,
-0.00260109826922417,
-0.00260961870662868,
-0.00261816033162177,
-0.00262672314420342,
-0.00263530714437366,
-0.00264391256496310,
-0.00265253917314112,
-0.00266118720173836,
-0.00266985641792417,
-0.00267854705452919,
-0.00268725911155343,
-0.00269599282182753,
-0.00270474795252085,
-0.00271352450363338,
-0.00272232270799577,
-0.00273114256560802,
-0.00273998407647014,
-0.00274884724058211,
-0.00275773205794394,
-0.00276663852855563,
-0.00277556688524783,
-0.00278451712802053,
-0.00279348902404308,
-0.00280248280614615,
-0.00281149870716035,
-0.00282053649425507,
-0.00282959616743028,
-0.00283867795951664,
-0.00284778163768351,
-0.00285690743476152,
-0.00286605535075068,
-0.00287522538565099,
-0.00288441777229309,
-0.00289363227784634,
-0.00290286913514137,
-0.00291212811134756,
-0.00292140943929553,
-0.00293071311898530,
-0.00294003915041685,
-0.00294938776642084,
-0.00295875873416662,
-0.00296815228648484,
-0.00297756819054484,
-0.00298700667917728,
-0.00299646775238216,
-0.00300595164299011,
-0.00301545811817050,
-0.00302498717792332,
-0.00303453905507922,
-0.00304411374963820,
-0.00305371126160026,
-0.00306333159096539,
-0.00307297473773360,
-0.00308264070190489,
-0.00309232971630991,
-0.00310204154811800,
-0.00311177643015981,
-0.00312153436243534,
-0.00313131534494460,
-0.00314111961051822,
-0.00315094692632556,
-0.00316079752519727,
-0.00317067117430270,
-0.00318056810647249,
-0.00319048832170665,
-0.00320043182000518,
-0.00321039860136807,
-0.00322038889862597,
-0.00323040271177888,
-0.00324043980799615,
-0.00325050042010844,
-0.00326058454811573,
-0.00327069242484868,
-0.00328082381747663,
-0.00329097872599959,
-0.00330115738324821,
-0.00331135978922248,
-0.00332158594392240,
-0.00333183584734797,
-0.00334210949949920,
-0.00335240713320673,
-0.00336272851563990,
-0.00337307387962937,
-0.00338344322517514,
-0.00339383655227721,
-0.00340425386093557,
-0.00341469538398087,
-0.00342516088858247,
-0.00343565060757101,
-0.00344616454094648,
-0.00345670268870890,
-0.00346726505085826,
-0.00347785162739456,
-0.00348846265114844,
-0.00349909788928926,
-0.00350975757464767,
-0.00352044170722365,
-0.00353115028701723,
-0.00354188354685903,
-0.00355264125391841,
-0.00356342364102602,
-0.00357423047535121,
-0.00358506198972464,
-0.00359591818414629,
-0.00360679929144681,
-0.00361770507879555,
-0.00362863554619253,
-0.00363959092646837,
-0.00365057121962309,
-0.00366157642565668,
-0.00367260654456913,
-0.00368366180919111,
-0.00369474198669195,
-0.00370584730990231,
-0.00371697777882218,
-0.00372813316062093,
-0.00373931392095983,
-0.00375051982700825,
-0.00376175087876618,
-0.00377300730906427,
-0.00378428911790252,
-0.00379559630528092,
-0.00380692887119949,
-0.00381828681565821,
-0.00382967037148774,
-0.00384107930585742,
-0.00385251385159791,
-0.00386397400870919,
-0.00387545977719128,
-0.00388697115704417,
-0.00389850838109851,
-0.00391007121652365,
-0.00392165966331959,
-0.00393327418714762,
-0.00394491432234645,
-0.00395658053457737,
-0.00396827282384038,
-0.00397999072447419,
-0.00399173470214009,
-0.00400350475683808,
-0.00401530088856816,
-0.00402712309733033,
-0.00403897138312459,
-0.00405084621161223,
-0.00406274711713195,
-0.00407467456534505,
-0.00408662809059024,
-0.00409860815852881,
-0.00411061430349946,
-0.00412264699116349,
-0.00413470622152090,
-0.00414679199457169,
-0.00415890431031585,
-0.00417104316875339,
-0.00418320856988430,
-0.00419540097936988,
-0.00420761993154883,
-0.00421986542642117,
-0.00423213792964816,
-0.00424443697556853,
-0.00425676302984357,
-0.00426911609247327,
-0.00428149616345763,
-0.00429390324279666,
-0.00430633733049035,
-0.00431879842653871,
-0.00433128653094173,
-0.00434380164369941,
-0.00435634423047304,
-0.00436891382560134,
-0.00438151089474559,
-0.00439413543790579,
-0.00440678698942065,
-0.00441946601495147,
-0.00443217251449823,
-0.00444490648806095,
-0.00445766793563962,
-0.00447045685723424,
-0.00448327371850610,
-0.00449611805379391,
-0.00450898986309767,
-0.00452188961207867,
-0.00453481683507562,
-0.00454777199774981,
-0.00456075510010123,
-0.00457376614212990,
-0.00458680512383580,
-0.00459987204521894,
-0.00461296690627933,
-0.00462608970701695,
-0.00463924044743180,
-0.00465241959318519,
-0.00466562667861581,
-0.00467886216938496,
-0.00469212559983134,
-0.00470541743561626,
-0.00471873767673969,
-0.00473208632320166,
-0.00474546337500215,
-0.00475886883214116,
-0.00477230269461870,
-0.00478576496243477,
-0.00479925610125065,
-0.00481277564540505,
-0.00482632359489799,
-0.00483990041539073,
-0.00485350610688329,
-0.00486714020371437,
-0.00488080317154527,
-0.00489449501037598,
-0.00490821572020650,
-0.00492196530103684,
-0.00493574421852827,
-0.00494955200701952,
-0.00496338866651058,
-0.00497725466266274,
-0.00499114952981472,
-0.00500507373362780,
-0.00501902727410197,
-0.00503300968557596,
-0.00504702143371105,
-0.00506106251850724,
-0.00507513293996453,
-0.00508923316374421,
-0.00510336272418499,
-0.00511752162128687,
-0.00513171032071114,
-0.00514592835679650,
-0.00516017619520426,
-0.00517445337027311,
-0.00518876034766436,
-0.00520309712737799,
-0.00521746370941401,
-0.00523186009377241,
-0.00524628628045321,
-0.00526074273511767,
-0.00527522899210453,
-0.00528974505141377,
-0.00530429137870669,
-0.00531886750832200,
-0.00533347390592098,
-0.00534811057150364,
-0.00536277750506997,
-0.00537747470661998,
-0.00539220217615366,
-0.00540695991367102,
-0.00542174791917205,
-0.00543656619265676,
-0.00545141519978643,
-0.00546629447489977,
-0.00548120448365808,
-0.00549614522606134,
-0.00551111623644829,
-0.00552611798048019,
-0.00554115045815706,
-0.00555621366947889,
-0.00557130761444569,
-0.00558643275871873,
-0.00560158863663673,
-0.00561677524819970,
-0.00563199305906892,
-0.00564724160358310,
-0.00566252134740353,
-0.00567783229053021,
-0.00569317443296313,
-0.00570854777470231,
-0.00572395231574774,
-0.00573938805609942,
-0.00575485499575734,
-0.00577035360038281,
-0.00578588340431452,
-0.00580144440755248,
-0.00581703707575798,
-0.00583266140893102,
-0.00584831694141030,
-0.00586400413885713,
-0.00587972300127149,
-0.00589547352865338,
-0.00591125618666410,
-0.00592707050964236,
-0.00594291649758816,
-0.00595879461616278,
-0.00597470439970493,
-0.00599064631387591,
-0.00600661989301443,
-0.00602262560278177,
-0.00603866344317794,
-0.00605473341420293,
-0.00607083551585674,
-0.00608696974813938,
-0.00610313657671213,
-0.00611933553591371,
-0.00613556662574410,
-0.00615183031186461,
-0.00616812612861395,
-0.00618445454165340,
-0.00620081555098295,
-0.00621720915660262,
-0.00623363535851240,
-0.00625009415671229,
-0.00626658555120230,
-0.00628311000764370,
-0.00629966706037521,
-0.00631625670939684,
-0.00633287942036986,
-0.00634953519329429,
-0.00636622356250882,
-0.00638294499367476,
-0.00639969948679209,
-0.00641648704186082,
-0.00643330765888095,
-0.00645016133785248,
-0.00646704854443669,
-0.00648396881297231,
-0.00650092260912061,
-0.00651790946722031,
-0.00653492985293269,
-0.00655198376625776,
-0.00656907074153423,
-0.00658619124442339,
-0.00660334527492523,
-0.00662053329870105,
-0.00663775485008955,
-0.00665500992909074,
-0.00667229900136590,
-0.00668962160125375,
-0.00670697819441557,
-0.00672436831519008,
-0.00674179242923856,
-0.00675925053656101,
-0.00677674263715744,
-0.00679426873102784,
-0.00681182881817222,
-0.00682942289859057,
-0.00684705143794417,
-0.00686471397057176,
-0.00688241096213460,
-0.00690014194697142,
-0.00691790739074349,
-0.00693570729345083,
-0.00695354165509343,
-0.00697141047567129,
-0.00698931375518441,
-0.00700725149363279,
-0.00702522369101644,
-0.00704323081299663,
-0.00706127239391208,
-0.00707934889942408,
-0.00709746032953262,
-0.00711560621857643,
-0.00713378703221679,
-0.00715200277045369,
-0.00717025343328714,
-0.00718853902071714,
-0.00720685953274369,
-0.00722521543502808,
-0.00724360626190901,
-0.00726203247904778,
-0.00728049362078309,
-0.00729899015277624,
-0.00731752207502723,
-0.00733608938753605,
-0.00735469209030271,
-0.00737333018332720,
-0.00739200366660953,
-0.00741071254014969,
-0.00742945680394769,
-0.00744823692366481,
-0.00746705243363977,
-0.00748590379953384,
-0.00750479102134705,
-0.00752371409907937,
-0.00754267256706953,
-0.00756166689097881,
-0.00758069753646851,
-0.00759976403787732,
-0.00761886639520526,
-0.00763800460845232,
-0.00765717914327979,
-0.00767638999968767,
-0.00769563671201468,
-0.00771491974592209,
-0.00773423910140991,
-0.00775359477847815,
-0.00777298677712679,
-0.00779241509735584,
-0.00781187973916531,
-0.00783138070255518,
-0.00785091891884804,
-0.00787049345672131,
-0.00789010431617498,
-0.00790975149720907,
-0.00792943593114615,
-0.00794915668666363,
-0.00796891469508410,
-0.00798870902508497,
-0.00800854060798883,
-0.00802840944379568,
-0.00804831460118294,
-0.00806825701147318,
-0.00808823667466641,
-0.00810825359076262,
-0.00812830775976181,
-0.00814839918166399,
-0.00816852785646915,
-0.00818869378417730,
-0.00820889696478844,
-0.00822913739830256,
-0.00824941508471966,
-0.00826973002403975,
-0.00829008314758539,
-0.00831047352403402,
-0.00833090115338564,
-0.00835136696696281,
-0.00837187003344297,
-0.00839241128414869,
-0.00841298978775740,
-0.00843360647559166,
-0.00845426041632891,
-0.00847495254129171,
-0.00849568285048008,
-0.00851645134389401,
-0.00853725802153349,
-0.00855810195207596,
-0.00857898406684399,
-0.00859990436583757,
-0.00862086284905672,
-0.00864186044782400,
-0.00866289623081684,
-0.00868397019803524,
-0.00870508234947920,
-0.00872623268514872,
-0.00874742213636637,
-0.00876864977180958,
-0.00878991559147835,
-0.00881122052669525,
-0.00883256364613771,
-0.00885394588112831,
-0.00887536723166704,
-0.00889682676643133,
-0.00891832541674376,
-0.00893986318260431,
-0.00896144006401300,
-0.00898305606096983,
-0.00900471024215221,
-0.00902640353888273,
-0.00904813595116139,
-0.00906990841031075,
-0.00909171998500824,
-0.00911357067525387,
-0.00913546048104763,
-0.00915738940238953,
-0.00917935837060213,
-0.00920136645436287,
-0.00922341365367174,
-0.00924550089985132,
-0.00926762726157904,
-0.00928979367017746,
-0.00931199919432402,
-0.00933424476534128,
-0.00935653038322926,
-0.00937885604798794,
-0.00940122082829475,
-0.00942362565547228,
-0.00944607052952051,
-0.00946855545043945,
-0.00949108041822910,
-0.00951364543288946,
-0.00953625049442053,
-0.00955889560282230,
-0.00958158168941736,
-0.00960430782288313,
-0.00962707400321960,
-0.00964988023042679,
-0.00967272743582726,
-0.00969561468809843,
-0.00971854291856289,
-0.00974151119589806,
-0.00976452045142651,
-0.00978757068514824,
-0.00981066096574068,
-0.00983379222452641,
-0.00985696446150541,
-0.00988017767667770,
-0.00990343187004328,
-0.00992672704160214,
-0.00995006319135428,
-0.00997344031929970,
-0.00999685842543840,
-0.0100203175097704,
-0.0100438175722957,
-0.0100673595443368,
-0.0100909424945712,
-0.0101145664229989,
-0.0101382322609425,
-0.0101619390770793,
-0.0101856878027320,
-0.0102094775065780,
-0.0102333091199398,
-0.0102571826428175,
-0.0102810971438885,
-0.0103050535544753,
-0.0103290518745780,
-0.0103530921041965,
-0.0103771742433310,
-0.0104012982919812,
-0.0104254642501473,
-0.0104496721178293,
-0.0104739218950272,
-0.0104982135817409,
-0.0105225471779704,
-0.0105469236150384,
-0.0105713419616222,
-0.0105958031490445,
-0.0106203062459826,
-0.0106448512524366,
-0.0106694390997291,
-0.0106940697878599,
-0.0107187423855066,
-0.0107434578239918,
-0.0107682161033154,
-0.0107930172234774,
-0.0108178602531552,
-0.0108427461236715,
-0.0108676748350263,
-0.0108926463872194,
-0.0109176607802510,
-0.0109427189454436,
-0.0109678199514747,
-0.0109929637983441,
-0.0110181504860520,
-0.0110433809459209,
-0.0110686542466283,
-0.0110939703881741,
-0.0111193303018808,
-0.0111447330564260,
-0.0111701795831323,
-0.0111956698819995,
-0.0112212030217052,
-0.0112467799335718,
-0.0112724006175995,
-0.0112980650737882,
-0.0113237733021379,
-0.0113495253026485,
-0.0113753210753202,
-0.0114011606201530,
-0.0114270439371467,
-0.0114529710263014,
-0.0114789418876171,
-0.0115049565210938,
-0.0115310158580542,
-0.0115571189671755,
-0.0115832658484578,
-0.0116094574332237,
-0.0116356927901506,
-0.0116619728505611,
-0.0116882976144552,
-0.0117146661505103,
-0.0117410793900490,
-0.0117675373330712,
-0.0117940399795771,
-0.0118205863982439,
-0.0118471775203943,
-0.0118738133460283,
-0.0119004938751459,
-0.0119272191077471,
-0.0119539899751544,
-0.0119808055460453,
-0.0120076658204198,
-0.0120345707982779,
-0.0120615214109421,
-0.0120885167270899,
-0.0121155567467213,
-0.0121426424011588,
-0.0121697736904025,
-0.0121969496831298,
-0.0122241713106632,
-0.0122514385730028,
-0.0122787505388260,
-0.0123061081394553,
-0.0123335113748908,
-0.0123609602451324,
-0.0123884547501802,
-0.0124159948900342,
-0.0124435806646943,
-0.0124712120741606,
-0.0124988891184330,
-0.0125266127288342,
-0.0125543819740415,
-0.0125821968540549,
-0.0126100583001971,
-0.0126379653811455,
-0.0126659190282226,
-0.0126939183101058,
-0.0127219641581178,
-0.0127500556409359,
-0.0127781936898828,
-0.0128063783049583,
-0.0128346094861627,
-0.0128628863021731,
-0.0128912096843123,
-0.0129195796325803,
-0.0129479961469769,
-0.0129764592275023,
-0.0130049698054791,
-0.0130335269495845,
-0.0130621306598187,
-0.0130907809361815,
-0.0131194787099957,
-0.0131482230499387,
-0.0131770139560103,
-0.0132058523595333,
-0.0132347382605076,
-0.0132636707276106,
-0.0132926506921649,
-0.0133216781541705,
-0.0133507521823049,
-0.0133798737078905,
-0.0134090427309275,
-0.0134382592514157,
-0.0134675232693553,
-0.0134968347847462,
-0.0135261937975883,
-0.0135556003078818,
-0.0135850543156266,
-0.0136145567521453,
-0.0136441066861153,
-0.0136737041175365,
-0.0137033499777317,
-0.0137330433353782,
-0.0137627851217985,
-0.0137925744056702,
-0.0138224121183157,
-0.0138522982597351,
-0.0138822318986058,
-0.0139122139662504,
-0.0139422444626689,
-0.0139723233878613,
-0.0140024507418275,
-0.0140326265245676,
-0.0140628507360816,
-0.0140931233763695,
-0.0141234444454312,
-0.0141538148745894,
-0.0141842337325215,
-0.0142147010192275,
-0.0142452176660299,
-0.0142757827416062,
-0.0143063971772790,
-0.0143370600417256,
-0.0143677722662687,
-0.0143985338509083,
-0.0144293438643217,
-0.0144602032378316,
-0.0144911119714379,
-0.0145220700651407,
-0.0145530775189400,
-0.0145841343328357,
-0.0146152405068278,
-0.0146463960409164,
-0.0146776009351015,
-0.0147088561207056,
-0.0147401606664062,
-0.0147715145722032,
-0.0148029187694192,
-0.0148343723267317,
-0.0148658761754632,
-0.0148974293842912,
-0.0149290328845382,
-0.0149606866762042,
-0.0149923907592893,
-0.0150241442024708,
-0.0150559479370713,
-0.0150878019630909,
-0.0151197062805295,
-0.0151516608893871,
-0.0151836657896638,
-0.0152157209813595,
-0.0152478273957968,
-0.0152799841016531,
-0.0153121910989285,
-0.0153444493189454,
-0.0153767578303814,
-0.0154091175645590,
-0.0154415275901556,
-0.0154739888384938,
-0.0155065003782511,
-0.0155390631407499,
-0.0155716771259904,
-0.0156043423339725,
-0.0156370587646961,
-0.0156698264181614,
-0.0157026443630457,
-0.0157355144619942,
-0.0157684348523617,
-0.0158014073967934,
-0.0158344320952892,
-0.0158675070852041,
-0.0159006342291832,
-0.0159338135272264,
-0.0159670431166887,
-0.0160003248602152,
-0.0160336587578058,
-0.0160670448094606,
-0.0161004830151796,
-0.0161339733749628,
-0.0161675140261650,
-0.0162011068314314,
-0.0162347517907619,
-0.0162684489041567,
-0.0163021981716156,
-0.0163359995931387,
-0.0163698550313711,
-0.0164037626236677,
-0.0164377223700285,
-0.0164717342704535,
-0.0165057983249426,
-0.0165399145334959,
-0.0165740847587585,
-0.0166083071380854,
-0.0166425816714764,
-0.0166769102215767,
-0.0167112909257412,
-0.0167457237839699,
-0.0167802106589079,
-0.0168147496879101,
-0.0168493427336216,
-0.0168839879333973,
-0.0169186871498823,
-0.0169534403830767,
-0.0169882457703352,
-0.0170231051743031,
-0.0170580185949802,
-0.0170929841697216,
-0.0171280037611723,
-0.0171630773693323,
-0.0171982049942017,
-0.0172333847731352,
-0.0172686185687780,
-0.0173039063811302,
-0.0173392482101917,
-0.0173746440559626,
-0.0174100939184427,
-0.0174455977976322,
-0.0174811556935310,
-0.0175167676061392,
-0.0175524335354567,
-0.0175881534814835,
-0.0176239274442196,
-0.0176597572863102,
-0.0176956411451101,
-0.0177315790206194,
-0.0177675709128380,
-0.0178036186844111,
-0.0178397204726934,
-0.0178758762776852,
-0.0179120879620314,
-0.0179483536630869,
-0.0179846752434969,
-0.0180210508406162,
-0.0180574823170900,
-0.0180939678102732,
-0.0181305091828108,
-0.0181671045720577,
-0.0182037558406591,
-0.0182404629886150,
-0.0182772241532803,
-0.0183140411973000,
-0.0183509141206741,
-0.0183878429234028,
-0.0184248276054859,
-0.0184618663042784,
-0.0184989608824253,
-0.0185361113399267,
-0.0185733176767826,
-0.0186105798929930,
-0.0186478979885578,
-0.0186852719634771,
-0.0187227018177509,
-0.0187601875513792,
-0.0187977310270071,
-0.0188353303819895,
-0.0188729856163263,
-0.0189106967300177,
-0.0189484637230635,
-0.0189862884581089,
-0.0190241690725088,
-0.0190621055662632,
-0.0191000998020172,
-0.0191381499171257,
-0.0191762577742338,
-0.0192144215106964,
-0.0192526429891586,
-0.0192909203469753,
-0.0193292554467917,
-0.0193676464259624,
-0.0194060951471329,
-0.0194446016103029,
-0.0194831639528275,
-0.0195217840373516,
-0.0195604618638754,
-0.0195991974323988,
-0.0196379907429218,
-0.0196768399327993,
-0.0197157468646765,
-0.0197547115385532,
-0.0197937339544296,
-0.0198328141123056,
-0.0198719520121813,
-0.0199111476540566,
-0.0199504010379314,
-0.0199897121638060,
-0.0200290828943253,
-0.0200685113668442,
-0.0201079975813627,
-0.0201475415378809,
-0.0201871432363987,
-0.0202268045395613,
-0.0202665235847235,
-0.0203063022345305,
-0.0203461386263371,
-0.0203860327601433,
-0.0204259864985943,
-0.0204659979790449,
-0.0205060690641403,
-0.0205461978912354,
-0.0205863863229752,
-0.0206266343593597,
-0.0206669401377440,
-0.0207073055207729,
-0.0207477305084467,
-0.0207882132381201,
-0.0208287555724382,
-0.0208693575114012,
-0.0209100190550089,
-0.0209507402032614,
-0.0209915209561586,
-0.0210323613137007,
-0.0210732612758875,
-0.0211142208427191,
-0.0211552400141954,
-0.0211963187903166,
-0.0212374571710825,
-0.0212786551564932,
-0.0213199127465487,
-0.0213612299412489,
-0.0214026086032391,
-0.0214440468698740,
-0.0214855447411537,
-0.0215271040797234,
-0.0215687230229378,
-0.0216104015707970,
-0.0216521415859461,
-0.0216939412057400,
-0.0217358022928238,
-0.0217777229845524,
-0.0218197051435709,
-0.0218617469072342,
-0.0219038501381874,
-0.0219460148364306,
-0.0219882391393185,
-0.0220305249094963,
-0.0220728721469641,
-0.0221152808517218,
-0.0221577491611242,
-0.0222002789378166,
-0.0222428701817989,
-0.0222855228930712,
-0.0223282370716333,
-0.0223710127174854,
-0.0224138498306274,
-0.0224567484110594,
-0.0224997084587812,
-0.0225427299737930,
-0.0225858129560947,
-0.0226289592683315,
-0.0226721670478582,
-0.0227154362946749,
-0.0227587670087814,
-0.0228021610528231,
-0.0228456165641546,
-0.0228891335427761,
-0.0229327138513327,
-0.0229763556271791,
-0.0230200607329607,
-0.0230638273060322,
-0.0231076572090387,
-0.0231515485793352,
-0.0231955032795668,
-0.0232395213097334,
-0.0232836008071899,
-0.0233277436345816,
-0.0233719497919083,
-0.0234162192791700,
-0.0234605502337217,
-0.0235049445182085,
-0.0235494021326303,
-0.0235939230769873,
-0.0236385073512793,
-0.0236831549555063,
-0.0237278658896685,
-0.0237726401537657,
-0.0238174777477980,
-0.0238623786717653,
-0.0239073429256678,
-0.0239523723721504,
-0.0239974651485682,
-0.0240426212549210,
-0.0240878406912088,
-0.0241331253200769,
-0.0241784732788801,
-0.0242238845676184,
-0.0242693610489368,
-0.0243149008601904,
-0.0243605058640242,
-0.0244061741977930,
-0.0244519077241421,
-0.0244977045804262,
-0.0245435666292906,
-0.0245894938707352,
-0.0246354844421148,
-0.0246815402060747,
-0.0247276611626148,
-0.0247738473117352,
-0.0248200967907906,
-0.0248664114624262,
-0.0249127913266420,
-0.0249592363834381,
-0.0250057466328144,
-0.0250523220747709,
-0.0250989627093077,
-0.0251456685364246,
-0.0251924395561218,
-0.0252392757683992,
-0.0252861790359020,
-0.0253331474959850,
-0.0253801811486483,
-0.0254272799938917,
-0.0254744458943605,
-0.0255216769874096,
-0.0255689732730389,
-0.0256163366138935,
-0.0256637651473284,
-0.0257112607359886,
-0.0257588215172291,
-0.0258064493536949,
-0.0258541423827410,
-0.0259019024670124,
-0.0259497296065092,
-0.0259976219385862,
-0.0260455813258886,
-0.0260936077684164,
-0.0261416994035244,
-0.0261898580938578,
-0.0262380838394165,
-0.0262863766402006,
-0.0263347364962101,
-0.0263831634074450,
-0.0264316573739052,
-0.0264802183955908,
-0.0265288464725018,
-0.0265775416046381,
-0.0266263037919998,
-0.0266751330345869,
-0.0267240311950445,
-0.0267729964107275,
-0.0268220286816359,
-0.0268711280077696,
-0.0269202962517738,
-0.0269695315510035,
-0.0270188357681036,
-0.0270682070404291,
-0.0271176453679800,
-0.0271671526134014,
-0.0272167287766933,
-0.0272663719952106,
-0.0273160841315985,
-0.0273658633232117,
-0.0274157114326954,
-0.0274656284600496,
-0.0275156144052744,
-0.0275656674057245,
-0.0276157893240452,
-0.0276659801602364,
-0.0277162399142981,
-0.0277665685862303,
-0.0278169661760330,
-0.0278674326837063,
-0.0279179681092501,
-0.0279685724526644,
-0.0280192457139492,
-0.0280699878931046,
-0.0281207989901304,
-0.0281716790050268,
-0.0282226298004389,
-0.0282736495137215,
-0.0283247381448746,
-0.0283758975565434,
-0.0284271258860827,
-0.0284784231334925,
-0.0285297911614180,
-0.0285812281072140,
-0.0286327358335257,
-0.0286843124777079,
-0.0287359599024057,
-0.0287876762449741,
-0.0288394633680582,
-0.0288913212716579,
-0.0289432499557734,
-0.0289952475577593,
-0.0290473159402609,
-0.0290994551032782,
-0.0291516650468111,
-0.0292039457708597,
-0.0292562972754240,
-0.0293087195605040,
-0.0293612126260996,
-0.0294137764722109,
-0.0294664110988379,
-0.0295191165059805,
-0.0295718926936388,
-0.0296247396618128,
-0.0296776574105024,
-0.0297306459397078,
-0.0297837071120739,
-0.0298368390649557,
-0.0298900417983532,
-0.0299433171749115,
-0.0299966633319855,
-0.0300500821322203,
-0.0301035717129707,
-0.0301571339368820,
-0.0302107669413090,
-0.0302644725888968,
-0.0303182490170002,
-0.0303720980882645,
-0.0304260198026896,
-0.0304800122976303,
-0.0305340774357319,
-0.0305882152169943,
-0.0306424256414175,
-0.0306967087090015,
-0.0307510625571013,
-0.0308054890483618,
-0.0308599881827831,
-0.0309145599603653,
-0.0309692043811083,
-0.0310239214450121,
-0.0310787111520767,
-0.0311335753649473,
-0.0311885122209787,
-0.0312435217201710,
-0.0312986038625240,
-0.0313537605106831,
-0.0314089879393578,
-0.0314642898738384,
-0.0315196663141251,
-0.0315751135349274,
-0.0316306352615356,
-0.0316862314939499,
-0.0317419022321701,
-0.0317976437509060,
-0.0318534597754478,
-0.0319093503057957,
-0.0319653153419495,
-0.0320213548839092,
-0.0320774689316750,
-0.0321336537599564,
-0.0321899130940437,
-0.0322462469339371,
-0.0323026552796364,
-0.0323591381311417,
-0.0324156954884529,
-0.0324723273515701,
-0.0325290337204933,
-0.0325858145952225,
-0.0326426699757576,
-0.0326995998620987,
-0.0327566042542458,
-0.0328136831521988,
-0.0328708365559578,
-0.0329280681908131,
-0.0329853743314743,
-0.0330427549779415,
-0.0331002101302147,
-0.0331577397882938,
-0.0332153439521790,
-0.0332730263471603,
-0.0333307832479477,
-0.0333886146545410,
-0.0334465205669403,
-0.0335045047104359,
-0.0335625633597374,
-0.0336206965148449,
-0.0336789079010487,
-0.0337371937930584,
-0.0337955541908741,
-0.0338539928197861,
-0.0339125059545040,
-0.0339710973203182,
-0.0340297631919384,
-0.0340885072946548,
-0.0341473259031773,
-0.0342062227427959,
-0.0342651940882206,
-0.0343242436647415,
-0.0343833677470684,
-0.0344425700604916,
-0.0345018468797207,
-0.0345612019300461,
-0.0346206352114677,
-0.0346801429986954,
-0.0347397290170193,
-0.0347993932664394,
-0.0348591320216656,
-0.0349189490079880,
-0.0349788442254067,
-0.0350388176739216,
-0.0350988656282425,
-0.0351589918136597,
-0.0352191962301731,
-0.0352794788777828,
-0.0353398397564888,
-0.0354002788662910,
-0.0354607924818993,
-0.0355213843286037,
-0.0355820544064045,
-0.0356428027153015,
-0.0357036292552948,
-0.0357645340263844,
-0.0358255170285702,
-0.0358865782618523,
-0.0359477177262306,
-0.0360089354217052,
-0.0360702313482761,
-0.0361316055059433,
-0.0361930578947067,
-0.0362545922398567,
-0.0363162048161030,
-0.0363778956234455,
-0.0364396646618843,
-0.0365015119314194,
-0.0365634374320507,
-0.0366254448890686,
-0.0366875305771828,
-0.0367496944963932,
-0.0368119403719902,
-0.0368742644786835,
-0.0369366668164730,
-0.0369991473853588,
-0.0370617099106312,
-0.0371243506669998,
-0.0371870733797550,
-0.0372498743236065,
-0.0373127534985542,
-0.0373757146298885,
-0.0374387539923191,
-0.0375018753111362,
-0.0375650748610497,
-0.0376283563673496,
-0.0376917161047459,
-0.0377551577985287,
-0.0378186814486980,
-0.0378822833299637,
-0.0379459671676159,
-0.0380097292363644,
-0.0380735732614994,
-0.0381374992430210,
-0.0382015034556389,
-0.0382655896246433,
-0.0383297577500343,
-0.0383940078318119,
-0.0384583361446857,
-0.0385227464139462,
-0.0385872386395931,
-0.0386518128216267,
-0.0387164689600468,
-0.0387812070548534,
-0.0388460233807564,
-0.0389109216630459,
-0.0389759019017220,
-0.0390409640967846,
-0.0391061082482338,
-0.0391713343560696,
-0.0392366424202919,
-0.0393020324409008,
-0.0393675044178963,
-0.0394330583512783,
-0.0394986942410469,
-0.0395644120872021,
-0.0396302118897438,
-0.0396960973739624,
-0.0397620648145676,
-0.0398281142115593,
-0.0398942455649376,
-0.0399604588747025,
-0.0400267541408539,
-0.0400931350886822,
-0.0401595979928970,
-0.0402261428534985,
-0.0402927696704865,
-0.0403594821691513,
-0.0404262766242027,
-0.0404931530356407,
-0.0405601151287556,
-0.0406271591782570,
-0.0406942889094353,
-0.0407615005970001,
-0.0408287942409515,
-0.0408961735665798,
-0.0409636348485947,
-0.0410311818122864,
-0.0410988107323647,
-0.0411665253341198,
-0.0412343256175518,
-0.0413022078573704,
-0.0413701757788658,
-0.0414382256567478,
-0.0415063612163067,
-0.0415745824575424,
-0.0416428856551647,
-0.0417112745344639,
-0.0417797490954399,
-0.0418483056128025,
-0.0419169478118420,
-0.0419856756925583,
-0.0420544892549515,
-0.0421233847737312,
-0.0421923659741879,
-0.0422614328563213,
-0.0423305854201317,
-0.0423998236656189,
-0.0424691475927830,
-0.0425385572016239,
-0.0426080524921417,
-0.0426776334643364,
-0.0427473001182079,
-0.0428170487284660,
-0.0428868867456913,
-0.0429568104445934,
-0.0430268198251724,
-0.0430969148874283,
-0.0431670956313610,
-0.0432373620569706,
-0.0433077141642571,
-0.0433781519532204,
-0.0434486754238606,
-0.0435192883014679,
-0.0435899868607521,
-0.0436607711017132,
-0.0437316410243511,
-0.0438025966286659,
-0.0438736416399479,
-0.0439447723329067,
-0.0440159887075424,
-0.0440872944891453,
-0.0441586859524250,
-0.0442301630973816,
-0.0443017296493053,
-0.0443733818829060,
-0.0444451235234737,
-0.0445169508457184,
-0.0445888675749302,
-0.0446608699858189,
-0.0447329618036747,
-0.0448051393032074,
-0.0448774062097073,
-0.0449497587978840,
-0.0450222007930279,
-0.0450947321951389,
-0.0451673492789269,
-0.0452400557696819,
-0.0453128516674042,
-0.0453857332468033,
-0.0454587042331696,
-0.0455317646265030,
-0.0456049144268036,
-0.0456781499087811,
-0.0457514747977257,
-0.0458248890936375,
-0.0458983927965164,
-0.0459719859063625,
-0.0460456684231758,
-0.0461194366216660,
-0.0461932942271233,
-0.0462672412395477,
-0.0463412776589394,
-0.0464154034852982,
-0.0464896187186241,
-0.0465639233589172,
-0.0466383174061775,
-0.0467128008604050,
-0.0467873774468899,
-0.0468620434403420,
-0.0469367988407612,
-0.0470116436481476,
-0.0470865778625011,
-0.0471616014838219,
-0.0472367145121098,
-0.0473119206726551,
-0.0473872162401676,
-0.0474626012146473,
-0.0475380793213844,
-0.0476136468350887,
-0.0476893037557602,
-0.0477650538086891,
-0.0478408932685852,
-0.0479168221354485,
-0.0479928441345692,
-0.0480689555406570,
-0.0481451600790024,
-0.0482214540243149,
-0.0482978411018848,
-0.0483743175864220,
-0.0484508872032166,
-0.0485275462269783,
-0.0486042983829975,
-0.0486811399459839,
-0.0487580746412277,
-0.0488351024687290,
-0.0489122197031975,
-0.0489894300699234,
-0.0490667335689068,
-0.0491441264748573,
-0.0492216125130653,
-0.0492991916835308,
-0.0493768639862537,
-0.0494546256959438,
-0.0495324805378914,
-0.0496104285120964,
-0.0496884696185589,
-0.0497666038572788,
-0.0498448312282562,
-0.0499231517314911,
-0.0500015616416931,
-0.0500800646841526,
-0.0501586608588696,
-0.0502373501658440,
-0.0503161326050758,
-0.0503950081765652,
-0.0504739806056023,
-0.0505530461668968,
-0.0506322048604488,
-0.0507114566862583,
-0.0507908016443253,
-0.0508702397346497,
-0.0509497709572315,
-0.0510293990373611,
-0.0511091202497482,
-0.0511889345943928,
-0.0512688420712948,
-0.0513488464057446,
-0.0514289438724518,
-0.0515091344714165,
-0.0515894219279289,
-0.0516698025166988,
-0.0517502762377262,
-0.0518308468163013,
-0.0519115105271339,
-0.0519922710955143,
-0.0520731247961521,
-0.0521540753543377,
-0.0522351190447807,
-0.0523162595927715,
-0.0523974932730198,
-0.0524788238108158,
-0.0525602474808693,
-0.0526417680084705,
-0.0527233853936195,
-0.0528050959110260,
-0.0528869032859802,
-0.0529688075184822,
-0.0530508048832417,
-0.0531328991055489,
-0.0532150901854038,
-0.0532973781228066,
-0.0533797629177570,
-0.0534622408449650,
-0.0535448156297207,
-0.0536274872720242,
-0.0537102557718754,
-0.0537931211292744,
-0.0538760833442211,
-0.0539591424167156,
-0.0540422983467579,
-0.0541255511343479,
-0.0542089007794857,
-0.0542923472821713,
-0.0543758906424046,
-0.0544595308601856,
-0.0545432679355145,
-0.0546271018683910,
-0.0547110326588154,
-0.0547950640320778,
-0.0548791922628880,
-0.0549634173512459,
-0.0550477392971516,
-0.0551321581006050,
-0.0552166774868965,
-0.0553012937307358,
-0.0553860068321228,
-0.0554708205163479,
-0.0555557310581207,
-0.0556407384574413,
-0.0557258464396000,
-0.0558110512793064,
-0.0558963567018509,
-0.0559817589819431,
-0.0560672618448734,
-0.0561528615653515,
-0.0562385618686676,
-0.0563243590295315,
-0.0564102567732334,
-0.0564962513744831,
-0.0565823465585709,
-0.0566685423254967,
-0.0567548349499702,
-0.0568412281572819,
-0.0569277219474316,
-0.0570143125951290,
-0.0571010038256645,
-0.0571877956390381,
-0.0572746880352497,
-0.0573616810142994,
-0.0574487708508968,
-0.0575359612703323,
-0.0576232522726059,
-0.0577106438577175,
-0.0577981360256672,
-0.0578857287764549,
-0.0579734221100807,
-0.0580612160265446,
-0.0581491105258465,
-0.0582371056079865,
-0.0583252012729645,
-0.0584133975207806,
-0.0585016943514347,
-0.0585900917649269,
-0.0586785897612572,
-0.0587671883404255,
-0.0588558912277222,
-0.0589446946978569,
-0.0590335987508297,
-0.0591226033866406,
-0.0592117123305798,
-0.0593009218573570,
-0.0593902319669724,
-0.0594796463847160,
-0.0595691613852978,
-0.0596587769687176,
-0.0597484968602657,
-0.0598383173346520,
-0.0599282421171665,
-0.0600182674825192,
-0.0601083971560001,
-0.0601986274123192,
-0.0602889619767666,
-0.0603793971240521,
-0.0604699365794659,
-0.0605605766177177,
-0.0606513209640980,
-0.0607421696186066,
-0.0608331188559532,
-0.0609241724014282,
-0.0610153302550316,
-0.0611065886914730,
-0.0611979514360428,
-0.0612894184887409,
-0.0613809898495674,
-0.0614726655185223,
-0.0615644417703152,
-0.0616563223302364,
-0.0617483071982861,
-0.0618403963744640,
-0.0619325898587704,
-0.0620248876512051,
-0.0621172897517681,
-0.0622097961604595,
-0.0623024068772793,
-0.0623951219022274,
-0.0624879412353039,
-0.0625808686017990,
-0.0626738965511322,
-0.0627670288085938,
-0.0628602653741837,
-0.0629536062479019,
-0.0630470514297485,
-0.0631406083703041,
-0.0632342696189880,
-0.0633280351758003,
-0.0634219050407410,
-0.0635158792138100,
-0.0636099576950073,
-0.0637041404843330,
-0.0637984350323677,
-0.0638928338885307,
-0.0639873370528221,
-0.0640819445252419,
-0.0641766563057900,
-0.0642714798450470,
-0.0643664076924324,
-0.0644614398479462,
-0.0645565837621689,
-0.0646518319845200,
-0.0647471845149994,
-0.0648426413536072,
-0.0649382099509239,
-0.0650338828563690,
-0.0651296600699425,
-0.0652255490422249,
-0.0653215423226357,
-0.0654176399111748,
-0.0655138492584229,
-0.0656101629137993,
-0.0657065883278847,
-0.0658031180500984,
-0.0658997595310211,
-0.0659965053200722,
-0.0660933554172516,
-0.0661903172731400,
-0.0662873834371567,
-0.0663845613598824,
-0.0664818435907364,
-0.0665792375802994,
-0.0666767358779907,
-0.0667743459343910,
-0.0668720602989197,
-0.0669698864221573,
-0.0670678243041039,
-0.0671658664941788,
-0.0672640204429627,
-0.0673622786998749,
-0.0674606487154961,
-0.0675591304898262,
-0.0676577165722847,
-0.0677564144134522,
-0.0678552240133286,
-0.0679541379213333,
-0.0680531635880470,
-0.0681523010134697,
-0.0682515427470207,
-0.0683508962392807,
-0.0684503614902496,
-0.0685499310493469,
-0.0686496123671532,
-0.0687494054436684,
-0.0688493102788925,
-0.0689493268728256,
-0.0690494477748871,
-0.0691496804356575,
-0.0692500248551369,
-0.0693504810333252,
-0.0694510489702225,
-0.0695517212152481,
-0.0696525052189827,
-0.0697534009814262,
-0.0698544085025787,
-0.0699555277824402,
-0.0700567588210106,
-0.0701581016182900,
-0.0702595561742783,
-0.0703611224889755,
-0.0704628005623817,
-0.0705645903944969,
-0.0706664919853210,
-0.0707685053348541,
-0.0708706304430962,
-0.0709728673100472,
-0.0710752159357071,
-0.0711776763200760,
-0.0712802484631538,
-0.0713829323649406,
-0.0714857280254364,
-0.0715886354446411,
-0.0716916546225548,
-0.0717947855591774,
-0.0718980282545090,
-0.0720013827085495,
-0.0721048489212990,
-0.0722084343433380,
-0.0723121315240860,
-0.0724159404635429,
-0.0725198611617088,
-0.0726238936185837,
-0.0727280452847481,
-0.0728323087096214,
-0.0729366838932037,
-0.0730411708354950,
-0.0731457769870758,
-0.0732504948973656,
-0.0733553245663643,
-0.0734602659940720,
-0.0735653266310692,
-0.0736704990267754,
-0.0737757831811905,
-0.0738811865448952,
-0.0739867016673088,
-0.0740923285484314,
-0.0741980746388435,
-0.0743039324879646,
-0.0744099020957947,
-0.0745159909129143,
-0.0746221914887428,
-0.0747285112738609,
-0.0748349428176880,
-0.0749414935708046,
-0.0750481560826302,
-0.0751549378037453,
-0.0752618312835693,
-0.0753688365221024,
-0.0754759609699249,
-0.0755832046270371,
-0.0756905600428581,
-0.0757980346679688,
-0.0759056210517883,
-0.0760133266448975,
-0.0761211439967156,
-0.0762290805578232,
-0.0763371288776398,
-0.0764452964067459,
-0.0765535831451416,
-0.0766619816422463,
-0.0767704993486404,
-0.0768791362643242,
-0.0769878849387169,
-0.0770967528223991,
-0.0772057399153709,
-0.0773148387670517,
-0.0774240568280220,
-0.0775333940982819,
-0.0776428505778313,
-0.0777524188160896,
-0.0778621062636375,
-0.0779719129204750,
-0.0780818387866020,
-0.0781918764114380,
-0.0783020332455635,
-0.0784123092889786,
-0.0785227045416832,
-0.0786332190036774,
-0.0787438526749611,
-0.0788546055555344,
-0.0789654701948166,
-0.0790764540433884,
-0.0791875571012497,
-0.0792987793684006,
-0.0794101208448410,
-0.0795215815305710,
-0.0796331614255905,
-0.0797448605298996,
-0.0798566788434982,
-0.0799686163663864,
-0.0800806730985642,
-0.0801928490400314,
-0.0803051441907883,
-0.0804175585508347,
-0.0805300921201706,
-0.0806427448987961,
-0.0807555168867111,
-0.0808684080839157,
-0.0809814184904099,
-0.0810945481061935,
-0.0812078043818474,
-0.0813211798667908,
-0.0814346745610237,
-0.0815482884645462,
-0.0816620215773583,
-0.0817758738994598,
-0.0818898528814316,
-0.0820039510726929,
-0.0821181684732437,
-0.0822325050830841,
-0.0823469609022141,
-0.0824615433812141,
-0.0825762450695038,
-0.0826910659670830,
-0.0828060135245323,
-0.0829210802912712,
-0.0830362662672997,
-0.0831515714526177,
-0.0832670032978058,
-0.0833825543522835,
-0.0834982320666313,
-0.0836140289902687,
-0.0837299451231957,
-0.0838459879159927,
-0.0839621499180794,
-0.0840784385800362,
-0.0841948464512825,
-0.0843113735318184,
-0.0844280272722244,
-0.0845448002219200,
-0.0846616998314858,
-0.0847787186503410,
-0.0848958641290665,
-0.0850131288170815,
-0.0851305201649666,
-0.0852480307221413,
-0.0853656679391861,
-0.0854834318161011,
-0.0856013149023056,
-0.0857193246483803,
-0.0858374536037445,
-0.0859557092189789,
-0.0860740914940834,
-0.0861925929784775,
-0.0863112211227417,
-0.0864299759268761,
-0.0865488499403000,
-0.0866678506135941,
-0.0867869779467583,
-0.0869062244892120,
-0.0870255976915360,
-0.0871450975537300,
-0.0872647240757942,
-0.0873844698071480,
-0.0875043421983719,
-0.0876243412494659,
-0.0877444669604302,
-0.0878647118806839,
-0.0879850834608078,
-0.0881055817008019,
-0.0882262066006661,
-0.0883469581604004,
-0.0884678363800049,
-0.0885888412594795,
-0.0887099653482437,
-0.0888312160968781,
-0.0889525935053825,
-0.0890740975737572,
-0.0891957283020020,
-0.0893174856901169,
-0.0894393697381020,
-0.0895613804459572,
-0.0896835178136826,
-0.0898057818412781,
-0.0899281725287437,
-0.0900506898760796,
-0.0901733338832855,
-0.0902961045503616,
-0.0904190018773079,
-0.0905420258641243,
-0.0906651765108109,
-0.0907884612679482,
-0.0909118726849556,
-0.0910354107618332,
-0.0911590754985809,
-0.0912828668951988,
-0.0914067849516869,
-0.0915308296680450,
-0.0916550084948540,
-0.0917793139815331,
-0.0919037461280823,
-0.0920283049345017,
-0.0921529904007912,
-0.0922778099775314,
-0.0924027562141419,
-0.0925278291106224,
-0.0926530361175537,
-0.0927783697843552,
-0.0929038301110268,
-0.0930294245481491,
-0.0931551456451416,
-0.0932809934020042,
-0.0934069752693176,
-0.0935330837965012,
-0.0936593189835548,
-0.0937856882810593,
-0.0939121842384338,
-0.0940388143062592,
-0.0941655710339546,
-0.0942924544215202,
-0.0944194719195366,
-0.0945466160774231,
-0.0946738943457604,
-0.0948012992739677,
-0.0949288383126259,
-0.0950565040111542,
-0.0951843038201332,
-0.0953122302889824,
-0.0954402908682823,
-0.0955684855580330,
-0.0956968069076538,
-0.0958252623677254,
-0.0959538444876671,
-0.0960825607180595,
-0.0962114110589027,
-0.0963403880596161,
-0.0964694991707802,
-0.0965987443923950,
-0.0967281162738800,
-0.0968576222658157,
-0.0969872623682022,
-0.0971170291304588,
-0.0972469300031662,
-0.0973769649863243,
-0.0975071340799332,
-0.0976374298334122,
-0.0977678596973419,
-0.0978984236717224,
-0.0980291217565537,
-0.0981599539518356,
-0.0982909128069878,
-0.0984220057725906,
-0.0985532328486443,
-0.0986845940351486,
-0.0988160893321037,
-0.0989477187395096,
-0.0990794822573662,
-0.0992113798856735,
-0.0993434116244316,
-0.0994755700230598,
-0.0996078625321388,
-0.0997402891516686,
-0.0998728498816490,
-0.100005544722080,
-0.100138373672962,
-0.100271336734295,
-0.100404433906078,
-0.100537672638893,
-0.100671045482159,
-0.100804552435875,
-0.100938193500042,
-0.101071968674660,
-0.101205877959728,
-0.101339921355248,
-0.101474098861218,
-0.101608410477638,
-0.101742856204510,
-0.101877443492413,
-0.102012164890766,
-0.102147020399570,
-0.102282010018826,
-0.102417133748531,
-0.102552399039269,
-0.102687798440456,
-0.102823331952095,
-0.102958999574184,
-0.103094808757305,
-0.103230752050877,
-0.103366829454899,
-0.103503048419952,
-0.103639401495457,
-0.103775888681412,
-0.103912517428398,
-0.104049280285835,
-0.104186177253723,
-0.104323215782642,
-0.104460388422012,
-0.104597702622414,
-0.104735150933266,
-0.104872733354568,
-0.105010457336903,
-0.105148315429688,
-0.105286315083504,
-0.105424448847771,
-0.105562724173069,
-0.105701133608818,
-0.105839684605598,
-0.105978369712830,
-0.106117196381092,
-0.106256164610386,
-0.106395266950130,
-0.106534510850906,
-0.106673888862133,
-0.106813408434391,
-0.106953069567680,
-0.107092864811420,
-0.107232801616192,
-0.107372879981995,
-0.107513092458248,
-0.107653446495533,
-0.107793942093849,
-0.107934571802616,
-0.108075343072414,
-0.108216255903244,
-0.108357310295105,
-0.108498498797417,
-0.108639828860760,
-0.108781300485134,
-0.108922913670540,
-0.109064668416977,
-0.109206564724445,
-0.109348595142365,
-0.109490767121315,
-0.109633080661297,
-0.109775535762310,
-0.109918132424355,
-0.110060870647430,
-0.110203750431538,
-0.110346771776676,
-0.110489934682846,
-0.110633239150047,
-0.110776685178280,
-0.110920272767544,
-0.111064001917839,
-0.111207872629166,
-0.111351884901524,
-0.111496038734913,
-0.111640334129334,
-0.111784771084785,
-0.111929349601269,
-0.112074069678783,
-0.112218931317329,
-0.112363934516907,
-0.112509079277515,
-0.112654365599155,
-0.112799800932407,
-0.112945377826691,
-0.113091096282005,
-0.113236956298351,
-0.113382957875729,
-0.113529108464718,
-0.113675400614738,
-0.113821834325790,
-0.113968409597874,
-0.114115133881569,
-0.114261999726295,
-0.114409007132053,
-0.114556163549423,
-0.114703461527824,
-0.114850901067257,
-0.114998489618301,
-0.115146219730377,
-0.115294091403484,
-0.115442112088203,
-0.115590274333954,
-0.115738585591316,
-0.115887038409710,
-0.116035632789135,
-0.116184376180172,
-0.116333261132240,
-0.116482295095921,
-0.116631470620632,
-0.116780795156956,
-0.116930261254311,
-0.117079876363277,
-0.117229633033276,
-0.117379538714886,
-0.117529593408108,
-0.117679789662361,
-0.117830134928226,
-0.117980621755123,
-0.118131257593632,
-0.118282042443752,
-0.118432968854904,
-0.118584044277668,
-0.118735268712044,
-0.118886634707451,
-0.119038149714470,
-0.119189813733101,
-0.119341626763344,
-0.119493581354618,
-0.119645684957504,
-0.119797937572002,
-0.119950339198112,
-0.120102882385254,
-0.120255574584007,
-0.120408415794373,
-0.120561406016350,
-0.120714545249939,
-0.120867833495140,
-0.121021263301373,
-0.121174842119217,
-0.121328569948673,
-0.121482446789742,
-0.121636472642422,
-0.121790647506714,
-0.121944971382618,
-0.122099444270134,
-0.122254066169262,
-0.122408837080002,
-0.122563757002354,
-0.122718825936317,
-0.122874043881893,
-0.123029410839081,
-0.123184926807880,
-0.123340591788292,
-0.123496405780315,
-0.123652368783951,
-0.123808480799198,
-0.123964749276638,
-0.124121166765690,
-0.124277733266354,
-0.124434448778629,
-0.124591313302517,
-0.124748326838017,
-0.124905496835709,
-0.125062808394432,
-0.125220283865929,
-0.125377908349037,
-0.125535681843758,
-0.125693604350090,
-0.125851675868034,
-0.126009896397591,
-0.126168265938759,
-0.126326799392700,
-0.126485481858253,
-0.126644313335419,
-0.126803293824196,
-0.126962423324585,
-0.127121701836586,
-0.127281144261360,
-0.127440735697746,
-0.127600476145744,
-0.127760365605354,
-0.127920418977737,
-0.128080621361732,
-0.128240972757339,
-0.128401473164558,
-0.128562137484550,
-0.128722950816154,
-0.128883913159370,
-0.129045024514198,
-0.129206299781799,
-0.129367724061012,
-0.129529297351837,
-0.129691019654274,
-0.129852905869484,
-0.130014941096306,
-0.130177125334740,
-0.130339473485947,
-0.130501970648766,
-0.130664616823196,
-0.130827426910400,
-0.130990386009216,
-0.131153494119644,
-0.131316766142845,
-0.131480187177658,
-0.131643772125244,
-0.131807506084442,
-0.131971389055252,
-0.132135435938835,
-0.132299631834030,
-0.132463991641998,
-0.132628500461578,
-0.132793158292770,
-0.132957980036736,
-0.133122950792313,
-0.133288085460663,
-0.133453369140625,
-0.133618816733360,
-0.133784413337708,
-0.133950173854828,
-0.134116083383560,
-0.134282156825066,
-0.134448379278183,
-0.134614765644074,
-0.134781301021576,
-0.134948000311852,
-0.135114848613739,
-0.135281860828400,
-0.135449022054672,
-0.135616347193718,
-0.135783821344376,
-0.135951459407806,
-0.136119246482849,
-0.136287197470665,
-0.136455312371254,
-0.136623576283455,
-0.136792004108429,
-0.136960580945015,
-0.137129321694374,
-0.137298226356506,
-0.137467280030251,
-0.137636497616768,
-0.137805864214897,
-0.137975394725800,
-0.138145089149475,
-0.138314932584763,
-0.138484939932823,
-0.138655111193657,
-0.138825431466103,
-0.138995915651321,
-0.139166563749313,
-0.139337360858917,
-0.139508321881294,
-0.139679446816444,
-0.139850735664368,
-0.140022173523903,
-0.140193775296211,
-0.140365540981293,
-0.140537455677986,
-0.140709534287453,
-0.140881776809692,
-0.141054183244705,
-0.141226738691330,
-0.141399458050728,
-0.141572341322899,
-0.141745388507843,
-0.141918599605560,
-0.142091959714890,
-0.142265483736992,
-0.142439171671867,
-0.142613023519516,
-0.142787039279938,
-0.142961204051971,
-0.143135532736778,
-0.143310025334358,
-0.143484681844711,
-0.143659502267838,
-0.143834486603737,
-0.144009634852409,
-0.144184932112694,
-0.144360393285751,
-0.144536018371582,
-0.144711807370186,
-0.144887760281563,
-0.145063877105713,
-0.145240157842636,
-0.145416602492332,
-0.145593211054802,
-0.145769983530045,
-0.145946919918060,
-0.146124005317688,
-0.146301254630089,
-0.146478667855263,
-0.146656244993210,
-0.146833986043930,
-0.147011891007423,
-0.147189959883690,
-0.147368192672730,
-0.147546589374542,
-0.147725149989128,
-0.147903874516487,
-0.148082762956619,
-0.148261815309525,
-0.148441031575203,
-0.148620426654816,
-0.148799985647202,
-0.148979708552361,
-0.149159595370293,
-0.149339646100998,
-0.149519860744476,
-0.149700239300728,
-0.149880781769753,
-0.150061488151550,
-0.150242358446121,
-0.150423392653465,
-0.150604590773582,
-0.150785967707634,
-0.150967508554459,
-0.151149213314056,
-0.151331081986427,
-0.151513114571571,
-0.151695311069489,
-0.151877671480179,
-0.152060210704803,
-0.152242913842201,
-0.152425780892372,
-0.152608811855316,
-0.152792006731033,
-0.152975380420685,
-0.153158918023109,
-0.153342619538307,
-0.153526484966278,
-0.153710529208183,
-0.153894737362862,
-0.154079109430313,
-0.154263645410538,
-0.154448360204697,
-0.154633238911629,
-0.154818281531334,
-0.155003488063812,
-0.155188873410225,
-0.155374422669411,
-0.155560135841370,
-0.155746027827263,
-0.155932083725929,
-0.156118303537369,
-0.156304702162743,
-0.156491264700890,
-0.156677991151810,
-0.156864896416664,
-0.157051965594292,
-0.157239198684692,
-0.157426610589027,
-0.157614186406136,
-0.157801926136017,
-0.157989844679832,
-0.158177927136421,
-0.158366188406944,
-0.158554613590240,
-0.158743202686310,
-0.158931970596313,
-0.159120902419090,
-0.159310013055801,
-0.159499287605286,
-0.159688740968704,
-0.159878358244896,
-0.160068154335022,
-0.160258114337921,
-0.160448238253593,
-0.160638540983200,
-0.160829007625580,
-0.161019653081894,
-0.161210462450981,
-0.161401450634003,
-0.161592617630959,
-0.161783948540688,
-0.161975458264351,
-0.162167131900787,
-0.162358984351158,
-0.162551000714302,
-0.162743195891380,
-0.162935554981232,
-0.163128092885017,
-0.163320809602737,
-0.163513690233231,
-0.163706749677658,
-0.163899973034859,
-0.164093375205994,
-0.164286956191063,
-0.164480701088905,
-0.164674624800682,
-0.164868712425232,
-0.165062978863716,
-0.165257424116135,
-0.165452033281326,
-0.165646821260452,
-0.165841788053513,
-0.166036918759346,
-0.166232228279114,
-0.166427716612816,
-0.166623368859291,
-0.166819199919701,
-0.167015209794045,
-0.167211398482323,
-0.167407751083374,
-0.167604282498360,
-0.167800992727280,
-0.167997881770134,
-0.168194934725761,
-0.168392166495323,
-0.168589577078819,
-0.168787166476250,
-0.168984919786453,
-0.169182851910591,
-0.169380962848663,
-0.169579252600670,
-0.169777721166611,
-0.169976353645325,
-0.170175164937973,
-0.170374155044556,
-0.170573323965073,
-0.170772671699524,
-0.170972198247910,
-0.171171888709068,
-0.171371757984161,
-0.171571806073189,
-0.171772032976151,
-0.171972438693047,
-0.172173023223877,
-0.172373786568642,
-0.172574728727341,
-0.172775849699974,
-0.172977134585381,
-0.173178598284721,
-0.173380240797997,
-0.173582062125206,
-0.173784062266350,
-0.173986241221428,
-0.174188598990440,
-0.174391135573387,
-0.174593850970268,
-0.174796745181084,
-0.174999818205833,
-0.175203070044518,
-0.175406500697136,
-0.175610110163689,
-0.175813898444176,
-0.176017865538597,
-0.176222011446953,
-0.176426336169243,
-0.176630839705467,
-0.176835522055626,
-0.177040383219719,
-0.177245423197746,
-0.177450641989708,
-0.177656054496765,
-0.177861645817757,
-0.178067415952683,
-0.178273364901543,
-0.178479492664337,
-0.178685799241066,
-0.178892284631729,
-0.179098948836327,
-0.179305791854858,
-0.179512828588486,
-0.179720044136047,
-0.179927438497543,
-0.180135011672974,
-0.180342763662338,
-0.180550694465637,
-0.180758818984032,
-0.180967122316360,
-0.181175604462624,
-0.181384265422821,
-0.181593105196953,
-0.181802138686180,
-0.182011350989342,
-0.182220742106438,
-0.182430312037468,
-0.182640075683594,
-0.182850018143654,
-0.183060139417648,
-0.183270439505577,
-0.183480933308601,
-0.183691605925560,
-0.183902457356453,
-0.184113502502441,
-0.184324726462364,
-0.184536129236221,
-0.184747710824013,
-0.184959486126900,
-0.185171440243721,
-0.185383573174477,
-0.185595899820328,
-0.185808405280113,
-0.186021104454994,
-0.186233982443810,
-0.186447039246559,
-0.186660289764404,
-0.186873719096184,
-0.187087327241898,
-0.187301129102707,
-0.187515109777451,
-0.187729284167290,
-0.187943637371063,
-0.188158184289932,
-0.188372910022736,
-0.188587814569473,
-0.188802912831306,
-0.189018189907074,
-0.189233660697937,
-0.189449310302734,
-0.189665153622627,
-0.189881175756454,
-0.190097391605377,
-0.190313786268234,
-0.190530374646187,
-0.190747141838074,
-0.190964102745056,
-0.191181242465973,
-0.191398575901985,
-0.191616103053093,
-0.191833809018135,
-0.192051708698273,
-0.192269787192345,
-0.192488059401512,
-0.192706510424614,
-0.192925155162811,
-0.193143993616104,
-0.193363010883331,
-0.193582221865654,
-0.193801611661911,
-0.194021195173264,
-0.194240972399712,
-0.194460928440094,
-0.194681078195572,
-0.194901421666145,
-0.195121943950653,
-0.195342659950256,
-0.195563569664955,
-0.195784658193588,
-0.196005940437317,
-0.196227416396141,
-0.196449071168900,
-0.196670919656754,
-0.196892961859703,
-0.197115197777748,
-0.197337612509727,
-0.197560220956802,
-0.197783023118973,
-0.198006018996239,
-0.198229193687439,
-0.198452562093735,
-0.198676124215126,
-0.198899880051613,
-0.199123829603195,
-0.199347957968712,
-0.199572280049324,
-0.199796795845032,
-0.200021505355835,
-0.200246408581734,
-0.200471505522728,
-0.200696781277657,
-0.200922250747681,
-0.201147913932800,
-0.201373770833015,
-0.201599821448326,
-0.201826065778732,
-0.202052503824234,
-0.202279135584831,
-0.202505946159363,
-0.202732950448990,
-0.202960148453712,
-0.203187540173531,
-0.203415125608444,
-0.203642904758453,
-0.203870877623558,
-0.204099044203758,
-0.204327404499054,
-0.204555958509445,
-0.204784706234932,
-0.205013647675514,
-0.205242782831192,
-0.205472111701965,
-0.205701634287834,
-0.205931350588799,
-0.206161260604858,
-0.206391364336014,
-0.206621661782265,
-0.206852152943611,
-0.207082837820053,
-0.207313716411591,
-0.207544788718224,
-0.207776054739952,
-0.208007514476776,
-0.208239182829857,
-0.208471044898033,
-0.208703100681305,
-0.208935350179672,
-0.209167793393135,
-0.209400430321693,
-0.209633260965347,
-0.209866285324097,
-0.210099518299103,
-0.210332944989204,
-0.210566565394402,
-0.210800379514694,
-0.211034387350082,
-0.211268588900566,
-0.211502999067307,
-0.211737602949142,
-0.211972400546074,
-0.212207391858101,
-0.212442576885223,
-0.212677970528603,
-0.212913557887077,
-0.213149338960648,
-0.213385313749313,
-0.213621497154236,
-0.213857874274254,
-0.214094445109367,
-0.214331224560738,
-0.214568197727203,
-0.214805364608765,
-0.215042725205421,
-0.215280294418335,
-0.215518057346344,
-0.215756013989449,
-0.215994179248810,
-0.216232538223267,
-0.216471105813980,
-0.216709867119789,
-0.216948822140694,
-0.217187985777855,
-0.217427343130112,
-0.217666894197464,
-0.217906653881073,
-0.218146607279778,
-0.218386769294739,
-0.218627125024796,
-0.218867689371109,
-0.219108447432518,
-0.219349399209023,
-0.219590559601784,
-0.219831913709641,
-0.220073476433754,
-0.220315232872963,
-0.220557197928429,
-0.220799356698990,
-0.221041724085808,
-0.221284285187721,
-0.221527054905891,
-0.221770018339157,
-0.222013190388680,
-0.222256556153297,
-0.222500130534172,
-0.222743898630142,
-0.222987875342369,
-0.223232060670853,
-0.223476439714432,
-0.223721027374268,
-0.223965808749199,
-0.224210798740387,
-0.224455997347832,
-0.224701389670372,
-0.224946990609169,
-0.225192785263062,
-0.225438788533211,
-0.225685000419617,
-0.225931406021118,
-0.226178020238876,
-0.226424843072891,
-0.226671859622002,
-0.226919084787369,
-0.227166518568993,
-0.227414146065712,
-0.227661982178688,
-0.227910026907921,
-0.228158280253410,
-0.228406727313995,
-0.228655382990837,
-0.228904247283936,
-0.229153320193291,
-0.229402586817741,
-0.229652062058449,
-0.229901745915413,
-0.230151638388634,
-0.230401724576950,
-0.230652019381523,
-0.230902522802353,
-0.231153234839439,
-0.231404155492783,
-0.231655269861221,
-0.231906592845917,
-0.232158124446869,
-0.232409864664078,
-0.232661813497543,
-0.232913970947266,
-0.233166337013245,
-0.233418896794319,
-0.233671665191650,
-0.233924642205238,
-0.234177827835083,
-0.234431222081184,
-0.234684824943542,
-0.234938636422157,
-0.235192656517029,
-0.235446885228157,
-0.235701322555542,
-0.235955968499184,
-0.236210823059082,
-0.236465886235237,
-0.236721158027649,
-0.236976638436317,
-0.237232327461243,
-0.237488225102425,
-0.237744331359863,
-0.238000646233559,
-0.238257169723511,
-0.238513901829720,
-0.238770842552185,
-0.239027991890907,
-0.239285349845886,
-0.239542916417122,
-0.239800691604614,
-0.240058675408363,
-0.240316867828369,
-0.240575268864632,
-0.240833878517151,
-0.241092711687088,
-0.241351753473282,
-0.241611003875732,
-0.241870462894440,
-0.242130130529404,
-0.242390006780624,
-0.242650091648102,
-0.242910400032997,
-0.243170917034149,
-0.243431642651558,
-0.243692576885223,
-0.243953719735146,
-0.244215086102486,
-0.244476661086082,
-0.244738444685936,
-0.245000436902046,
-0.245262652635574,
-0.245525076985359,
-0.245787709951401,
-0.246050551533699,
-0.246313616633415,
-0.246576890349388,
-0.246840372681618,
-0.247104063630104,
-0.247367978096008,
-0.247632101178169,
-0.247896432876587,
-0.248160988092422,
-0.248425751924515,
-0.248690724372864,
-0.248955920338631,
-0.249221324920654,
-0.249486938118935,
-0.249752774834633,
-0.250018835067749,
-0.250285089015961,
-0.250551581382751,
-0.250818282365799,
-0.251085191965103,
-0.251352310180664,
-0.251619637012482,
-0.251887202262878,
-0.252154976129532,
-0.252422958612442,
-0.252691149711609,
-0.252959549427032,
-0.253228187561035,
-0.253497034311295,
-0.253766089677811,
-0.254035353660584,
-0.254304856061935,
-0.254574567079544,
-0.254844486713409,
-0.255114644765854,
-0.255385011434555,
-0.255655586719513,
-0.255926370620728,
-0.256197392940521,
-0.256468623876572,
-0.256740063428879,
-0.257011741399765,
-0.257283627986908,
-0.257555723190308,
-0.257828027009964,
-0.258100569248199,
-0.258373320102692,
-0.258646279573441,
-0.258919477462769,
-0.259192883968353,
-0.259466499090195,
-0.259740352630615,
-0.260014414787293,
-0.260288685560226,
-0.260563194751740,
-0.260837912559509,
-0.261112838983536,
-0.261388003826141,
-0.261663377285004,
-0.261938989162445,
-0.262214809656143,
-0.262490838766098,
-0.262767106294632,
-0.263043582439423,
-0.263320267200470,
-0.263597190380096,
-0.263874322175980,
-0.264151692390442,
-0.264429271221161,
-0.264707058668137,
-0.264985084533691,
-0.265263319015503,
-0.265541791915894,
-0.265820473432541,
-0.266099393367767,
-0.266378521919251,
-0.266657859086990,
-0.266937434673309,
-0.267217218875885,
-0.267497241497040,
-0.267777472734451,
-0.268057942390442,
-0.268338620662689,
-0.268619537353516,
-0.268900662660599,
-0.269181996583939,
-0.269463568925858,
-0.269745349884033,
-0.270027369260788,
-0.270309597253799,
-0.270592063665390,
-0.270874738693237,
-0.271157652139664,
-0.271440774202347,
-0.271724134683609,
-0.272007703781128,
-0.272291511297226,
-0.272575527429581,
-0.272859781980515,
-0.273144274950027,
-0.273428976535797,
-0.273713916540146,
-0.273999065160751,
-0.274284452199936,
-0.274570047855377,
-0.274855881929398,
-0.275141924619675,
-0.275428205728531,
-0.275714695453644,
-0.276001423597336,
-0.276288390159607,
-0.276575565338135,
-0.276862978935242,
-0.277150601148605,
-0.277438461780548,
-0.277726560831070,
-0.278014868497849,
-0.278303414583206,
-0.278592169284821,
-0.278881162405014,
-0.279170393943787,
-0.279459834098816,
-0.279749512672424,
-0.280039399862289,
-0.280329525470734,
-0.280619889497757,
-0.280910462141037,
-0.281201273202896,
-0.281492322683334,
-0.281783580780029,
-0.282075077295303,
-0.282366812229157,
-0.282658755779266,
-0.282950937747955,
-0.283243358135223,
-0.283535987138748,
-0.283828854560852,
-0.284121960401535,
-0.284415274858475,
-0.284708827733994,
-0.285002619028091,
-0.285296618938446,
-0.285590857267380,
-0.285885334014893,
-0.286180019378662,
-0.286474943161011,
-0.286770105361939,
-0.287065505981445,
-0.287361115217209,
-0.287656962871552,
-0.287953048944473,
-0.288249373435974,
-0.288545906543732,
-0.288842678070068,
-0.289139688014984,
-0.289436936378479,
-0.289734393358231,
-0.290032088756561,
-0.290330022573471,
-0.290628194808960,
-0.290926575660706,
-0.291225194931030,
-0.291524052619934,
-0.291823148727417,
-0.292122483253479,
-0.292422026395798,
-0.292721807956696,
-0.293021827936173,
-0.293322086334229,
-0.293622583150864,
-0.293923288583756,
-0.294224232435226,
-0.294525414705277,
-0.294826835393906,
-0.295128494501114,
-0.295430392026901,
-0.295732498168945,
-0.296034842729569,
-0.296337425708771,
-0.296640247106552,
-0.296943306922913,
-0.297246605157852,
-0.297550112009048,
-0.297853857278824,
-0.298157840967178,
-0.298462063074112,
-0.298766523599625,
-0.299071222543716,
-0.299376159906387,
-0.299681335687637,
-0.299986749887466,
-0.300292372703552,
-0.300598233938217,
-0.300904333591461,
-0.301210671663284,
-0.301517248153687,
-0.301824063062668,
-0.302131116390228,
-0.302438408136368,
-0.302745938301086,
-0.303053706884384,
-0.303361713886261,
-0.303669959306717,
-0.303978443145752,
-0.304287165403366,
-0.304596126079559,
-0.304905295372009,
-0.305214703083038,
-0.305524349212647,
-0.305834233760834,
-0.306144356727600,
-0.306454718112946,
-0.306765317916870,
-0.307076156139374,
-0.307387232780457,
-0.307698547840118,
-0.308010101318359,
-0.308321893215179,
-0.308633923530579,
-0.308946192264557,
-0.309258699417114,
-0.309571444988251,
-0.309884428977966,
-0.310197681188583,
-0.310511171817780,
-0.310824900865555,
-0.311138868331909,
-0.311453074216843,
-0.311767518520355,
-0.312082201242447,
-0.312397122383118,
-0.312712281942368,
-0.313027679920197,
-0.313343316316605,
-0.313659191131592,
-0.313975304365158,
-0.314291656017303,
-0.314608246088028,
-0.314925104379654,
-0.315242201089859,
-0.315559536218643,
-0.315877109766006,
-0.316194921731949,
-0.316512972116470,
-0.316831260919571,
-0.317149788141251,
-0.317468583583832,
-0.317787617444992,
-0.318106889724731,
-0.318426400423050,
-0.318746149539948,
-0.319066137075424,
-0.319386363029480,
-0.319706857204437,
-0.320027589797974,
-0.320348560810089,
-0.320669770240784,
-0.320991218090057,
-0.321312904357910,
-0.321634858846664,
-0.321957051753998,
-0.322279483079910,
-0.322602152824402,
-0.322925060987473,
-0.323248237371445,
-0.323571652173996,
-0.323895305395126,
-0.324219197034836,
-0.324543356895447,
-0.324867755174637,
-0.325192391872406,
-0.325517266988754,
-0.325842380523682,
-0.326167762279511,
-0.326493382453918,
-0.326819241046906,
-0.327145338058472,
-0.327471703290939,
-0.327798306941986,
-0.328125149011612,
-0.328452259302139,
-0.328779608011246,
-0.329107195138931,
-0.329435020685196,
-0.329763114452362,
-0.330091446638107,
-0.330420017242432,
-0.330748856067657,
-0.331077933311462,
-0.331407248973846,
-0.331736832857132,
-0.332066655158997,
-0.332396715879440,
-0.332727044820786,
-0.333057612180710,
-0.333388417959213,
-0.333719491958618,
-0.334050804376602,
-0.334382355213165,
-0.334714174270630,
-0.335046231746674,
-0.335378527641296,
-0.335711091756821,
-0.336043894290924,
-0.336376965045929,
-0.336710274219513,
-0.337043821811676,
-0.337377637624741,
-0.337711691856384,
-0.338045984506607,
-0.338380545377731,
-0.338715344667435,
-0.339050412178040,
-0.339385718107224,
-0.339721292257309,
-0.340057104825974,
-0.340393155813217,
-0.340729475021362,
-0.341066032648087,
-0.341402858495712,
-0.341739922761917,
-0.342077255249023,
-0.342414826154709,
-0.342752665281296,
-0.343090742826462,
-0.343429088592529,
-0.343767672777176,
-0.344106495380402,
-0.344445586204529,
-0.344784915447235,
-0.345124512910843,
-0.345464348793030,
-0.345804452896118,
-0.346144795417786,
-0.346485406160355,
-0.346826255321503,
-0.347167372703552,
-0.347508758306503,
-0.347850382328033,
-0.348192274570465,
-0.348534405231476,
-0.348876804113388,
-0.349219441413879,
-0.349562346935272,
-0.349905490875244,
-0.350248903036118,
-0.350592553615570,
-0.350936472415924,
-0.351280659437180,
-0.351625084877014,
-0.351969778537750,
-0.352314710617065,
-0.352659910917282,
-0.353005349636078,
-0.353351056575775,
-0.353697031736374,
-0.354043245315552,
-0.354389727115631,
-0.354736447334290,
-0.355083435773850,
-0.355430692434311,
-0.355778187513351,
-0.356125950813293,
-0.356473982334137,
-0.356822252273560,
-0.357170790433884,
-0.357519596815109,
-0.357868641614914,
-0.358217954635620,
-0.358567535877228,
-0.358917355537415,
-0.359267443418503,
-0.359617799520493,
-0.359968394041061,
-0.360319256782532,
-0.360670387744904,
-0.361021757125855,
-0.361373394727707,
-0.361725300550461,
-0.362077444791794,
-0.362429857254028,
-0.362782537937164,
-0.363135457038879,
-0.363488644361496,
-0.363842099905014,
-0.364195823669434,
-0.364549785852432,
-0.364904016256332,
-0.365258514881134,
-0.365613281726837,
-0.365968286991119,
-0.366323560476303,
-0.366679102182388,
-0.367034912109375,
-0.367390960454941,
-0.367747277021408,
-0.368103861808777,
-0.368460714817047,
-0.368817806243897,
-0.369175165891647,
-0.369532793760300,
-0.369890689849854,
-0.370248854160309,
-0.370607256889343,
-0.370965927839279,
-0.371324867010117,
-0.371684074401855,
-0.372043550014496,
-0.372403264045715,
-0.372763246297836,
-0.373123496770859,
-0.373484015464783,
-0.373844802379608,
-0.374205857515335,
-0.374567151069641,
-0.374928712844849,
-0.375290542840958,
-0.375652641057968,
-0.376015007495880,
-0.376377642154694,
-0.376740545034409,
-0.377103686332703,
-0.377467095851898,
-0.377830773591995,
-0.378194719552994,
-0.378558933734894,
-0.378923416137695,
-0.379288166761398,
-0.379653185606003,
-0.380018472671509,
-0.380383998155594,
-0.380749791860580,
-0.381115853786469,
-0.381482183933258,
-0.381848782300949,
-0.382215648889542,
-0.382582783699036,
-0.382950186729431,
-0.383317857980728,
-0.383685797452927,
-0.384054005146027,
-0.384422481060028,
-0.384791225194931,
-0.385160237550736,
-0.385529518127441,
-0.385899066925049,
-0.386268883943558,
-0.386638939380646,
-0.387009263038635,
-0.387379854917526,
-0.387750715017319,
-0.388121843338013,
-0.388493239879608,
-0.388864904642105,
-0.389236837625504,
-0.389609038829803,
-0.389981508255005,
-0.390354245901108,
-0.390727251768112,
-0.391100525856018,
-0.391474068164825,
-0.391847908496857,
-0.392222017049789,
-0.392596393823624,
-0.392971038818359,
-0.393345952033997,
-0.393721133470535,
-0.394096583127975,
-0.394472301006317,
-0.394848287105560,
-0.395224541425705,
-0.395601063966751,
-0.395977854728699,
-0.396354913711548,
-0.396732240915298,
-0.397109836339951,
-0.397487699985504,
-0.397865831851959,
-0.398244261741638,
-0.398622959852219,
-0.399001926183701,
-0.399381160736084,
-0.399760663509369,
-0.400140434503555,
-0.400520473718643,
-0.400900781154633,
-0.401281356811523,
-0.401662230491638,
-0.402043372392654,
-0.402424782514572,
-0.402806460857391,
-0.403188407421112,
-0.403570622205734,
-0.403953105211258,
-0.404335886240006,
-0.404718935489655,
-0.405102252960205,
-0.405485838651657,
-0.405869692564011,
-0.406253814697266,
-0.406638205051422,
-0.407022893428803,
-0.407407850027084,
-0.407793074846268,
-0.408178567886353,
-0.408564329147339,
-0.408950388431549,
-0.409336715936661,
-0.409723311662674,
-0.410110175609589,
-0.410497307777405,
-0.410884737968445,
-0.411272436380386,
-0.411660403013229,
-0.412048637866974,
-0.412437170743942,
-0.412825971841812,
-0.413215041160584,
-0.413604378700256,
-0.413993984460831,
-0.414383888244629,
-0.414774060249329,
-0.415164500474930,
-0.415555208921433,
-0.415946215391159,
-0.416337490081787,
-0.416729032993317,
-0.417120873928070,
-0.417512983083725,
-0.417905360460281,
-0.418298006057739,
-0.418690949678421,
-0.419084161520004,
-0.419477641582489,
-0.419871419668198,
-0.420265465974808,
-0.420659780502319,
-0.421054363250732,
-0.421449244022369,
-0.421844393014908,
-0.422239810228348,
-0.422635525465012,
-0.423031508922577,
-0.423427760601044,
-0.423824310302734,
-0.424221128225327,
-0.424618214368820,
-0.425015598535538,
-0.425413250923157,
-0.425811171531677,
-0.426209390163422,
-0.426607877016068,
-0.427006632089615,
-0.427405685186386,
-0.427805006504059,
-0.428204625844955,
-0.428604513406754,
-0.429004669189453,
-0.429405122995377,
-0.429805845022202,
-0.430206865072250,
-0.430608153343201,
-0.431009709835053,
-0.431411564350128,
-0.431813687086105,
-0.432216107845306,
-0.432618796825409,
-0.433021754026413,
-0.433425009250641,
-0.433828532695770,
-0.434232354164124,
-0.434636443853378,
-0.435040801763535,
-0.435445457696915,
-0.435850381851196,
-0.436255604028702,
-0.436661094427109,
-0.437066882848740,
-0.437472939491272,
-0.437879294157028,
-0.438285917043686,
-0.438692837953568,
-0.439100027084351,
-0.439507484436035,
-0.439915239810944,
-0.440323263406754,
-0.440731585025787,
-0.441140174865723,
-0.441549062728882,
-0.441958218812943,
-0.442367672920227,
-0.442777395248413,
-0.443187415599823,
-0.443597704172134,
-0.444008290767670,
-0.444419145584106,
-0.444830298423767,
-0.445241719484329,
-0.445653438568115,
-0.446065425872803,
-0.446477711200714,
-0.446890294551849,
-0.447303146123886,
-0.447716295719147,
-0.448129713535309,
-0.448543429374695,
-0.448957413434982,
-0.449371695518494,
-0.449786245822907,
-0.450201094150543,
-0.450616210699081,
-0.451031625270844,
-0.451447337865829,
-0.451863318681717,
-0.452279597520828,
-0.452696144580841,
-0.453112989664078,
-0.453530132770538,
-0.453947544097900,
-0.454365253448486,
-0.454783231019974,
-0.455201506614685,
-0.455620080232620,
-0.456038922071457,
-0.456458061933517,
-0.456877470016480,
-0.457297176122665,
-0.457717180252075,
-0.458137452602387,
-0.458558022975922,
-0.458978891372681,
-0.459400027990341,
-0.459821462631226,
-0.460243165493012,
-0.460665166378021,
-0.461087465286255,
-0.461510032415390,
-0.461932897567749,
-0.462356060743332,
-0.462779492139816,
-0.463203221559525,
-0.463627249002457,
-0.464051544666290,
-0.464476138353348,
-0.464901030063629,
-0.465326189994812,
-0.465751647949219,
-0.466177403926849,
-0.466603457927704,
-0.467029780149460,
-0.467456400394440,
-0.467883318662643,
-0.468310505151749,
-0.468737989664078,
-0.469165772199631,
-0.469593852758408,
-0.470022201538086,
-0.470450848340988,
-0.470879793167114,
-0.471309006214142,
-0.471738517284393,
-0.472168326377869,
-0.472598433494568,
-0.473028808832169,
-0.473459482192993,
-0.473890453577042,
-0.474321722984314,
-0.474753260612488,
-0.475185096263886,
-0.475617229938507,
-0.476049661636353,
-0.476482391357422,
-0.476915389299393,
-0.477348685264587,
-0.477782279253006,
-0.478216171264648,
-0.478650361299515,
-0.479084819555283,
-0.479519575834274,
-0.479954630136490,
-0.480389982461929,
-0.480825632810593,
-0.481261551380157,
-0.481697767972946,
-0.482134282588959,
-0.482571095228195,
-0.483008205890656,
-0.483445584774017,
-0.483883261680603,
-0.484321236610413,
-0.484759509563446,
-0.485198080539703,
-0.485636949539185,
-0.486076116561890,
-0.486515551805496,
-0.486955285072327,
-0.487395316362381,
-0.487835645675659,
-0.488276273012161,
-0.488717198371887,
-0.489158421754837,
-0.489599913358688,
-0.490041702985764,
-0.490483790636063,
-0.490926176309586,
-0.491368860006332,
-0.491811841726303,
-0.492255121469498,
-0.492698699235916,
-0.493142575025558,
-0.493586748838425,
-0.494031190872192,
-0.494475930929184,
-0.494920969009399,
-0.495366305112839,
-0.495811939239502,
-0.496257871389389,
-0.496704101562500,
-0.497150629758835,
-0.497597455978394,
-0.498044580221176,
-0.498492002487183,
-0.498939722776413,
-0.499387741088867,
-0.499836057424545,
-0.500284671783447,
-0.500733554363251,
-0.501182734966278,
-0.501632213592529,
-0.502081990242004,
-0.502532064914703,
-0.502982437610626,
-0.503433108329773,
-0.503884077072144,
-0.504335343837738,
-0.504786908626556,
-0.505238771438599,
-0.505690932273865,
-0.506143391132355,
-0.506596148014069,
-0.507049202919006,
-0.507502555847168,
-0.507956206798554,
-0.508410155773163,
-0.508864402770996,
-0.509318947792053,
-0.509773790836334,
-0.510228931903839,
-0.510684370994568,
-0.511140108108521,
-0.511596143245697,
-0.512052476406097,
-0.512509107589722,
-0.512966036796570,
-0.513423264026642,
-0.513880789279938,
-0.514338672161102,
-0.514796853065491,
-0.515255331993103,
-0.515714108943939,
-0.516173183917999,
-0.516632556915283,
-0.517092227935791,
-0.517552196979523,
-0.518012464046478,
-0.518473029136658,
-0.518933892250061,
-0.519395053386688,
-0.519856512546539,
-0.520318269729614,
-0.520780324935913,
-0.521242678165436,
-0.521705329418182,
-0.522168278694153,
-0.522631525993347,
-0.523095071315765,
-0.523558974266052,
-0.524023175239563,
-0.524487674236298,
-0.524952471256256,
-0.525417566299439,
-0.525882959365845,
-0.526348650455475,
-0.526814639568329,
-0.527280926704407,
-0.527747511863709,
-0.528214395046234,
-0.528681576251984,
-0.529149055480957,
-0.529616832733154,
-0.530084967613220,
-0.530553400516510,
-0.531022131443024,
-0.531491160392761,
-0.531960487365723,
-0.532430112361908,
-0.532900035381317,
-0.533370256423950,
-0.533840775489807,
-0.534311592578888,
-0.534782767295837,
-0.535254240036011,
-0.535726010799408,
-0.536198079586029,
-0.536670446395874,
-0.537143111228943,
-0.537616074085236,
-0.538089334964752,
-0.538562893867493,
-0.539036810398102,
-0.539511024951935,
-0.539985537528992,
-0.540460348129273,
-0.540935456752777,
-0.541410863399506,
-0.541886568069458,
-0.542362570762634,
-0.542838931083679,
-0.543315589427948,
-0.543792545795441,
-0.544269800186157,
-0.544747352600098,
-0.545225203037262,
-0.545703351497650,
-0.546181857585907,
-0.546660661697388,
-0.547139763832092,
-0.547619163990021,
-0.548098862171173,
-0.548578858375549,
-0.549059152603149,
-0.549539804458618,
-0.550020754337311,
-0.550502002239227,
-0.550983548164368,
-0.551465392112732,
-0.551947534084320,
-0.552430033683777,
-0.552912831306458,
-0.553395926952362,
-0.553879320621491,
-0.554363012313843,
-0.554847002029419,
-0.555331349372864,
-0.555815994739533,
-0.556300938129425,
-0.556786179542542,
-0.557271718978882,
-0.557757556438446,
-0.558243751525879,
-0.558730244636536,
-0.559217035770416,
-0.559704124927521,
-0.560191512107849,
-0.560679256916046,
-0.561167299747467,
-0.561655640602112,
-0.562144279479981,
-0.562633216381073,
-0.563122510910034,
-0.563612103462219,
-0.564101994037628,
-0.564592182636261,
-0.565082669258118,
-0.565573513507843,
-0.566064655780792,
-0.566556096076965,
-0.567047834396362,
-0.567539870738983,
-0.568032264709473,
-0.568524956703186,
-0.569017946720123,
-0.569511234760284,
-0.570004880428314,
-0.570498824119568,
-0.570993065834045,
-0.571487605571747,
-0.571982443332672,
-0.572477638721466,
-0.572973132133484,
-0.573468923568726,
-0.573965013027191,
-0.574461460113525,
-0.574958205223084,
-0.575455248355866,
-0.575952589511871,
-0.576450288295746,
-0.576948285102844,
-0.577446579933167,
-0.577945172786713,
-0.578444063663483,
-0.578943312168121,
-0.579442858695984,
-0.579942703247070,
-0.580442845821381,
-0.580943346023560,
-0.581444144248962,
-0.581945240497589,
-0.582446694374085,
-0.582948446273804,
-0.583450496196747,
-0.583952844142914,
-0.584455549716950,
-0.584958553314209,
-0.585461854934692,
-0.585965454578400,
-0.586469411849976,
-0.586973667144775,
-0.587478220462799,
-0.587983071804047,
-0.588488280773163,
-0.588993787765503,
-0.589499592781067,
-0.590005755424500,
-0.590512216091156,
-0.591018974781036,
-0.591526031494141,
-0.592033445835114,
-0.592541158199310,
-0.593049168586731,
-0.593557536602020,
-0.594066202640533,
-0.594575166702271,
-0.595084428787231,
-0.595594048500061,
-0.596103966236115,
-0.596614181995392,
-0.597124755382538,
-0.597635626792908,
-0.598146796226502,
-0.598658323287964,
-0.599170148372650,
-0.599682271480560,
-0.600194752216339,
-0.600707530975342,
-0.601220607757568,
-0.601733982563019,
-0.602247714996338,
-0.602761745452881,
-0.603276073932648,
-0.603790760040283,
-0.604305744171143,
-0.604821026325226,
-0.605336666107178,
-0.605852603912354,
-0.606368839740753,
-0.606885433197022,
-0.607402324676514,
-0.607919514179230,
-0.608437061309815,
-0.608954906463623,
-0.609473049640656,
-0.609991550445557,
-0.610510349273682,
-0.611029446125031,
-0.611548900604248,
-0.612068653106690,
-0.612588703632355,
-0.613109111785889,
-0.613629817962647,
-0.614150822162628,
-0.614672183990479,
-0.615193843841553,
-0.615715861320496,
-0.616238176822662,
-0.616760790348053,
-0.617283761501312,
-0.617807030677795,
-0.618330597877502,
-0.618854522705078,
-0.619378745555878,
-0.619903266429901,
-0.620428144931793,
-0.620953321456909,
-0.621478855609894,
-0.622004687786102,
-0.622530817985535,
-0.623057305812836,
-0.623584091663361,
-0.624111175537109,
-0.624638617038727,
-0.625166356563568,
-0.625694453716278,
-0.626222848892212,
-0.626751542091370,
-0.627280592918396,
-0.627809941768646,
-0.628339648246765,
-0.628869652748108,
-0.629399955272675,
-0.629930615425110,
-0.630461573600769,
-0.630992889404297,
-0.631524503231049,
-0.632056415081024,
-0.632588684558868,
-0.633121252059937,
-0.633654177188873,
-0.634187400341034,
-0.634720921516419,
-0.635254800319672,
-0.635788977146149,
-0.636323511600494,
-0.636858344078064,
-0.637393474578857,
-0.637928962707520,
-0.638464748859406,
-0.639000892639160,
-0.639537334442139,
-0.640074133872986,
-0.640611231327057,
-0.641148626804352,
-0.641686379909515,
-0.642224431037903,
-0.642762839794159,
-0.643301546573639,
-0.643840610980988,
-0.644379973411560,
-0.644919633865356,
-0.645459651947022,
-0.645999968051910,
-0.646540641784668,
-0.647081613540649,
-0.647622942924500,
-0.648164570331574,
-0.648706495761871,
-0.649248778820038,
-0.649791359901428,
-0.650334298610687,
-0.650877535343170,
-0.651421129703522,
-0.651965022087097,
-0.652509272098541,
-0.653053820133209,
-0.653598725795746,
-0.654143929481506,
-0.654689431190491,
-0.655235290527344,
-0.655781447887421,
-0.656327962875366,
-0.656874775886536,
-0.657421946525574,
-0.657969415187836,
-0.658517241477966,
-0.659065365791321,
-0.659613847732544,
-0.660162627696991,
-0.660711765289307,
-0.661261200904846,
-0.661810994148254,
-0.662361085414887,
-0.662911534309387,
-0.663462281227112,
-0.664013385772705,
-0.664564788341522,
-0.665116488933563,
-0.665668547153473,
-0.666220903396606,
-0.666773617267609,
-0.667326629161835,
-0.667879998683929,
-0.668433666229248,
-0.668987691402435,
-0.669542014598846,
-0.670096695423126,
-0.670651674270630,
-0.671207010746002,
-0.671762645244598,
-0.672318637371063,
-0.672874927520752,
-0.673431575298309,
-0.673988521099091,
-0.674545824527741,
-0.675103425979614,
-0.675661385059357,
-0.676219642162323,
-0.676778256893158,
-0.677337229251862,
-0.677896499633789,
-0.678456127643585,
-0.679016053676605,
-0.679576337337494,
-0.680136919021606,
-0.680697858333588,
-0.681259095668793,
-0.681820690631867,
-0.682382583618164,
-0.682944834232330,
-0.683507382869721,
-0.684070289134979,
-0.684633493423462,
-0.685197055339813,
-0.685760915279388,
-0.686325132846832,
-0.686889648437500,
-0.687454521656036,
-0.688019752502441,
-0.688585281372070,
-0.689151167869568,
-0.689717352390289,
-0.690283894538879,
-0.690850734710693,
-0.691417932510376,
-0.691985428333283,
-0.692553281784058,
-0.693121433258057,
-0.693689942359924,
-0.694258809089661,
-0.694827973842621,
-0.695397496223450,
-0.695967316627502,
-0.696537494659424,
-0.697107970714569,
-0.697678804397583,
-0.698249936103821,
-0.698821425437927,
-0.699393272399902,
-0.699965417385101,
-0.700537919998169,
-0.701110720634460,
-0.701683878898621,
-0.702257335186005,
-0.702831149101257,
-0.703405320644379,
-0.703979790210724,
-0.704554617404938,
-0.705129742622376,
-0.705705225467682,
-0.706281006336212,
-0.706857144832611,
-0.707433640956879,
-0.708010435104370,
-0.708587586879730,
-0.709165036678314,
-0.709742844104767,
-0.710320949554443,
-0.710899412631989,
-0.711478233337402,
-0.712057352066040,
-0.712636828422546,
-0.713216602802277,
-0.713796734809876,
-0.714377224445343,
-0.714958012104034,
-0.715539157390595,
-0.716120600700378,
-0.716702401638031,
-0.717284560203552,
-0.717867016792297,
-0.718449831008911,
-0.719032943248749,
-0.719616413116455,
-0.720200240612030,
-0.720784366130829,
-0.721368849277496,
-0.721953630447388,
-0.722538769245148,
-0.723124265670776,
-0.723710060119629,
-0.724296212196350,
-0.724882662296295,
-0.725469470024109,
-0.726056635379791,
-0.726644098758698,
-0.727231919765472,
-0.727820038795471,
-0.728408515453339,
-0.728997349739075,
-0.729586482048035,
-0.730175971984863,
-0.730765819549561,
-0.731355965137482,
-0.731946468353272,
-0.732537269592285,
-0.733128428459168,
-0.733719944953919,
-0.734311759471893,
-0.734903931617737,
-0.735496461391449,
-0.736089289188385,
-0.736682474613190,
-0.737275958061218,
-0.737869799137116,
-0.738463997840881,
-0.739058494567871,
-0.739653348922730,
-0.740248560905457,
-0.740844070911408,
-0.741439938545227,
-0.742036163806915,
-0.742632687091827,
-0.743229568004608,
-0.743826806545258,
-0.744424343109131,
-0.745022237300873,
-0.745620429515839,
-0.746218979358673,
-0.746817886829376,
-0.747417092323303,
-0.748016655445099,
-0.748616576194763,
-0.749216794967651,
-0.749817371368408,
-0.750418305397034,
-0.751019537448883,
-0.751621127128601,
-0.752223074436188,
-0.752825319766998,
-0.753427922725678,
-0.754030883312225,
-0.754634141921997,
-0.755237758159638,
-0.755841732025147,
-0.756446003913879,
-0.757050633430481,
-0.757655620574951,
-0.758260905742645,
-0.758866548538208,
-0.759472548961639,
-0.760078847408295,
-0.760685503482819,
-0.761292517185211,
-0.761899828910828,
-0.762507498264313,
-0.763115525245667,
-0.763723850250244,
-0.764332532882690,
-0.764941573143005,
-0.765550911426544,
-0.766160607337952,
-0.766770660877228,
-0.767381012439728,
-0.767991721630096,
-0.768602788448334,
-0.769214153289795,
-0.769825875759125,
-0.770437955856323,
-0.771050333976746,
-0.771663069725037,
-0.772276163101196,
-0.772889554500580,
-0.773503303527832,
-0.774117410182953,
-0.774731814861298,
-0.775346577167511,
-0.775961697101593,
-0.776577115058899,
-0.777192890644074,
-0.777809023857117,
-0.778425514698029,
-0.779042303562164,
-0.779659450054169,
-0.780276954174042,
-0.780894756317139,
-0.781512916088104,
-0.782131433486939,
-0.782750248908997,
-0.783369421958923,
-0.783988952636719,
-0.784608840942383,
-0.785229027271271,
-0.785849571228027,
-0.786470472812653,
-0.787091672420502,
-0.787713229656220,
-0.788335144519806,
-0.788957357406616,
-0.789579927921295,
-0.790202856063843,
-0.790826141834259,
-0.791449725627899,
-0.792073667049408,
-0.792697966098785,
-0.793322563171387,
-0.793947517871857,
-0.794572830200195,
-0.795198500156403,
-0.795824468135834,
-0.796450793743134,
-0.797077476978302,
-0.797704458236694,
-0.798331797122955,
-0.798959493637085,
-0.799587547779083,
-0.800215899944305,
-0.800844609737396,
-0.801473677158356,
-0.802103042602539,
-0.802732765674591,
-0.803362846374512,
-0.803993284702301,
-0.804624021053314,
-0.805255115032196,
-0.805886566638947,
-0.806518316268921,
-0.807150423526764,
-0.807782888412476,
-0.808415710926056,
-0.809048831462860,
-0.809682309627533,
-0.810316145420075,
-0.810950338840485,
-0.811584830284119,
-0.812219679355621,
-0.812854886054993,
-0.813490390777588,
-0.814126253128052,
-0.814762473106384,
-0.815399050712585,
-0.816035926342011,
-0.816673159599304,
-0.817310750484467,
-0.817948698997498,
-0.818586945533752,
-0.819225549697876,
-0.819864511489868,
-0.820503830909729,
-0.821143448352814,
-0.821783423423767,
-0.822423756122589,
-0.823064446449280,
-0.823705434799194,
-0.824346780776978,
-0.824988484382629,
-0.825630486011505,
-0.826272845268250,
-0.826915562152863,
-0.827558636665344,
-0.828202009201050,
-0.828845739364624,
-0.829489827156067,
-0.830134272575378,
-0.830779016017914,
-0.831424117088318,
-0.832069575786591,
-0.832715392112732,
-0.833361506462097,
-0.834007978439331,
-0.834654808044434,
-0.835301995277405,
-0.835949480533600,
-0.836597323417664,
-0.837245523929596,
-0.837894082069397,
-0.838542938232422,
-0.839192152023315,
-0.839841723442078,
-0.840491652488709,
-0.841141939163208,
-0.841792523860931,
-0.842443466186523,
-0.843094766139984,
-0.843746423721314,
-0.844398379325867,
-0.845050692558289,
-0.845703363418579,
-0.846356391906738,
-0.847009718418121,
-0.847663402557373,
-0.848317444324493,
-0.848971843719482,
-0.849626541137695,
-0.850281596183777,
-0.850937008857727,
-0.851592779159546,
-0.852248907089233,
-0.852905333042145,
-0.853562116622925,
-0.854219257831574,
-0.854876756668091,
-0.855534553527832,
-0.856192708015442,
-0.856851220130920,
-0.857510089874268,
-0.858169257640839,
-0.858828783035278,
-0.859488666057587,
-0.860148906707764,
-0.860809504985809,
-0.861470401287079,
-0.862131655216217,
-0.862793266773224,
-0.863455235958099,
-0.864117562770844,
-0.864780187606812,
-0.865443170070648,
-0.866106510162354,
-0.866770207881928,
-0.867434203624725,
-0.868098556995392,
-0.868763267993927,
-0.869428336620331,
-0.870093762874603,
-0.870759487152100,
-0.871425569057465,
-0.872092008590698,
-0.872758805751801,
-0.873425960540772,
-0.874093413352966,
-0.874761223793030,
-0.875429391860962,
-0.876097917556763,
-0.876766741275787,
-0.877435922622681,
-0.878105461597443,
-0.878775358200073,
-0.879445612430573,
-0.880116164684296,
-0.880787074565888,
-0.881458342075348,
-0.882129967212677,
-0.882801949977875,
-0.883474230766296,
-0.884146869182587,
-0.884819865226746,
-0.885493218898773,
-0.886166930198669,
-0.886840939521790,
-0.887515306472778,
-0.888190031051636,
-0.888865113258362,
-0.889540553092957,
-0.890216290950775,
-0.890892386436462,
-0.891568839550018,
-0.892245650291443,
-0.892922818660736,
-0.893600344657898,
-0.894278168678284,
-0.894956350326538,
-0.895634889602661,
-0.896313786506653,
-0.896993041038513,
-0.897672593593597,
-0.898352503776550,
-0.899032771587372,
-0.899713397026062,
-0.900394380092621,
-0.901075720787048,
-0.901757359504700,
-0.902439355850220,
-0.903121709823608,
-0.903804421424866,
-0.904487490653992,
-0.905170857906342,
-0.905854582786560,
-0.906538665294647,
-0.907223105430603,
-0.907907903194428,
-0.908593058586121,
-0.909278512001038,
-0.909964323043823,
-0.910650491714478,
-0.911337018013001,
-0.912023901939392,
-0.912711143493652,
-0.913398683071137,
-0.914086580276489,
-0.914774835109711,
-0.915463447570801,
-0.916152417659760,
-0.916841745376587,
-0.917531371116638,
-0.918221354484558,
-0.918911695480347,
-0.919602394104004,
-0.920293450355530,
-0.920984864234924,
-0.921676576137543,
-0.922368645668030,
-0.923061072826386,
-0.923753857612610,
-0.924447000026703,
-0.925140500068665,
-0.925834298133850,
-0.926528453826904,
-0.927222967147827,
-0.927917838096619,
-0.928613066673279,
-0.929308652877808,
-0.930004596710205,
-0.930700838565826,
-0.931397438049316,
-0.932094395160675,
-0.932791709899902,
-0.933489382266998,
-0.934187412261963,
-0.934885799884796,
-0.935584485530853,
-0.936283528804779,
-0.936982929706574,
-0.937682688236237,
-0.938382804393768,
-0.939083278179169,
-0.939784109592438,
-0.940485239028931,
-0.941186726093292,
-0.941888570785523,
-0.942590773105621,
-0.943293333053589,
-0.943996250629425,
-0.944699525833130,
-0.945403099060059,
-0.946107029914856,
-0.946811318397522,
-0.947515964508057,
-0.948220968246460,
-0.948926329612732,
-0.949632048606873,
-0.950338065624237,
-0.951044440269470,
-0.951751172542572,
-0.952458262443543,
-0.953165709972382,
-0.953873515129089,
-0.954581677913666,
-0.955290198326111,
-0.955999016761780,
-0.956708192825317,
-0.957417726516724,
-0.958127617835999,
-0.958837866783142,
-0.959548473358154,
-0.960259437561035,
-0.960970759391785,
-0.961682379245758,
-0.962394356727600,
-0.963106691837311,
-0.963819384574890,
-0.964532434940338,
-0.965245842933655,
-0.965959608554840,
-0.966673731803894,
-0.967388153076172,
-0.968102931976318,
-0.968818068504334,
-0.969533562660217,
-0.970249414443970,
-0.970965623855591,
-0.971682190895081,
-0.972399115562439,
-0.973116397857666,
-0.973833978176117,
-0.974551916122437,
-0.975270211696625,
-0.975988864898682,
-0.976707875728607,
-0.977427244186401,
-0.978146970272064,
-0.978867053985596,
-0.979587495326996,
-0.980308234691620,
-0.981029331684113,
-0.981750786304474,
-0.982472598552704,
-0.983194768428803,
-0.983917295932770,
-0.984640181064606,
-0.985363423824310,
-0.986087024211884,
-0.986810922622681,
-0.987535178661346,
-0.988259792327881,
-0.988984763622284,
-0.989710092544556,
-0.990435779094696,
-0.991161823272705,
-0.991888225078583,
-0.992614984512329,
-0.993342101573944,
-0.994069576263428,
-0.994797348976135,
-0.995525479316711,
-0.996253967285156,
-0.996982812881470,
-0.997712016105652,
-0.998441576957703,
-0.999171495437622,
-0.999901771545410,
-1.00063240528107,
-1.00136339664459,
-1.00209474563599,
-1.00282645225525,
-1.00355851650238,
-1.00429093837738,
-1.00502371788025,
-1.00575685501099,
-1.00649023056030,
-1.00722396373749,
-1.00795805454254,
-1.00869250297546,
-1.00942730903625,
-1.01016247272491,
-1.01089799404144,
-1.01163387298584,
-1.01237010955811,
-1.01310670375824,
-1.01384365558624,
-1.01458096504211,
-1.01531863212585,
-1.01605665683746,
-1.01679503917694,
-1.01753377914429,
-1.01827287673950,
-1.01901233196259,
-1.01975214481354,
-1.02049231529236,
-1.02123284339905,
-1.02197372913361,
-1.02271497249603,
-1.02345657348633,
-1.02419853210449,
-1.02494072914124,
-1.02568328380585,
-1.02642619609833,
-1.02716946601868,
-1.02791309356689,
-1.02865707874298,
-1.02940142154694,
-1.03014612197876,
-1.03089118003845,
-1.03163659572601,
-1.03238236904144,
-1.03312849998474,
-1.03387498855591,
-1.03462183475494,
-1.03536903858185,
-1.03611660003662,
-1.03686451911926,
-1.03761279582977,
-1.03836143016815,
-1.03911042213440,
-1.03985977172852,
-1.04060947895050,
-1.04135954380035,
-1.04210996627808,
-1.04286074638367,
-1.04361188411713,
-1.04436337947845,
-1.04511523246765,
-1.04586744308472,
-1.04662001132965,
-1.04737293720245,
-1.04812610149384,
-1.04887962341309,
-1.04963350296021,
-1.05038774013519,
-1.05114233493805,
-1.05189728736877,
-1.05265259742737,
-1.05340826511383,
-1.05416429042816,
-1.05492067337036,
-1.05567741394043,
-1.05643451213837,
-1.05719196796417,
-1.05794978141785,
-1.05870795249939,
-1.05946648120880,
-1.06022536754608,
-1.06098461151123,
-1.06174421310425,
-1.06250417232513,
-1.06326448917389,
-1.06402516365051,
-1.06478619575500,
-1.06554758548737,
-1.06630933284760,
-1.06707143783569,
-1.06783390045166,
-1.06859672069550,
-1.06935989856720,
-1.07012343406677,
-1.07088732719421,
-1.07165157794952,
-1.07241618633270,
-1.07318115234375,
-1.07394647598267,
-1.07471215724945,
-1.07547819614410,
-1.07624459266663,
-1.07701134681702,
-1.07777845859528,
-1.07854580879211,
-1.07931351661682,
-1.08008158206940,
-1.08085000514984,
-1.08161878585815,
-1.08238792419434,
-1.08315742015839,
-1.08392727375031,
-1.08469748497009,
-1.08546805381775,
-1.08623898029327,
-1.08701026439667,
-1.08778190612793,
-1.08855390548706,
-1.08932626247406,
-1.09009897708893,
-1.09087204933167,
-1.09164547920227,
-1.09241926670074,
-1.09319341182709,
-1.09396791458130,
-1.09474277496338,
-1.09551799297333,
-1.09629356861115,
-1.09706950187683,
-1.09784579277039,
-1.09862244129181,
-1.09939944744110,
-1.10017681121826,
-1.10095453262329,
-1.10173261165619,
-1.10251104831696,
-1.10328984260559,
-1.10406899452209,
-1.10484850406647,
-1.10562837123871,
-1.10640859603882,
-1.10718917846680,
-1.10797011852264,
-1.10875141620636,
-1.10953307151794,
-1.11031508445740,
-1.11109745502472,
-1.11188018321991,
-1.11266326904297,
-1.11344671249390,
-1.11423051357269,
-1.11501467227936,
-1.11579918861389,
-1.11658406257629,
-1.11736929416657,
-1.11815488338470,
-1.11894083023071,
-1.11972713470459,
-1.12051379680634,
-1.12130081653595,
-1.12208819389343,
-1.12287592887878,
-1.12366390228271,
-1.12445223331451,
-1.12524092197418,
-1.12602996826172,
-1.12681937217712,
-1.12760913372040,
-1.12839925289154,
-1.12918972969055,
-1.12998056411743,
-1.13077175617218,
-1.13156330585480,
-1.13235521316528,
-1.13314747810364,
-1.13394010066986,
-1.13473308086395,
-1.13552641868591,
-1.13632011413574,
-1.13711416721344,
-1.13790857791901,
-1.13870334625244,
-1.13949847221375,
-1.14029395580292,
-1.14108979701996,
-1.14188599586487,
-1.14268255233765,
-1.14347946643829,
-1.14427673816681,
-1.14507436752319,
-1.14587235450745,
-1.14667069911957,
-1.14746940135956,
-1.14826846122742,
-1.14906787872314,
-1.14986765384674,
-1.15066778659821,
-1.15146827697754,
-1.15226912498474,
-1.15307033061981,
-1.15387189388275,
-1.15467381477356,
-1.15547609329224,
-1.15627872943878,
-1.15708172321320,
-1.15788507461548,
-1.15868878364563,
-1.15949285030365,
-1.16029727458954,
-1.16110205650330,
-1.16190719604492,
-1.16271269321442,
-1.16351854801178,
-1.16432476043701,
-1.16513133049011,
-1.16593825817108,
-1.16674554347992,
-1.16755318641663,
-1.16836118698120,
-1.16916954517365,
-1.16997826099396,
-1.17078733444214,
-1.17159676551819,
-1.17240655422211,
-1.17321670055389,
-1.17402720451355,
-1.17483806610107,
-1.17564928531647,
-1.17646086215973,
-1.17727279663086,
-1.17808508872986,
-1.17889773845673,
-1.17971074581146,
-1.18052411079407,
-1.18133783340454,
-1.18215191364288,
-1.18296635150909,
-1.18378114700317,
-1.18459630012512,
-1.18541181087494,
-1.18622767925262,
-1.18704390525818,
-1.18786048889160,
-1.18867743015289,
-1.18949472904205,
-1.19031238555908,
-1.19113039970398,
-1.19194877147675,
-1.19276750087738,
-1.19358658790588,
-1.19440603256226,
-1.19522583484650,
-1.19604599475861,
-1.19686651229858,
-1.19768738746643,
-1.19850862026215,
-1.19933021068573,
-1.20015215873718,
-1.20097446441650,
-1.20179712772369,
-1.20262014865875,
-1.20344352722168,
-1.20426726341248,
-1.20509135723114,
-1.20591580867767,
-1.20674061775208,
-1.20756578445435,
-1.20839130878448,
-1.20921719074249,
-1.21004343032837,
-1.21087002754211,
-1.21169698238373,
-1.21252429485321,
-1.21335196495056,
-1.21417999267578,
-1.21500837802887,
-1.21583712100983,
-1.21666622161865,
-1.21749567985535,
-1.21832549571991,
-1.21915566921234,
-1.21998620033264,
-1.22081708908081,
-1.22164833545685,
-1.22247993946075,
-1.22331190109253,
-1.22414422035217,
-1.22497689723969,
-1.22580993175507,
-1.22664332389832,
-1.22747707366943,
-1.22831118106842,
-1.22914564609528,
-1.22998046875000,
-1.23081564903259,
-1.23165118694305,
-1.23248708248138,
-1.23332333564758,
-1.23415994644165,
-1.23499691486359,
-1.23583424091339,
-1.23667192459106,
-1.23750996589661,
-1.23834836483002,
-1.23918712139130,
-1.24002623558044,
-1.24086558818817,
-1.24170529842377,
-1.24254536628723,
-1.24338579177856,
-1.24422657489777,
-1.24506771564484,
-1.24590921401978,
-1.24675107002258,
-1.24759328365326,
-1.24843585491180,
-1.24927878379822,
-1.25012207031250,
-1.25096571445465,
-1.25180971622467,
-1.25265407562256,
-1.25349879264832,
-1.25434386730194,
-1.25518929958344,
-1.25603508949280,
-1.25688123703003,
-1.25772774219513,
-1.25857460498810,
-1.25942182540894,
-1.26026940345764,
-1.26111733913422,
-1.26196563243866,
-1.26281428337097,
-1.26366329193115,
-1.26451265811920,
-1.26536238193512,
-1.26621246337891,
-1.26706290245056,
-1.26791369915009,
-1.26876485347748,
-1.26961636543274,
-1.27046823501587,
-1.27132046222687,
-1.27217304706573,
-1.27302598953247,
-1.27387928962708,
-1.27473294734955,
-1.27558696269989,
-1.27644133567810,
-1.27729606628418,
-1.27815115451813,
-1.27900660037994,
-1.27986240386963,
-1.28071856498718,
-1.28157508373261,
-1.28243196010590,
-1.28328919410706,
-1.28414678573608,
-1.28500473499298,
-1.28586304187775,
-1.28672170639038,
-1.28758072853088,
-1.28844010829926,
-1.28929984569550,
-1.29015994071960,
-1.29102039337158,
-1.29188120365143,
-1.29274237155914,
-1.29360389709473,
-1.29446578025818,
-1.29532802104950,
-1.29619061946869,
-1.29705357551575,
-1.29791688919067,
-1.29878056049347,
-1.29964458942413,
-1.30050897598267,
-1.30137372016907,
-1.30223882198334,
-1.30310428142548,
-1.30397009849548,
-1.30483627319336,
-1.30570280551910,
-1.30656969547272,
-1.30743694305420,
-1.30830454826355,
-1.30917251110077,
-1.31004083156586,
-1.31090950965881,
-1.31177854537964,
-1.31264793872833,
-1.31351768970490,
-1.31438779830933,
-1.31525826454163,
-1.31612908840179,
-1.31700026988983,
-1.31787180900574,
-1.31874370574951,
-1.31961596012115,
-1.32048857212067,
-1.32136154174805,
-1.32223486900330,
-1.32310855388641,
-1.32398259639740,
-1.32485699653625,
-1.32573175430298,
-1.32660686969757,
-1.32748234272003,
-1.32835817337036,
-1.32923436164856,
-1.33011090755463,
-1.33098781108856,
-1.33186507225037,
-1.33274269104004,
-1.33362066745758,
-1.33449900150299,
-1.33537769317627,
-1.33625674247742,
-1.33713614940643,
-1.33801591396332,
-1.33889603614807,
-1.33977651596069,
-1.34065735340118,
-1.34153854846954,
-1.34242010116577,
-1.34330201148987,
-1.34418427944183,
-1.34506690502167,
-1.34594988822937,
-1.34683322906494,
-1.34771692752838,
-1.34860098361969,
-1.34948539733887,
-1.35037016868591,
-1.35125529766083,
-1.35214078426361,
-1.35302662849426,
-1.35391283035278,
-1.35479938983917,
-1.35568630695343,
-1.35657358169556,
-1.35746121406555,
-1.35834920406342,
-1.35923755168915,
-1.36012625694275,
-1.36101531982422,
-1.36190474033356,
-1.36279451847076,
-1.36368465423584,
-1.36457514762878,
-1.36546599864960,
-1.36635720729828,
-1.36724877357483,
-1.36814069747925,
-1.36903297901154,
-1.36992561817169,
-1.37081861495972,
-1.37171196937561,
-1.37260568141937,
-1.37349975109100,
-1.37439417839050,
-1.37528896331787,
-1.37618410587311,
-1.37707960605621,
-1.37797546386719,
-1.37887167930603,
-1.37976825237274,
-1.38066518306732,
-1.38156247138977,
-1.38246011734009,
-1.38335812091827,
-1.38425648212433,
-1.38515520095825,
-1.38605427742004,
-1.38695371150970,
-1.38785350322723,
-1.38875365257263,
-1.38965415954590,
-1.39055502414703,
-1.39145624637604,
-1.39235782623291,
-1.39325976371765,
-1.39416205883026,
-1.39506471157074,
-1.39596772193909,
-1.39687108993530,
-1.39777481555939,
-1.39867889881134,
-1.39958333969116,
-1.40048813819885,
-1.40139329433441,
-1.40229880809784,
-1.40320467948914,
-1.40411090850830,
-1.40501749515533,
-1.40592443943024,
-1.40683174133301,
-1.40773940086365,
-1.40864741802216,
-1.40955579280853,
-1.41046452522278,
-1.41137361526489,
-1.41228306293488,
-1.41319286823273,
-1.41410303115845,
-1.41501355171204,
-1.41592442989349,
-1.41683566570282,
-1.41774725914001,
-1.41865921020508,
-1.41957151889801,
-1.42048418521881,
-1.42139720916748,
-1.42231059074402,
-1.42322432994843,
-1.42413842678070,
-1.42505288124084,
-1.42596769332886,
-1.42688286304474,
-1.42779839038849,
-1.42871427536011,
-1.42963051795959,
-1.43054711818695,
-1.43146407604218,
-1.43238139152527,
-1.43329906463623,
-1.43421709537506,
-1.43513548374176,
-1.43605422973633,
-1.43697333335876,
-1.43789279460907,
-1.43881261348724,
-1.43973278999329,
-1.44065332412720,
-1.44157421588898,
-1.44249546527863,
-1.44341707229614,
-1.44433903694153,
-1.44526135921478,
-1.44618403911591,
-1.44710707664490,
-1.44803047180176,
-1.44895422458649,
-1.44987833499908,
-1.45080280303955,
-1.45172762870789,
-1.45265281200409,
-1.45357835292816,
-1.45450425148010,
-1.45543050765991,
-1.45635712146759,
-1.45728409290314,
-1.45821142196655,
-1.45913910865784,
-1.46006715297699,
-1.46099555492401,
-1.46192431449890,
-1.46285343170166,
-1.46378290653229,
-1.46471273899078,
-1.46564292907715,
-1.46657347679138,
-1.46750438213348,
-1.46843564510345,
-1.46936726570129,
-1.47029924392700,
-1.47123157978058,
-1.47216427326202,
-1.47309732437134,
-1.47403073310852,
-1.47496449947357,
-1.47589862346649,
-1.47683310508728,
-1.47776794433594,
-1.47870314121246,
-1.47963869571686,
-1.48057460784912,
-1.48151087760925,
-1.48244750499725,
-1.48338449001312,
-1.48432183265686,
-1.48525953292847,
-1.48619759082794,
-1.48713600635529,
-1.48807477951050,
-1.48901391029358,
-1.48995339870453,
-1.49089324474335,
-1.49183344841003,
-1.49277400970459,
-1.49371492862701,
-1.49465620517731,
-1.49559783935547,
-1.49653983116150,
-1.49748206138611,
-1.49842464923859,
-1.49936759471893,
-1.50031089782715,
-1.50125455856323,
-1.50219857692719,
-1.50314295291901,
-1.50408768653870,
-1.50503277778625,
-1.50597822666168,
-1.50692403316498,
-1.50787019729614,
-1.50881671905518,
-1.50976359844208,
-1.51071083545685,
-1.51165843009949,
-1.51260638237000,
-1.51355469226837,
-1.51450335979462,
-1.51545238494873,
-1.51640176773071,
-1.51735150814056,
-1.51830160617828,
-1.51925206184387,
-1.52020287513733,
-1.52115404605865,
-1.52210557460785,
-1.52305746078491,
-1.52400970458984,
-1.52496230602264,
-1.52591526508331,
-1.52686858177185,
-1.52782225608826,
-1.52877628803253,
-1.52973067760468,
-1.53068542480469,
-1.53164052963257,
-1.53259599208832,
-1.53355181217194,
-1.53450798988342,
-1.53546452522278,
-1.53642141819000,
-1.53737866878510,
-1.53833627700806,
-1.53929424285889,
-1.54025256633759,
-1.54121124744415,
-1.54217028617859,
-1.54312968254089,
-1.54408943653107,
-1.54504954814911,
-1.54601001739502,
-1.54697084426880,
-1.54793202877045,
-1.54889357089996,
-1.54985535144806,
-1.55081748962402,
-1.55177998542786,
-1.55274283885956,
-1.55370604991913,
-1.55466961860657,
-1.55563354492188,
-1.55659782886505,
-1.55756247043610,
-1.55852746963501,
-1.55949282646179,
-1.56045854091644,
-1.56142461299896,
-1.56239104270935,
-1.56335783004761,
-1.56432497501373,
-1.56529247760773,
-1.56626033782959,
-1.56722855567932,
-1.56819713115692,
-1.56916606426239,
-1.57013535499573,
-1.57110500335693,
-1.57207500934601,
-1.57304537296295,
-1.57401609420776,
-1.57498717308044,
-1.57595860958099,
-1.57693040370941,
-1.57790255546570,
-1.57887506484985,
-1.57984793186188,
-1.58082115650177,
-1.58179473876953,
-1.58276867866516,
-1.58374297618866,
-1.58471751213074,
-1.58569240570068,
-1.58666765689850,
-1.58764326572418,
-1.58861923217773,
-1.58959555625916,
-1.59057223796844,
-1.59154927730560,
-1.59252667427063,
-1.59350442886353,
-1.59448254108429,
-1.59546101093292,
-1.59643983840942,
-1.59741902351379,
-1.59839856624603,
-1.59937846660614,
-1.60035872459412,
-1.60133934020996,
-1.60232031345367,
-1.60330164432526,
-1.60428333282471,
-1.60526537895203,
-1.60624778270721,
-1.60723054409027,
-1.60821366310120,
-1.60919713973999,
-1.61018097400665,
-1.61116516590118,
-1.61214971542358,
-1.61313450336456,
-1.61411964893341,
-1.61510515213013,
-1.61609101295471,
-1.61707723140717,
-1.61806380748749,
-1.61905074119568,
-1.62003803253174,
-1.62102568149567,
-1.62201368808746,
-1.62300205230713,
-1.62399077415466,
-1.62497985363007,
-1.62596929073334,
-1.62695908546448,
-1.62794923782349,
-1.62893974781036,
-1.62993061542511,
-1.63092184066772,
-1.63191342353821,
-1.63290536403656,
-1.63389766216278,
-1.63489031791687,
-1.63588321208954,
-1.63687646389008,
-1.63787007331848,
-1.63886404037476,
-1.63985836505890,
-1.64085304737091,
-1.64184808731079,
-1.64284348487854,
-1.64383924007416,
-1.64483535289764,
-1.64583182334900,
-1.64682865142822,
-1.64782583713532,
-1.64882338047028,
-1.64982128143311,
-1.65081954002380,
-1.65181815624237,
-1.65281713008881,
-1.65381646156311,
-1.65481615066528,
-1.65581607818604,
-1.65681636333466,
-1.65781700611115,
-1.65881800651550,
-1.65981936454773,
-1.66082108020782,
-1.66182315349579,
-1.66282558441162,
-1.66382837295532,
-1.66483151912689,
-1.66583502292633,
-1.66683888435364,
-1.66784310340881,
-1.66884768009186,
-1.66985261440277,
-1.67085790634155,
-1.67186355590820,
-1.67286956310272,
-1.67387580871582,
-1.67488241195679,
-1.67588937282562,
-1.67689669132233,
-1.67790436744690,
-1.67891240119934,
-1.67992079257965,
-1.68092954158783,
-1.68193864822388,
-1.68294811248779,
-1.68395793437958,
-1.68496811389923,
-1.68597865104675,
-1.68698954582214,
-1.68800079822540,
-1.68901240825653,
-1.69002425670624,
-1.69103646278381,
-1.69204902648926,
-1.69306194782257,
-1.69407522678375,
-1.69508886337280,
-1.69610285758972,
-1.69711720943451,
-1.69813191890717,
-1.69914698600769,
-1.70016241073608,
-1.70117819309235,
-1.70219433307648,
-1.70321083068848,
-1.70422768592834,
-1.70524477958679,
-1.70626223087311,
-1.70728003978729,
-1.70829820632935,
-1.70931673049927,
-1.71033561229706,
-1.71135485172272,
-1.71237444877625,
-1.71339440345764,
-1.71441471576691,
-1.71543538570404,
-1.71645641326904,
-1.71747779846191,
-1.71849942207336,
-1.71952140331268,
-1.72054374217987,
-1.72156643867493,
-1.72258949279785,
-1.72361290454865,
-1.72463667392731,
-1.72566080093384,
-1.72668528556824,
-1.72771012783051,
-1.72873532772064,
-1.72976088523865,
-1.73078680038452,
-1.73181295394897,
-1.73283946514130,
-1.73386633396149,
-1.73489356040955,
-1.73592114448547,
-1.73694908618927,
-1.73797738552094,
-1.73900604248047,
-1.74003505706787,
-1.74106442928314,
-1.74209415912628,
-1.74312424659729,
-1.74415457248688,
-1.74518525600433,
-1.74621629714966,
-1.74724769592285,
-1.74827945232391,
-1.74931156635284,
-1.75034403800964,
-1.75137686729431,
-1.75241005420685,
-1.75344359874725,
-1.75447750091553,
-1.75551164150238,
-1.75654613971710,
-1.75758099555969,
-1.75861620903015,
-1.75965178012848,
-1.76068770885468,
-1.76172399520874,
-1.76276063919067,
-1.76379764080048,
-1.76483500003815,
-1.76587259769440,
-1.76691055297852,
-1.76794886589050,
-1.76898753643036,
-1.77002656459808,
-1.77106595039368,
-1.77210569381714,
-1.77314579486847,
-1.77418625354767,
-1.77522706985474,
-1.77626812458038,
-1.77730953693390,
-1.77835130691528,
-1.77939343452454,
-1.78043591976166,
-1.78147876262665,
-1.78252196311951,
-1.78356552124023,
-1.78460943698883,
-1.78565371036530,
-1.78669822216034,
-1.78774309158325,
-1.78878831863403,
-1.78983390331268,
-1.79087984561920,
-1.79192614555359,
-1.79297280311584,
-1.79401981830597,
-1.79506719112396,
-1.79611480236053,
-1.79716277122498,
-1.79821109771729,
-1.79925978183746,
-1.80030882358551,
-1.80135822296143,
-1.80240797996521,
-1.80345809459686,
-1.80450856685638,
-1.80555927753448,
-1.80661034584045,
-1.80766177177429,
-1.80871355533600,
-1.80976569652557,
-1.81081819534302,
-1.81187105178833,
-1.81292426586151,
-1.81397783756256,
-1.81503164768219,
-1.81608581542969,
-1.81714034080505,
-1.81819522380829,
-1.81925046443939,
-1.82030606269836,
-1.82136201858521,
-1.82241833209991,
-1.82347488403320,
-1.82453179359436,
-1.82558906078339,
-1.82664668560028,
-1.82770466804504,
-1.82876300811768,
-1.82982170581818,
-1.83088076114655,
-1.83194005489349,
-1.83299970626831,
-1.83405971527100,
-1.83512008190155,
-1.83618080615997,
-1.83724188804626,
-1.83830332756042,
-1.83936500549316,
-1.84042704105377,
-1.84148943424225,
-1.84255218505859,
-1.84361529350281,
-1.84467875957489,
-1.84574258327484,
-1.84680676460266,
-1.84787118434906,
-1.84893596172333,
-1.85000109672546,
-1.85106658935547,
-1.85213243961334,
-1.85319864749908,
-1.85426521301270,
-1.85533201694489,
-1.85639917850494,
-1.85746669769287,
-1.85853457450867,
-1.85960280895233,
-1.86067140102386,
-1.86174035072327,
-1.86280965805054,
-1.86387920379639,
-1.86494910717011,
-1.86601936817169,
-1.86708998680115,
-1.86816096305847,
-1.86923229694366,
-1.87030398845673,
-1.87137591838837,
-1.87244820594788,
-1.87352085113525,
-1.87459385395050,
-1.87566721439362,
-1.87674093246460,
-1.87781488895416,
-1.87888920307159,
-1.87996387481689,
-1.88103890419006,
-1.88211429119110,
-1.88319003582001,
-1.88426613807678,
-1.88534247875214,
-1.88641917705536,
-1.88749623298645,
-1.88857364654541,
-1.88965141773224,
-1.89072954654694,
-1.89180803298950,
-1.89288675785065,
-1.89396584033966,
-1.89504528045654,
-1.89612507820129,
-1.89720523357391,
-1.89828574657440,
-1.89936649799347,
-1.90044760704041,
-1.90152907371521,
-1.90261089801788,
-1.90369307994843,
-1.90477561950684,
-1.90585851669312,
-1.90694165229797,
-1.90802514553070,
-1.90910899639130,
-1.91019320487976,
-1.91127777099609,
-1.91236269474030,
-1.91344785690308,
-1.91453337669373,
-1.91561925411224,
-1.91670548915863,
-1.91779208183289,
-1.91887903213501,
-1.91996622085571,
-1.92105376720428,
-1.92214167118073,
-1.92322993278503,
-1.92431855201721,
-1.92540752887726,
-1.92649674415588,
-1.92758631706238,
-1.92867624759674,
-1.92976653575897,
-1.93085718154907,
-1.93194818496704,
-1.93303942680359,
-1.93413102626801,
-1.93522298336029,
-1.93631529808044,
-1.93740797042847,
-1.93850100040436,
-1.93959426879883,
-1.94068789482117,
-1.94178187847137,
-1.94287621974945,
-1.94397091865540,
-1.94506585597992,
-1.94616115093231,
-1.94725680351257,
-1.94835281372070,
-1.94944918155670,
-1.95054590702057,
-1.95164287090302,
-1.95274019241333,
-1.95383787155151,
-1.95493590831757,
-1.95603430271149,
-1.95713293552399,
-1.95823192596436,
-1.95933127403259,
-1.96043097972870,
-1.96153104305267,
-1.96263146400452,
-1.96373212337494,
-1.96483314037323,
-1.96593451499939,
-1.96703624725342,
-1.96813833713532,
-1.96924066543579,
-1.97034335136414,
-1.97144639492035,
-1.97254979610443,
-1.97365355491638,
-1.97475767135620,
-1.97586202621460,
-1.97696673870087,
-1.97807180881500,
-1.97917723655701,
-1.98028302192688,
-1.98138904571533,
-1.98249542713165,
-1.98360216617584,
-1.98470926284790,
-1.98581671714783,
-1.98692440986633,
-1.98803246021271,
-1.98914086818695,
-1.99024963378906,
-1.99135875701904,
-1.99246811866760,
-1.99357783794403,
-1.99468791484833,
-1.99579834938049,
-1.99690914154053,
-1.99802017211914,
-1.99913156032562,
-2.00024318695068,
-2.00135517120361,
-2.00246763229370,
-2.00358033180237,
-2.00469350814819,
-2.00580692291260,
-2.00692057609558,
-2.00803470611572,
-2.00914907455444,
-2.01026391983032,
-2.01137900352478,
-2.01249432563782,
-2.01361012458801,
-2.01472616195679,
-2.01584267616272,
-2.01695942878723,
-2.01807641983032,
-2.01919388771057,
-2.02031159400940,
-2.02142977714539,
-2.02254819869995,
-2.02366685867310,
-2.02478599548340,
-2.02590537071228,
-2.02702498435974,
-2.02814507484436,
-2.02926540374756,
-2.03038620948792,
-2.03150725364685,
-2.03262853622437,
-2.03375029563904,
-2.03487229347229,
-2.03599476814270,
-2.03711748123169,
-2.03824043273926,
-2.03936386108398,
-2.04048752784729,
-2.04161167144775,
-2.04273605346680,
-2.04386067390442,
-2.04498577117920,
-2.04611110687256,
-2.04723668098450,
-2.04836273193359,
-2.04948902130127,
-2.05061578750610,
-2.05174279212952,
-2.05287003517151,
-2.05399775505066,
-2.05512571334839,
-2.05625414848328,
-2.05738282203674,
-2.05851173400879,
-2.05964112281799,
-2.06077075004578,
-2.06190061569214,
-2.06303095817566,
-2.06416153907776,
-2.06529259681702,
-2.06642389297485,
-2.06755542755127,
-2.06868743896484,
-2.06981968879700,
-2.07095217704773,
-2.07208514213562,
-2.07321834564209,
-2.07435202598572,
-2.07548594474793,
-2.07662010192871,
-2.07775473594666,
-2.07888960838318,
-2.08002495765686,
-2.08116054534912,
-2.08229637145996,
-2.08343267440796,
-2.08456921577454,
-2.08570599555969,
-2.08684325218201,
-2.08798074722290,
-2.08911871910095,
-2.09025692939758,
-2.09139537811279,
-2.09253430366516,
-2.09367346763611,
-2.09481287002563,
-2.09595274925232,
-2.09709286689758,
-2.09823322296143,
-2.09937405586243,
-2.10051512718201,
-2.10165667533875,
-2.10279846191406,
-2.10394048690796,
-2.10508298873901,
-2.10622572898865,
-2.10736870765686,
-2.10851216316223,
-2.10965585708618,
-2.11080002784729,
-2.11194443702698,
-2.11308908462524,
-2.11423420906067,
-2.11537957191467,
-2.11652517318726,
-2.11767125129700,
-2.11881756782532,
-2.11996412277222,
-2.12111115455627,
-2.12225842475891,
-2.12340617179871,
-2.12455415725708,
-2.12570238113403,
-2.12685108184814,
-2.12800002098084,
-2.12914919853210,
-2.13029885292053,
-2.13144874572754,
-2.13259887695313,
-2.13374948501587,
-2.13490033149719,
-2.13605165481567,
-2.13720321655273,
-2.13835501670837,
-2.13950729370117,
-2.14065980911255,
-2.14181256294251,
-2.14296579360962,
-2.14411926269531,
-2.14527297019959,
-2.14642715454102,
-2.14758157730103,
-2.14873647689819,
-2.14989161491394,
-2.15104699134827,
-2.15220284461975,
-2.15335893630981,
-2.15451526641846,
-2.15567207336426,
-2.15682911872864,
-2.15798640251160,
-2.15914416313171,
-2.16030216217041,
-2.16146039962769,
-2.16261911392212,
-2.16377806663513,
-2.16493725776672,
-2.16609692573547,
-2.16725683212280,
-2.16841721534729,
-2.16957783699036,
-2.17073869705200,
-2.17190003395081,
-2.17306160926819,
-2.17422342300415,
-2.17538571357727,
-2.17654824256897,
-2.17771100997925,
-2.17887425422668,
-2.18003773689270,
-2.18120145797730,
-2.18236565589905,
-2.18353009223938,
-2.18469476699829,
-2.18585991859436,
-2.18702530860901,
-2.18819093704224,
-2.18935704231262,
-2.19052338600159,
-2.19168996810913,
-2.19285702705383,
-2.19402432441711,
-2.19519186019897,
-2.19635987281799,
-2.19752812385559,
-2.19869661331177,
-2.19986557960510,
-2.20103478431702,
-2.20220422744751,
-2.20337414741516,
-2.20454430580139,
-2.20571470260620,
-2.20688557624817,
-2.20805668830872,
-2.20922803878784,
-2.21039986610413,
-2.21157193183899,
-2.21274423599243,
-2.21391701698303,
-2.21509003639221,
-2.21626329421997,
-2.21743702888489,
-2.21861100196838,
-2.21978521347046,
-2.22095990180969,
-2.22213482856751,
-2.22330999374390,
-2.22448563575745,
-2.22566151618958,
-2.22683763504028,
-2.22801423072815,
-2.22919106483459,
-2.23036813735962,
-2.23154568672180,
-2.23272347450256,
-2.23390150070190,
-2.23508000373840,
-2.23625874519348,
-2.23743772506714,
-2.23861718177795,
-2.23979687690735,
-2.24097681045532,
-2.24215722084045,
-2.24333786964417,
-2.24451875686646,
-2.24570012092590,
-2.24688172340393,
-2.24806356430054,
-2.24924588203430,
-2.25042843818665,
-2.25161123275757,
-2.25279450416565,
-2.25397801399231,
-2.25516176223755,
-2.25634598731995,
-2.25753045082092,
-2.25871515274048,
-2.25990033149719,
-2.26108574867249,
-2.26227140426636,
-2.26345753669739,
-2.26464390754700,
-2.26583051681519,
-2.26701736450195,
-2.26820468902588,
-2.26939225196838,
-2.27058005332947,
-2.27176833152771,
-2.27295684814453,
-2.27414560317993,
-2.27533483505249,
-2.27652430534363,
-2.27771401405334,
-2.27890419960022,
-2.28009462356567,
-2.28128528594971,
-2.28247642517090,
-2.28366780281067,
-2.28485941886902,
-2.28605127334595,
-2.28724360466003,
-2.28843617439270,
-2.28962898254395,
-2.29082226753235,
-2.29201579093933,
-2.29320955276489,
-2.29440379142761,
-2.29559826850891,
-2.29679298400879,
-2.29798817634583,
-2.29918360710144,
-2.30037927627563,
-2.30157518386841,
-2.30277156829834,
-2.30396819114685,
-2.30516505241394,
-2.30636239051819,
-2.30755996704102,
-2.30875778198242,
-2.30995607376099,
-2.31115460395813,
-2.31235337257385,
-2.31355237960815,
-2.31475186347961,
-2.31595158576965,
-2.31715154647827,
-2.31835198402405,
-2.31955265998840,
-2.32075357437134,
-2.32195496559143,
-2.32315659523010,
-2.32435846328735,
-2.32556056976318,
-2.32676315307617,
-2.32796597480774,
-2.32916903495789,
-2.33037257194519,
-2.33157634735107,
-2.33278036117554,
-2.33398461341858,
-2.33518934249878,
-2.33639430999756,
-2.33759951591492,
-2.33880519866943,
-2.34001111984253,
-2.34121727943420,
-2.34242367744446,
-2.34363055229187,
-2.34483766555786,
-2.34604501724243,
-2.34725284576416,
-2.34846091270447,
-2.34966921806335,
-2.35087776184082,
-2.35208678245544,
-2.35329604148865,
-2.35450553894043,
-2.35571551322937,
-2.35692572593689,
-2.35813617706299,
-2.35934686660767,
-2.36055803298950,
-2.36176943778992,
-2.36298108100891,
-2.36419320106506,
-2.36540555953980,
-2.36661815643311,
-2.36783099174500,
-2.36904430389404,
-2.37025785446167,
-2.37147164344788,
-2.37268590927124,
-2.37390041351318,
-2.37511515617371,
-2.37633013725281,
-2.37754559516907,
-2.37876129150391,
-2.37997722625732,
-2.38119339942932,
-2.38241004943848,
-2.38362693786621,
-2.38484406471252,
-2.38606166839600,
-2.38727951049805,
-2.38849759101868,
-2.38971590995789,
-2.39093470573425,
-2.39215373992920,
-2.39337301254272,
-2.39459252357483,
-2.39581251144409,
-2.39703273773193,
-2.39825320243835,
-2.39947390556335,
-2.40069508552551,
-2.40191650390625,
-2.40313816070557,
-2.40436029434204,
-2.40558266639709,
-2.40680527687073,
-2.40802812576294,
-2.40925145149231,
-2.41047501564026,
-2.41169881820679,
-2.41292285919189,
-2.41414737701416,
-2.41537213325501,
-2.41659712791443,
-2.41782236099243,
-2.41904807090759,
-2.42027401924133,
-2.42150020599365,
-2.42272663116455,
-2.42395353317261,
-2.42518067359924,
-2.42640805244446,
-2.42763566970825,
-2.42886376380920,
-2.43009209632874,
-2.43132066726685,
-2.43254947662354,
-2.43377876281738,
-2.43500828742981,
-2.43623805046082,
-2.43746805191040,
-2.43869853019714,
-2.43992924690247,
-2.44116020202637,
-2.44239139556885,
-2.44362306594849,
-2.44485497474670,
-2.44608712196350,
-2.44731950759888,
-2.44855237007141,
-2.44978547096252,
-2.45101881027222,
-2.45225238800049,
-2.45348644256592,
-2.45472073554993,
-2.45595526695251,
-2.45719003677368,
-2.45842528343201,
-2.45966076850891,
-2.46089649200439,
-2.46213245391846,
-2.46336889266968,
-2.46460556983948,
-2.46584248542786,
-2.46707963943481,
-2.46831727027893,
-2.46955513954163,
-2.47079324722290,
-2.47203159332275,
-2.47327017784119,
-2.47450923919678,
-2.47574853897095,
-2.47698807716370,
-2.47822785377502,
-2.47946810722351,
-2.48070859909058,
-2.48194932937622,
-2.48319029808044,
-2.48443174362183,
-2.48567342758179,
-2.48691534996033,
-2.48815751075745,
-2.48940014839172,
-2.49064302444458,
-2.49188613891602,
-2.49312949180603,
-2.49437308311462,
-2.49561715126038,
-2.49686145782471,
-2.49810600280762,
-2.49935078620911,
-2.50059604644775,
-2.50184154510498,
-2.50308728218079,
-2.50433325767517,
-2.50557947158813,
-2.50682616233826,
-2.50807309150696,
-2.50932025909424,
-2.51056766510010,
-2.51181554794312,
-2.51306366920471,
-2.51431202888489,
-2.51556062698364,
-2.51680946350098,
-2.51805877685547,
-2.51930832862854,
-2.52055811882019,
-2.52180814743042,
-2.52305841445923,
-2.52430915832520,
-2.52556014060974,
-2.52681136131287,
-2.52806282043457,
-2.52931475639343,
-2.53056693077087,
-2.53181934356689,
-2.53307199478149,
-2.53432488441467,
-2.53557825088501,
-2.53683185577393,
-2.53808569908142,
-2.53933978080750,
-2.54059410095215,
-2.54184889793396,
-2.54310393333435,
-2.54435920715332,
-2.54561471939087,
-2.54687047004700,
-2.54812669754028,
-2.54938316345215,
-2.55063986778259,
-2.55189681053162,
-2.55315399169922,
-2.55441164970398,
-2.55566954612732,
-2.55692768096924,
-2.55818605422974,
-2.55944466590881,
-2.56070375442505,
-2.56196308135986,
-2.56322264671326,
-2.56448245048523,
-2.56574249267578,
-2.56700301170349,
-2.56826376914978,
-2.56952476501465,
-2.57078599929810,
-2.57204747200012,
-2.57330942153931,
-2.57457160949707,
-2.57583403587341,
-2.57709670066834,
-2.57835960388184,
-2.57962298393250,
-2.58088660240173,
-2.58215045928955,
-2.58341455459595,
-2.58467888832092,
-2.58594369888306,
-2.58720874786377,
-2.58847403526306,
-2.58973956108093,
-2.59100532531738,
-2.59227132797241,
-2.59353780746460,
-2.59480452537537,
-2.59607148170471,
-2.59733867645264,
-2.59860610961914,
-2.59987401962280,
-2.60114216804504,
-2.60241055488586,
-2.60367918014526,
-2.60494804382324,
-2.60621714591980,
-2.60748672485352,
-2.60875654220581,
-2.61002659797668,
-2.61129689216614,
-2.61256742477417,
-2.61383843421936,
-2.61510968208313,
-2.61638116836548,
-2.61765289306641,
-2.61892485618591,
-2.62019705772400,
-2.62146973609924,
-2.62274265289307,
-2.62401580810547,
-2.62528920173645,
-2.62656283378601,
-2.62783670425415,
-2.62911105155945,
-2.63038563728333,
-2.63166046142578,
-2.63293552398682,
-2.63421082496643,
-2.63548636436462,
-2.63676238059998,
-2.63803863525391,
-2.63931512832642,
-2.64059185981751,
-2.64186882972717,
-2.64314603805542,
-2.64442372322083,
-2.64570164680481,
-2.64697980880737,
-2.64825820922852,
-2.64953684806824,
-2.65081572532654,
-2.65209507942200,
-2.65337467193604,
-2.65465450286865,
-2.65593457221985,
-2.65721487998962,
-2.65849542617798,
-2.65977621078491,
-2.66105747222900,
-2.66233897209168,
-2.66362071037293,
-2.66490268707275,
-2.66618490219116,
-2.66746735572815,
-2.66875028610230,
-2.67003345489502,
-2.67131686210632,
-2.67260050773621,
-2.67388439178467,
-2.67516851425171,
-2.67645287513733,
-2.67773771286011,
-2.67902278900147,
-2.68030810356140,
-2.68159365653992,
-2.68287944793701,
-2.68416547775269,
-2.68545174598694,
-2.68673849105835,
-2.68802547454834,
-2.68931269645691,
-2.69060015678406,
-2.69188785552979,
-2.69317579269409,
-2.69446396827698,
-2.69575262069702,
-2.69704151153564,
-2.69833064079285,
-2.69962000846863,
-2.70090961456299,
-2.70219945907593,
-2.70348954200745,
-2.70478010177612,
-2.70607089996338,
-2.70736193656921,
-2.70865321159363,
-2.70994472503662,
-2.71123647689819,
-2.71252846717834,
-2.71382069587708,
-2.71511340141296,
-2.71640634536743,
-2.71769952774048,
-2.71899294853210,
-2.72028660774231,
-2.72158050537109,
-2.72287464141846,
-2.72416901588440,
-2.72546386718750,
-2.72675895690918,
-2.72805428504944,
-2.72934985160828,
-2.73064565658569,
-2.73194169998169,
-2.73323798179626,
-2.73453450202942,
-2.73583149909973,
-2.73712873458862,
-2.73842620849609,
-2.73972392082214,
-2.74102187156677,
-2.74232006072998,
-2.74361848831177,
-2.74491715431213,
-2.74621629714966,
-2.74751567840576,
-2.74881529808044,
-2.75011515617371,
-2.75141525268555,
-2.75271558761597,
-2.75401616096497,
-2.75531697273254,
-2.75661802291870,
-2.75791954994202,
-2.75922131538391,
-2.76052331924438,
-2.76182556152344,
-2.76312804222107,
-2.76443076133728,
-2.76573371887207,
-2.76703691482544,
-2.76834034919739,
-2.76964402198792,
-2.77094817161560,
-2.77225255966187,
-2.77355718612671,
-2.77486205101013,
-2.77616715431213,
-2.77747249603272,
-2.77877807617188,
-2.78008389472961,
-2.78138995170593,
-2.78269624710083,
-2.78400301933289,
-2.78531002998352,
-2.78661727905273,
-2.78792476654053,
-2.78923249244690,
-2.79054045677185,
-2.79184865951538,
-2.79315710067749,
-2.79446578025818,
-2.79577469825745,
-2.79708409309387,
-2.79839372634888,
-2.79970359802246,
-2.80101370811462,
-2.80232405662537,
-2.80363464355469,
-2.80494546890259,
-2.80625653266907,
-2.80756783485413,
-2.80887937545776,
-2.81019115447998,
-2.81150341033936,
-2.81281590461731,
-2.81412863731384,
-2.81544160842896,
-2.81675481796265,
-2.81806826591492,
-2.81938195228577,
-2.82069587707520,
-2.82201004028320,
-2.82332444190979,
-2.82463908195496,
-2.82595396041870,
-2.82726907730103,
-2.82858467102051,
-2.82990050315857,
-2.83121657371521,
-2.83253288269043,
-2.83384943008423,
-2.83516621589661,
-2.83648324012756,
-2.83780050277710,
-2.83911800384522,
-2.84043574333191,
-2.84175372123718,
-2.84307193756104,
-2.84439039230347,
-2.84570908546448,
-2.84702825546265,
-2.84834766387939,
-2.84966731071472,
-2.85098719596863,
-2.85230731964111,
-2.85362768173218,
-2.85494828224182,
-2.85626912117004,
-2.85759019851685,
-2.85891151428223,
-2.86023306846619,
-2.86155486106873,
-2.86287689208984,
-2.86419916152954,
-2.86552166938782,
-2.86684441566467,
-2.86816763877869,
-2.86949110031128,
-2.87081480026245,
-2.87213873863220,
-2.87346291542053,
-2.87478733062744,
-2.87611198425293,
-2.87743687629700,
-2.87876200675964,
-2.88008737564087,
-2.88141298294067,
-2.88273882865906,
-2.88406491279602,
-2.88539123535156,
-2.88671779632568,
-2.88804459571838,
-2.88937163352966,
-2.89069890975952,
-2.89202642440796,
-2.89335441589355,
-2.89468264579773,
-2.89601111412048,
-2.89733982086182,
-2.89866876602173,
-2.89999794960022,
-2.90132737159729,
-2.90265703201294,
-2.90398693084717,
-2.90531706809998,
-2.90664744377136,
-2.90797805786133,
-2.90930891036987,
-2.91064000129700,
-2.91197133064270,
-2.91330289840698,
-2.91463470458984,
-2.91596674919128,
-2.91729903221130,
-2.91863155364990,
-2.91996431350708,
-2.92129731178284,
-2.92263054847717,
-2.92396402359009,
-2.92529773712158,
-2.92663168907166,
-2.92796587944031,
-2.92930054664612,
-2.93063545227051,
-2.93197059631348,
-2.93330597877502,
-2.93464159965515,
-2.93597745895386,
-2.93731355667114,
-2.93864989280701,
-2.93998646736145,
-2.94132328033447,
-2.94266033172607,
-2.94399762153626,
-2.94533514976501,
-2.94667291641235,
-2.94801092147827,
-2.94934916496277,
-2.95068764686584,
-2.95202636718750,
-2.95336532592773,
-2.95470452308655,
-2.95604395866394,
-2.95738363265991,
-2.95872354507446,
-2.96006369590759,
-2.96140408515930,
-2.96274471282959,
-2.96408557891846,
-2.96542668342590,
-2.96676802635193,
-2.96810960769653,
-2.96945142745972,
-2.97079348564148,
-2.97213578224182,
-2.97347831726074,
-2.97482109069824,
-2.97616410255432,
-2.97750735282898,
-2.97885084152222,
-2.98019456863403,
-2.98153853416443,
-2.98288273811340,
-2.98422718048096,
-2.98557186126709,
-2.98691678047180,
-2.98826193809509,
-2.98960733413696,
-2.99095296859741,
-2.99229884147644,
-2.99364495277405,
-2.99499130249023,
-2.99633789062500,
-2.99768471717834,
-2.99903178215027,
-3.00037908554077,
-3.00172662734985,
-3.00307440757751,
-3.00442242622376,
-3.00577068328857,
-3.00711917877197,
-3.00846791267395,
-3.00981688499451,
-3.01116609573364,
-3.01251554489136,
-3.01386523246765,
-3.01521515846252,
-3.01656532287598,
-3.01791572570801,
-3.01926636695862,
-3.02061724662781,
-3.02196836471558,
-3.02331972122192,
-3.02467131614685,
-3.02602314949036,
-3.02737522125244,
-3.02872753143311,
-3.03008008003235,
-3.03143286705017,
-3.03278589248657,
-3.03413915634155,
-3.03549265861511,
-3.03684639930725,
-3.03820037841797,
-3.03955459594727,
-3.04090881347656,
-3.04226326942444,
-3.04361796379089,
-3.04497289657593,
-3.04632806777954,
-3.04768347740173,
-3.04903912544251,
-3.05039501190186,
-3.05175113677979,
-3.05310750007629,
-3.05446410179138,
-3.05582094192505,
-3.05717802047730,
-3.05853533744812,
-3.05989289283752,
-3.06125068664551,
-3.06260871887207,
-3.06396698951721,
-3.06532549858093,
-3.06668424606323,
-3.06804323196411,
-3.06940245628357,
-3.07076191902161,
-3.07212162017822,
-3.07348155975342,
-3.07484173774719,
-3.07620215415955,
-3.07756257057190,
-3.07892322540283,
-3.08028411865234,
-3.08164525032043,
-3.08300662040710,
-3.08436822891235,
-3.08573007583618,
-3.08709216117859,
-3.08845448493958,
-3.08981704711914,
-3.09117984771729,
-3.09254288673401,
-3.09390616416931,
-3.09526968002319,
-3.09663343429565,
-3.09799742698669,
-3.09936165809631,
-3.10072612762451,
-3.10209059715271,
-3.10345530509949,
-3.10482025146484,
-3.10618543624878,
-3.10755085945129,
-3.10891652107239,
-3.11028242111206,
-3.11164855957031,
-3.11301493644714,
-3.11438155174255,
-3.11574840545654,
-3.11711549758911,
-3.11848282814026,
-3.11985039710999,
-3.12121820449829,
-3.12258625030518,
-3.12395429611206,
-3.12532258033752,
-3.12669110298157,
-3.12805986404419,
-3.12942886352539,
-3.13079810142517,
-3.13216757774353,
-3.13353729248047,
-3.13490724563599,
-3.13627743721008,
-3.13764786720276,
-3.13901853561401,
-3.14038944244385,
-3.14176034927368,
-3.14313149452209,
-3.14450287818909,
-3.14587450027466,
-3.14724636077881,
-3.14861845970154,
-3.14999079704285,
-3.15136337280273,
-3.15273618698120,
-3.15410923957825,
-3.15548253059387,
-3.15685606002808,
-3.15822958946228,
-3.15960335731506,
-3.16097736358643,
-3.16235160827637,
-3.16372609138489,
-3.16510081291199,
-3.16647577285767,
-3.16785097122192,
-3.16922640800476,
-3.17060208320618,
-3.17197799682617,
-3.17335391044617,
-3.17473006248474,
-3.17610645294189,
-3.17748308181763,
-3.17885994911194,
-3.18023705482483,
-3.18161439895630,
-3.18299198150635,
-3.18436980247498,
-3.18574786186218,
-3.18712592124939,
-3.18850421905518,
-3.18988275527954,
-3.19126152992249,
-3.19264054298401,
-3.19401979446411,
-3.19539928436279,
-3.19677901268005,
-3.19815897941589,
-3.19953894615173,
-3.20091915130615,
-3.20229959487915,
-3.20368027687073,
-3.20506119728088,
-3.20644235610962,
-3.20782375335693,
-3.20920538902283,
-3.21058726310730,
-3.21196913719177,
-3.21335124969482,
-3.21473360061646,
-3.21611618995667,
-3.21749901771545,
-3.21888208389282,
-3.22026538848877,
-3.22164893150330,
-3.22303247451782,
-3.22441625595093,
-3.22580027580261,
-3.22718453407288,
-3.22856903076172,
-3.22995376586914,
-3.23133873939514,
-3.23272395133972,
-3.23410916328430,
-3.23549461364746,
-3.23688030242920,
-3.23826622962952,
-3.23965239524841,
-3.24103879928589,
-3.24242544174194,
-3.24381232261658,
-3.24519920349121,
-3.24658632278442,
-3.24797368049622,
-3.24936127662659,
-3.25074911117554,
-3.25213718414307,
-3.25352549552918,
-3.25491404533386,
-3.25630259513855,
-3.25769138336182,
-3.25908041000366,
-3.26046967506409,
-3.26185917854309,
-3.26324892044067,
-3.26463890075684,
-3.26602888107300,
-3.26741909980774,
-3.26880955696106,
-3.27020025253296,
-3.27159118652344,
-3.27298235893250,
-3.27437376976013,
-3.27576518058777,
-3.27715682983398,
-3.27854871749878,
-3.27994084358215,
-3.28133320808411,
-3.28272581100464,
-3.28411841392517,
-3.28551125526428,
-3.28690433502197,
-3.28829765319824,
-3.28969120979309,
-3.29108500480652,
-3.29247903823853,
-3.29387307167053,
-3.29526734352112,
-3.29666185379028,
-3.29805660247803,
-3.29945158958435,
-3.30084681510925,
-3.30224204063416,
-3.30363750457764,
-3.30503320693970,
-3.30642914772034,
-3.30782532691956,
-3.30922174453735,
-3.31061816215515,
-3.31201481819153,
-3.31341171264648,
-3.31480884552002,
-3.31620621681213,
-3.31760382652283,
-3.31900143623352,
-3.32039928436279,
-3.32179737091064,
-3.32319569587708,
-3.32459425926209,
-3.32599306106567,
-3.32739186286926,
-3.32879090309143,
-3.33019018173218,
-3.33158969879150,
-3.33298945426941,
-3.33438920974731,
-3.33578920364380,
-3.33718943595886,
-3.33858990669251,
-3.33999061584473,
-3.34139156341553,
-3.34279251098633,
-3.34419369697571,
-3.34559512138367,
-3.34699678421021,
-3.34839868545532,
-3.34980058670044,
-3.35120272636414,
-3.35260510444641,
-3.35400772094727,
-3.35541057586670,
-3.35681366920471,
-3.35821676254272,
-3.35962009429932,
-3.36102366447449,
-3.36242747306824,
-3.36383152008057,
-3.36523556709290,
-3.36663985252380,
-3.36804437637329,
-3.36944913864136,
-3.37085413932800,
-3.37225914001465,
-3.37366437911987,
-3.37506985664368,
-3.37647557258606,
-3.37788152694702,
-3.37928748130798,
-3.38069367408752,
-3.38210010528564,
-3.38350677490234,
-3.38491368293762,
-3.38632059097290,
-3.38772773742676,
-3.38913512229919,
-3.39054274559021,
-3.39195060729980,
-3.39335846900940,
-3.39476656913757,
-3.39617490768433,
-3.39758348464966,
-3.39899230003357,
-3.40040111541748,
-3.40181016921997,
-3.40321946144104,
-3.40462899208069,
-3.40603852272034,
-3.40744829177856,
-3.40885829925537,
-3.41026854515076,
-3.41167902946472,
-3.41308951377869,
-3.41450023651123,
-3.41591119766235,
-3.41732239723206,
-3.41873359680176,
-3.42014503479004,
-3.42155671119690,
-3.42296862602234,
-3.42438077926636,
-3.42579293251038,
-3.42720532417297,
-3.42861795425415,
-3.43003082275391,
-3.43144369125366,
-3.43285679817200,
-3.43427014350891,
-3.43568372726440,
-3.43709754943848,
-3.43851137161255,
-3.43992543220520,
-3.44133973121643,
-3.44275426864624,
-3.44416880607605,
-3.44558358192444,
-3.44699859619141,
-3.44841384887695,
-3.44982910156250,
-3.45124459266663,
-3.45266032218933,
-3.45407629013062,
-3.45549225807190,
-3.45690846443176,
-3.45832490921021,
-3.45974159240723,
-3.46115851402283,
-3.46257543563843,
-3.46399259567261,
-3.46540999412537,
-3.46682763099670,
-3.46824526786804,
-3.46966314315796,
-3.47108125686646,
-3.47249960899353,
-3.47391796112061,
-3.47533655166626,
-3.47675538063049,
-3.47817444801331,
-3.47959351539612,
-3.48101282119751,
-3.48243236541748,
-3.48385214805603,
-3.48527193069458,
-3.48669195175171,
-3.48811221122742,
-3.48953247070313,
-3.49095296859741,
-3.49237370491028,
-3.49379467964172,
-3.49521565437317,
-3.49663686752319,
-3.49805831909180,
-3.49948000907898,
-3.50090169906616,
-3.50232362747192,
-3.50374579429626,
-3.50516819953918,
-3.50659060478210,
-3.50801324844360,
-3.50943613052368,
-3.51085925102234,
-3.51228237152100,
-3.51370573043823,
-3.51512932777405,
-3.51655292510986,
-3.51797676086426,
-3.51940083503723,
-3.52082514762878,
-3.52224946022034,
-3.52367401123047,
-3.52509880065918,
-3.52652382850647,
-3.52794885635376,
-3.52937412261963,
-3.53079962730408,
-3.53222513198853,
-3.53365087509155,
-3.53507685661316,
-3.53650307655334,
-3.53792929649353,
-3.53935575485230,
-3.54078245162964,
-3.54220914840698,
-3.54363608360291,
-3.54506325721741,
-3.54649066925049,
-3.54791808128357,
-3.54934573173523,
-3.55077362060547,
-3.55220150947571,
-3.55362963676453,
-3.55505800247192,
-3.55648636817932,
-3.55791497230530,
-3.55934381484985,
-3.56077289581299,
-3.56220197677612,
-3.56363129615784,
-3.56506085395813,
-3.56649041175842,
-3.56792020797730,
-3.56935024261475,
-3.57078027725220,
-3.57221055030823,
-3.57364106178284,
-3.57507181167603,
-3.57650256156921,
-3.57793354988098,
-3.57936477661133,
-3.58079600334168,
-3.58222746849060,
-3.58365917205811,
-3.58509087562561,
-3.58652281761169,
-3.58795499801636,
-3.58938717842102,
-3.59081959724426,
-3.59225225448608,
-3.59368515014648,
-3.59511804580688,
-3.59655117988586,
-3.59798455238342,
-3.59941792488098,
-3.60085153579712,
-3.60228538513184,
-3.60371923446655,
-3.60515332221985,
-3.60658764839172,
-3.60802197456360,
-3.60945653915405,
-3.61089134216309,
-3.61232614517212,
-3.61376118659973,
-3.61519646644592,
-3.61663174629211,
-3.61806726455688,
-3.61950302124023,
-3.62093877792358,
-3.62237477302551,
-3.62381100654602,
-3.62524724006653,
-3.62668371200562,
-3.62812042236328,
-3.62955713272095,
-3.63099408149719,
-3.63243126869202,
-3.63386845588684,
-3.63530588150024,
-3.63674354553223,
-3.63818120956421,
-3.63961911201477,
-3.64105725288391,
-3.64249539375305,
-3.64393377304077,
-3.64537239074707,
-3.64681100845337,
-3.64824986457825,
-3.64968895912170,
-3.65112805366516,
-3.65256738662720,
-3.65400695800781,
-3.65544652938843,
-3.65688633918762,
-3.65832614898682,
-3.65976619720459,
-3.66120648384094,
-3.66264677047730,
-3.66408729553223,
-3.66552805900574,
-3.66696882247925,
-3.66840982437134,
-3.66985106468201,
-3.67129230499268,
-3.67273378372192,
-3.67417550086975,
-3.67561721801758,
-3.67705917358398,
-3.67850112915039,
-3.67994332313538,
-3.68138575553894,
-3.68282818794251,
-3.68427085876465,
-3.68571376800537,
-3.68715667724609,
-3.68859982490540,
-3.69004321098328,
-3.69148659706116,
-3.69293022155762,
-3.69437384605408,
-3.69581770896912,
-3.69726181030273,
-3.69870591163635,
-3.70015025138855,
-3.70159482955933,
-3.70303940773010,
-3.70448422431946,
-3.70592904090881,
-3.70737409591675,
-3.70881938934326,
-3.71026468276978,
-3.71171021461487,
-3.71315574645996,
-3.71460151672363,
-3.71604752540588,
-3.71749353408813,
-3.71893978118897,
-3.72038626670837,
-3.72183275222778,
-3.72327947616577,
-3.72472620010376,
-3.72617316246033,
-3.72762036323547,
-3.72906756401062,
-3.73051500320435,
-3.73196244239807,
-3.73341012001038,
-3.73485803604126,
-3.73630595207214,
-3.73775410652161,
-3.73920226097107,
-3.74065065383911,
-3.74209928512573,
-3.74354791641235,
-3.74499678611755,
-3.74644565582275,
-3.74789476394653,
-3.74934411048889,
-3.75079345703125,
-3.75224304199219,
-3.75369262695313,
-3.75514245033264,
-3.75659251213074,
-3.75804257392883,
-3.75949287414551,
-3.76094317436218,
-3.76239371299744,
-3.76384425163269,
-3.76529502868652,
-3.76674604415894,
-3.76819705963135,
-3.76964831352234,
-3.77109956741333,
-3.77255105972290,
-3.77400279045105,
-3.77545452117920,
-3.77690649032593,
-3.77835845947266,
-3.77981066703796,
-3.78126287460327,
-3.78271532058716,
-3.78416800498962,
-3.78562068939209,
-3.78707361221313,
-3.78852653503418,
-3.78997969627380,
-3.79143285751343,
-3.79288625717163,
-3.79433989524841,
-3.79579353332520,
-3.79724740982056,
-3.79870128631592,
-3.80015540122986,
-3.80160951614380,
-3.80306386947632,
-3.80451822280884,
-3.80597281455994,
-3.80742764472961,
-3.80888247489929,
-3.81033754348755,
-3.81179261207581,
-3.81324791908264,
-3.81470322608948,
-3.81615877151489,
-3.81761431694031,
-3.81907010078430,
-3.82052612304688,
-3.82198214530945,
-3.82343840599060,
-3.82489466667175,
-3.82635116577148,
-3.82780766487122,
-3.82926440238953,
-3.83072113990784,
-3.83217811584473,
-3.83363533020020,
-3.83509254455566,
-3.83654999732971,
-3.83800745010376,
-3.83946514129639,
-3.84092283248901,
-3.84238076210022,
-3.84383869171143,
-3.84529685974121,
-3.84675502777100,
-3.84821343421936,
-3.84967184066772,
-3.85113048553467,
-3.85258913040161,
-3.85404801368713,
-3.85550713539124,
-3.85696625709534,
-3.85842561721802,
-3.85988497734070,
-3.86134457588196,
-3.86280417442322,
-3.86426401138306,
-3.86572384834290,
-3.86718392372131,
-3.86864399909973,
-3.87010431289673,
-3.87156462669373,
-3.87302517890930,
-3.87448573112488,
-3.87594652175903,
-3.87740731239319,
-3.87886834144592,
-3.88032937049866,
-3.88179063796997,
-3.88325190544128,
-3.88471341133118,
-3.88617491722107,
-3.88763666152954,
-3.88909840583801,
-3.89056038856506,
-3.89202237129211,
-3.89348459243774,
-3.89494705200195,
-3.89640951156616,
-3.89787220954895,
-3.89933490753174,
-3.90079784393311,
-3.90226078033447,
-3.90372395515442,
-3.90518712997437,
-3.90665054321289,
-3.90811395645142,
-3.90957736968994,
-3.91104102134705,
-3.91250467300415,
-3.91396856307983,
-3.91543245315552,
-3.91689658164978,
-3.91836071014404,
-3.91982507705688,
-3.92128944396973,
-3.92275404930115,
-3.92421865463257,
-3.92568349838257,
-3.92714834213257,
-3.92861342430115,
-3.93007850646973,
-3.93154382705688,
-3.93300914764404,
-3.93447470664978,
-3.93594026565552,
-3.93740606307983,
-3.93887186050415,
-3.94033789634705,
-3.94180393218994,
-3.94327020645142,
-3.94473648071289,
-3.94620299339294,
-3.94766950607300,
-3.94913625717163,
-3.95060300827026,
-3.95206975936890,
-3.95353674888611,
-3.95500373840332,
-3.95647096633911,
-3.95793819427490,
-3.95940566062927,
-3.96087312698364,
-3.96234083175659,
-3.96380853652954,
-3.96527647972107,
-3.96674442291260,
-3.96821260452271,
-3.96968078613281,
-3.97114896774292,
-3.97261738777161,
-3.97408580780029,
-3.97555446624756,
-3.97702312469482,
-3.97849202156067,
-3.97996091842651,
-3.98143005371094,
-3.98289918899536,
-3.98436856269836,
-3.98583793640137,
-3.98730731010437,
-3.98877692222595,
-3.99024653434753,
-3.99171638488770,
-3.99318623542786,
-3.99465632438660,
-3.99612641334534,
-3.99759650230408,
-3.99906682968140,
-4.00053739547730,
-4.00200796127319,
-4.00347852706909,
-4.00494909286499,
-4.00642013549805,
-4.00789117813110,
-4.00936222076416,
-4.01083326339722,
-4.01230430603027,
-4.01377582550049,
-4.01524734497070,
-4.01671886444092,
-4.01819038391113,
-4.01966190338135,
-4.02113389968872,
-4.02260589599609,
-4.02407789230347,
-4.02554988861084,
-4.02702236175537,
-4.02849483489990,
-4.02996730804443,
-4.03143978118897,
-4.03291225433350,
-4.03438520431519,
-4.03585815429688,
-4.03733110427856,
-4.03880405426025,
-4.04027700424194,
-4.04175043106079,
-4.04322385787964,
-4.04469728469849,
-4.04617071151733,
-4.04764413833618,
-4.04911804199219,
-4.05059194564819,
-4.05206584930420,
-4.05353975296021,
-4.05501365661621,
-4.05648803710938,
-4.05796241760254,
-4.05943679809570,
-4.06091117858887,
-4.06238555908203,
-4.06386041641235,
-4.06533527374268,
-4.06681013107300,
-4.06828498840332,
-4.06975984573364,
-4.07123517990112,
-4.07271051406860,
-4.07418584823608,
-4.07566118240356,
-4.07713651657105,
-4.07861232757568,
-4.08008813858032,
-4.08156394958496,
-4.08303976058960,
-4.08451557159424,
-4.08599185943604,
-4.08746814727783,
-4.08894443511963,
-4.09042072296143,
-4.09189701080322,
-4.09337329864502,
-4.09485006332398,
-4.09632682800293,
-4.09780359268189,
-4.09928035736084,
-4.10075712203980,
-4.10223436355591,
-4.10371160507202,
-4.10518884658814,
-4.10666608810425,
-4.10814332962036,
-4.10962104797363,
-4.11109876632690,
-4.11257648468018,
-4.11405420303345,
-4.11553192138672,
-4.11700963973999,
-4.11848783493042,
-4.11996603012085,
-4.12144422531128,
-4.12292242050171,
-4.12440061569214,
-4.12587928771973,
-4.12735795974731,
-4.12883663177490,
-4.13031530380249,
-4.13179397583008,
-4.13327264785767,
-4.13475179672241,
-4.13623094558716,
-4.13771009445190,
-4.13918924331665,
-4.14066839218140,
-4.14214754104614,
-4.14362716674805,
-4.14510679244995,
-4.14658641815186,
-4.14806604385376,
-4.14954566955566,
-4.15102529525757,
-4.15250539779663,
-4.15398550033569,
-4.15546560287476,
-4.15694570541382,
-4.15842580795288,
-4.15990591049194,
-4.16138648986816,
-4.16286706924439,
-4.16434764862061,
-4.16582822799683,
-4.16730880737305,
-4.16878938674927,
-4.17027044296265,
-4.17175149917603,
-4.17323255538940,
-4.17471361160278,
-4.17619466781616,
-4.17767572402954,
-4.17915725708008,
-4.18063879013062,
-4.18212032318115,
-4.18360185623169,
-4.18508338928223,
-4.18656492233276,
-4.18804693222046,
-4.18952894210815,
-4.19101095199585,
-4.19249296188355,
-4.19397497177124,
-4.19545698165894,
-4.19693899154663,
-4.19842147827148,
-4.19990396499634,
-4.20138645172119,
-4.20286893844605,
-4.20435142517090,
-4.20583391189575,
-4.20731687545776,
-4.20879983901978,
-4.21028280258179,
-4.21176576614380,
-4.21324872970581,
-4.21473169326782,
-4.21621465682983,
-4.21769809722900,
-4.21918153762817,
-4.22066497802734,
-4.22214841842651,
-4.22363185882568,
-4.22511529922485,
-4.22659873962402,
-4.22808265686035,
-4.22956657409668,
-4.23105049133301,
-4.23253440856934,
-4.23401832580566,
-4.23550224304199,
-4.23698616027832,
-4.23847055435181,
-4.23995923995972,
-4.24218654632568,
-4.24287128448486,
-4.24619340896606,
-4.24561643600464,
-4.25053405761719,
-4.24785709381104,
-4.25124597549439,
-4.24905872344971,
-4.24626970291138,
-4.24938154220581,
-4.23249578475952,
-4.24874353408814,
-4.20635366439819,
-4.24792909622192,
-4.16295766830444,
-4.24252033233643,
-4.17368078231812,
-4.26464033126831,
-4.14904737472534,
-4.28827524185181,
-4.13068771362305,
-4.39835548400879,
-4.12333059310913,
-4.26282310485840,
-4.05759286880493,
-4.34411048889160,
-4.26688432693481,
-4.22456741333008,
-4.76027917861939,
-4.08250236511231,
-5.43543052673340,
-4.03710842132568,
-5.28371524810791,
-4.15645980834961,
-5.78961992263794,
-4.49025869369507,
-6.41181182861328,
-5.20756673812866,
-8.60256195068359,
-5.53817081451416,
26.9392089843750,
-7.84591436386108,
-30.4595489501953,
-12.0969829559326,
-3.08221220970154,
13.3848018646240,
10.9495410919189,
48.5289688110352,
32.9144248962402,
-15.7588062286377,
-0.349153041839600,
-0.781292438507080,
-13.9084806442261,
-14.0972366333008,
-54.3517723083496,
0.790834903717041,
59.6821899414063,
-44.3396453857422,
-16.0944061279297,
5.70932531356812,
2.17439794540405,
4.84311532974243,
-14.4090156555176,
31.9038925170898,
-27.4082031250000,
23.9800186157227,
12.7297153472900,
-52.3868904113770,
-15.4648761749268,
-11.0140447616577,
-15.1697998046875,
-52.6315574645996,
41.6278800964356,
31.1637268066406,
-32.8378639221191,
40.0957832336426,
31.0562667846680,
-22.9171409606934,
-54.9558868408203,
-7.10457468032837,
-18.0274810791016,
-14.9025173187256,
36.4758567810059,
-43.9849319458008,
-30.5716800689697,
5.05335235595703,
-35.7736015319824,
-4.75768184661865,
18.6046504974365,
-24.4997253417969,
0.0522370338439941,
49.7225418090820,
20.7230567932129,
41.0983734130859,
49.2214050292969,
55.0252990722656,
33.2417907714844,
-27.3901557922363,
-16.8656005859375,
5.65694141387939,
14.9300403594971,
15.2072982788086,
64.8196640014648,
-13.2164096832275,
4.85469913482666,
54.0829925537109,
-60.0157241821289,
9.88717937469482,
27.8120250701904,
29.1071434020996,
11.7082805633545,
-19.9756813049316,
48.2882118225098,
-17.6652202606201,
-49.7879066467285,
-12.1749458312988,
2.48234272003174,
52.6125450134277,
6.39780902862549,
-45.1225585937500,
29.8629684448242,
13.1679553985596,
-32.1842117309570,
-2.31591892242432,
32.0912666320801,
25.2400588989258,
-22.5875968933105,
30.9460506439209,
-11.7882337570190,
-23.5397300720215,
46.5229225158691,
-29.1739673614502,
30.0652561187744,
24.2947463989258,
-39.8393630981445,
5.52241897583008,
-38.1115608215332,
-7.91510868072510,
65.3200531005859,
-1.70755410194397,
4.17309236526489,
22.0694656372070,
-41.4797134399414,
16.1723804473877,
28.1840324401855,
26.3344116210938,
27.3679199218750,
-13.9621667861938,
7.18173980712891,
-10.8020038604736,
21.5335025787354,
35.5535278320313,
-47.2087554931641,
36.3846282958984,
30.4848155975342,
-21.0901908874512,
48.1425399780273,
-32.8453292846680,
-14.4393291473389,
9.95934581756592,
-47.4821853637695,
-15.7466964721680,
73.4372024536133,
-1.78488349914551,
-32.0309524536133,
65.0601043701172,
-2.14680099487305,
28.8578987121582,
3.43489789962769,
-14.5469198226929,
49.6382179260254,
44.8689079284668,
-13.6041851043701,
-3.94590449333191,
19.3995685577393,
-54.2783164978027,
-28.3898849487305,
6.73454856872559,
30.0382080078125,
9.60222148895264,
17.4200611114502,
-10.2129917144775,
4.24231863021851,
10.3164463043213,
-37.9153556823731,
16.3796367645264,
-23.7146167755127,
-10.2260341644287,
-9.68401718139648,
22.4457817077637,
45.4117279052734,
-11.3348026275635,
56.9796371459961,
-9.86338901519775,
-22.6914291381836,
90.7708969116211,
-5.52187013626099,
-37.5899314880371,
-11.7073230743408,
-1.47309970855713,
50.9735641479492,
17.5085906982422,
27.5478706359863,
37.8487091064453,
-10.1192893981934,
-58.4507179260254,
24.6897354125977,
8.22626304626465,
-38.0252227783203,
65.6377105712891,
2.97809171676636,
-20.5252037048340,
5.64750576019287,
-2.64566159248352,
9.65871715545654,
7.87186527252197,
32.0113525390625,
47.2705383300781,
-7.39634227752686,
17.7656326293945,
34.0230560302734,
-55.4530944824219,
29.2453079223633,
54.3610992431641,
9.35575866699219,
-12.1456651687622,
-37.2160110473633,
46.3289756774902,
-9.90006256103516,
-65.1661071777344,
23.6013832092285,
47.6516952514648,
-1.51801800727844,
18.5814704895020,
-32.8277015686035,
-30.1158428192139,
59.4227180480957,
-57.3968048095703,
39.2430267333984,
34.2403106689453,
-12.5524024963379,
32.3792190551758,
-51.5419692993164,
19.7374324798584,
-2.72233605384827,
39.4986534118652,
1.32845449447632,
-12.5883417129517,
48.0457878112793,
-27.8903617858887,
-20.3459682464600,
-25.5448474884033,
31.5947971343994,
35.1502151489258,
-3.37991714477539,
-12.5830421447754,
-10.4981994628906,
22.7390327453613,
24.4320850372314,
5.25825691223145,
-45.3204116821289,
4.00011920928955,
9.16945838928223,
-56.5967102050781,
-11.8328094482422,
28.6965560913086,
17.2843112945557,
6.85087966918945,
47.2897071838379,
-5.54755306243897,
-32.4747428894043,
48.5333557128906,
9.86152648925781,
7.47197914123535,
27.2131710052490,
-45.5067443847656,
16.1935634613037,
41.2232398986816,
-52.3740310668945,
10.3741455078125,
31.3089141845703,
-1.93109607696533,
-19.4943199157715,
-42.8717651367188,
-13.9533996582031,
-29.7602653503418,
-30.1876144409180,
18.2308597564697,
1.14473390579224,
-52.1790542602539,
24.8010807037354,
-20.2451782226563,
-61.2719573974609,
73.5298309326172,
15.7295837402344,
9.20408821105957,
-15.9727172851563,
-2.65994453430176,
37.5392189025879,
-52.7409210205078,
58.5831527709961,
31.2819976806641,
-44.3801116943359,
4.90258026123047,
3.94485616683960,
-37.0306015014648,
-18.5470638275147,
17.0799388885498,
30.2495021820068,
29.2134990692139,
4.82019853591919,
33.3511161804199,
-27.0348129272461,
23.3999214172363,
6.07450056076050,
-27.2983474731445,
37.0920104980469,
22.2385540008545,
49.8981361389160,
-9.69439697265625,
-1.86930060386658,
62.7852592468262,
19.3757419586182,
-26.6205177307129,
21.4993610382080,
-17.5127754211426,
-34.6080398559570,
56.0639152526856,
-28.2400703430176,
-30.0737228393555,
-21.4755687713623,
-8.29751396179199,
40.4286041259766,
-15.9480857849121,
4.89804029464722,
-36.2880210876465,
11.7032527923584,
15.6558227539063,
8.93527030944824,
60.5577735900879,
-56.6532592773438,
42.2714347839356,
35.6891517639160,
-3.34716796875000,
23.1807727813721,
-49.1387100219727,
34.2822608947754,
-21.7052478790283,
14.6481513977051,
33.8546180725098,
-67.9336776733398,
-20.5886478424072,
22.5034828186035,
29.6507835388184,
-63.9120330810547,
-33.7732925415039,
-12.4313449859619,
-36.8757667541504,
17.5551033020020,
7.96669578552246,
-10.4771051406860,
-0.940095901489258,
65.1168289184570,
-9.05950546264648,
-34.1903152465820,
36.8330039978027,
-5.67955303192139,
-13.5464534759521,
-18.6965942382813,
19.0252113342285,
40.6135406494141,
16.0664710998535,
-22.8519439697266,
10.1157655715942,
8.17700099945068,
-49.5624465942383,
65.7743148803711,
29.1304206848145,
-22.2370643615723,
19.7372627258301,
-21.8360519409180,
22.1601524353027,
10.5317144393921,
-66.2114410400391,
5.44521665573120,
-2.33450603485107,
-49.0079727172852,
49.6831092834473,
-2.27448511123657,
-1.19767928123474,
-10.5849056243896,
-55.5888557434082,
33.0468673706055,
-31.9533977508545,
24.4930210113525,
4.44312381744385,
-40.8159599304199,
34.2297439575195,
-33.8874206542969,
40.8925285339356,
35.5461807250977,
-11.8683719635010,
0.705768585205078,
20.1473045349121,
41.3837966918945,
2.17886209487915,
33.8349533081055,
9.23056125640869,
-39.0672836303711,
10.0631170272827,
28.7926177978516,
-56.6590919494629,
-8.62992858886719,
-12.9184103012085,
-70.8980407714844,
5.92291688919067,
6.73135375976563,
-27.7370491027832,
16.1419086456299,
31.6907272338867,
-59.5578727722168,
-17.0586490631104,
44.4171180725098,
5.61831235885620,
24.7960166931152,
57.0832862854004,
7.93701171875000,
-19.5262622833252,
89.1594390869141,
9.88194274902344,
-30.7514686584473,
46.5597534179688,
-43.0414466857910,
-15.5006713867188,
4.08998727798462,
-8.41531372070313,
10.6638412475586,
-13.4738273620605,
1.17269229888916,
50.0104293823242,
-4.05683231353760,
-23.2940025329590,
63.6328697204590,
-57.3349990844727,
-24.6999053955078,
74.7725219726563,
13.3115510940552,
-16.8700809478760,
-35.7460212707520,
-28.7629470825195,
-14.5434417724609,
68.4465637207031,
1.89004325866699,
-51.0601730346680,
42.2911720275879,
31.5009555816650,
-11.0407047271729,
-10.5305280685425,
44.5529937744141,
-19.1131572723389,
-16.0340957641602,
47.4349708557129,
-47.1195297241211,
26.8875389099121,
36.4969863891602,
-51.3997039794922,
-31.5315189361572,
-20.2503948211670,
34.0966072082520,
11.8777484893799,
33.1340446472168,
25.3719482421875,
-10.7632255554199,
45.9503250122070,
-29.6600914001465,
-9.61540412902832,
-0.803284645080566,
-53.5409469604492,
7.14341259002686,
-31.0412597656250,
-42.1375389099121,
17.1356620788574,
29.4329757690430,
-2.20388197898865,
9.49730110168457,
-2.93929910659790,
-44.5160522460938,
-16.5268669128418,
35.8902740478516,
18.1616973876953,
-61.3567161560059,
20.9435997009277,
2.46176719665527,
4.86137628555298,
46.7772407531738,
-28.5264549255371,
25.9548969268799,
-7.64263677597046,
15.8140373229980,
40.9894180297852,
-12.0397987365723,
-26.3353843688965,
1.21963310241699,
12.8342361450195,
-33.2545928955078,
21.1225852966309,
-48.3275680541992,
-34.1036529541016,
49.3121643066406,
-15.5349702835083,
40.6693229675293,
8.61123847961426,
-45.1780433654785,
15.9065647125244,
-40.7513160705566,
-14.6573915481567,
0.429886817932129,
4.16623592376709,
44.8247566223145,
30.7222404479980,
48.4793243408203,
-20.8400115966797,
-18.1486244201660,
-29.9379158020020,
14.9557046890259,
29.9821052551270,
6.10617446899414,
48.8926391601563,
-19.9755973815918,
8.18410491943359,
0.496086120605469,
-35.0985450744629,
8.18108558654785,
-5.08301210403442,
-67.1209869384766,
34.9884529113770,
6.40088081359863,
-35.3746376037598,
22.2977485656738,
-51.3824462890625,
3.22015476226807,
-23.9096488952637,
3.57452869415283,
43.2669258117676,
27.0498619079590,
23.9818649291992,
6.61959505081177,
49.6190185546875,
20.0515537261963,
29.8598899841309,
38.5686721801758,
-5.98092842102051,
-38.8064994812012,
-12.1531047821045,
-11.3990688323975,
-38.2565727233887,
-36.1641464233398,
-26.9436473846436,
-5.43043422698975,
-14.5679988861084,
-48.2407264709473,
-3.30516195297241,
4.25544929504395,
1.55964422225952,
47.8690147399902,
-12.4842624664307,
32.1350746154785,
18.4819927215576,
18.2281188964844,
48.8453750610352,
-3.25663471221924,
27.5547924041748,
42.4285850524902,
-12.2835178375244,
-30.2143554687500,
64.2547760009766,
5.48330307006836,
-3.20397472381592,
11.5258378982544,
9.67572402954102,
17.2865829467773,
-26.2054157257080,
-6.93700885772705,
-38.1617012023926,
13.0262489318848,
-31.4686279296875,
-52.5379333496094,
-0.731255054473877,
-16.4478454589844,
33.5799293518066,
-8.92671298980713,
-30.6737003326416,
63.7196006774902,
-8.14074707031250,
-40.2887992858887,
50.1143760681152,
-41.9877700805664,
-8.80143737792969,
53.1582908630371,
-13.5895404815674,
30.8059062957764,
8.70056533813477,
-26.5358428955078,
13.6507129669189,
21.0416965484619,
-16.5793476104736,
-34.4412002563477,
44.7587013244629,
13.6928539276123,
-35.9357185363770,
15.9392538070679,
13.3869075775146,
-3.24725866317749,
-18.1799335479736,
43.1724243164063,
36.3619689941406,
32.7905921936035,
14.5906009674072,
-39.2388458251953,
26.9198436737061,
-20.8504962921143,
12.6495609283447,
33.7231101989746,
24.8366317749023,
7.99161338806152,
-17.5783195495605,
13.6697931289673,
-20.0152873992920,
34.8162078857422,
-19.3272552490234,
-37.9405288696289,
31.0439548492432,
14.2863779067993,
-40.5402336120606,
-2.11934375762939,
38.0919189453125,
-11.5101442337036,
-5.93047618865967,
36.3462944030762,
16.1689910888672,
-46.4784545898438,
35.5362396240234,
4.81446695327759,
-21.6454620361328,
-14.3938083648682,
-22.4662971496582,
35.1263465881348,
11.2297296524048,
13.2148265838623,
-38.6230354309082,
29.3320007324219,
14.7978439331055,
-52.0982398986816,
24.9197559356689,
-36.4869384765625,
17.3196372985840,
18.7732849121094,
-46.5914115905762,
-0.367571830749512,
22.7740192413330,
-9.11990356445313,
-45.1363067626953,
-30.0215511322022,
-2.04478740692139,
6.09706163406372,
-62.5121078491211,
50.3831481933594,
1.11219024658203,
-29.6118202209473,
47.3212776184082,
-63.7463073730469,
7.14050436019898,
40.4603881835938,
-16.0079402923584,
-47.8637924194336,
47.5058517456055,
11.1811962127686,
-31.3219356536865,
5.35511112213135,
5.69040393829346,
27.9443588256836,
-31.5172424316406,
42.3686561584473,
-14.6855707168579,
-33.9506912231445,
17.2313137054443,
15.1921215057373,
36.9248352050781,
16.7287254333496,
17.4640998840332,
-50.4444274902344,
-18.6435203552246,
-9.67684936523438,
-13.1500740051270,
52.5321121215820,
25.5554046630859,
34.4419708251953,
6.72962331771851,
-6.02201557159424,
18.5696144104004,
-26.5435848236084,
-26.8513755798340,
-11.9966688156128,
-0.242864608764648,
-13.1754894256592,
-0.714519977569580,
46.6646385192871,
-5.62848186492920,
3.65492343902588,
54.9710083007813,
11.1602287292480,
-19.4132766723633,
-45.4949951171875,
3.36691522598267,
32.8793258666992,
-49.0222854614258,
33.6953887939453,
59.8555412292481,
-46.4436492919922,
36.3515701293945,
66.2831802368164,
-18.5186786651611,
-16.6702842712402,
3.63463640213013,
41.8375816345215,
38.3228149414063,
-50.1678314208984,
-22.9469680786133,
31.7066841125488,
-36.9280014038086,
-47.6451530456543,
-12.1909809112549,
-31.2021503448486,
-52.5770454406738,
-28.6866645812988,
-14.7693328857422,
-11.3422603607178,
10.9707298278809,
-20.5038394927979,
5.91078662872314,
-32.5570411682129,
-52.8900604248047,
62.5120887756348,
-9.44603824615479,
12.1094121932983,
11.0815925598145,
-17.3461055755615,
37.9702796936035,
-41.3965492248535,
1.77085876464844,
18.9146156311035,
-3.97207522392273,
-32.0345687866211,
12.9092521667480,
27.4138412475586,
-26.3047790527344,
27.5214557647705,
12.7335433959961,
46.4495429992676,
24.5922393798828,
-8.51954269409180,
23.3466014862061,
41.2100601196289,
54.3297882080078,
2.56944227218628,
5.27882003784180,
21.5247707366943,
-13.0667781829834,
-8.51568698883057,
29.3319244384766,
-12.9832305908203,
-57.4474296569824,
-6.70190191268921,
-19.2299652099609,
-36.0052909851074,
0.416480064392090,
23.2873344421387,
38.9731674194336,
22.8507633209229,
10.1552476882935,
-28.7932090759277,
7.65492725372314,
-10.8446931838989,
-45.7542724609375,
29.1343803405762,
19.7184867858887,
37.5542907714844,
30.9972000122070,
35.9285736083984,
10.3908395767212,
21.9438400268555,
15.8930053710938,
-41.3455963134766,
39.8292388916016,
0.728384494781494,
-1.54977416992188,
43.0209236145020,
46.6454658508301,
-29.2149295806885,
-16.2337303161621,
12.3780403137207,
-36.6877212524414,
58.0820388793945,
0.567758560180664,
2.75795888900757,
-22.4996871948242,
-36.1057968139648,
3.46154165267944,
-27.3498821258545,
66.9172821044922,
-37.1230354309082,
-17.4116439819336,
49.1760864257813,
-41.1472244262695,
62.6500892639160,
33.2405509948731,
-22.8296508789063,
15.4839458465576,
7.62145185470581,
36.9555244445801,
31.8364582061768,
1.64775562286377,
22.9223709106445,
40.9183197021484,
26.2687835693359,
27.6589965820313,
-4.99673461914063,
27.8601989746094,
30.2265987396240,
-49.0298728942871,
-25.4237918853760,
29.3223609924316,
14.4732780456543,
0.725495815277100,
11.5170106887817,
-60.0580825805664,
-27.8508148193359,
56.6199569702148,
37.0245857238770,
36.1917800903320,
-22.1989860534668,
-49.3303871154785,
21.0645389556885,
52.0809974670410,
20.7659778594971,
-34.3145599365234,
-14.5489406585693,
39.2163619995117,
24.0560836791992,
-16.2691345214844,
59.1018066406250,
52.0185127258301,
-61.1382827758789,
37.4191665649414,
55.5788612365723,
-42.0956420898438,
-20.1827507019043,
-16.8031139373779,
21.6749382019043,
29.2558040618897,
-37.4601554870606,
-25.3849601745605,
7.59809303283691,
-36.9904212951660,
-30.7917289733887,
54.2421379089356,
-18.0944366455078,
-13.9764442443848,
60.6580200195313,
25.9965953826904,
18.3178710937500,
26.0118961334229,
17.2543220520020,
-28.8657073974609,
21.7605590820313,
-4.34109592437744,
8.37021732330322,
31.4311027526855,
-34.5369529724121,
68.5484542846680,
18.0178146362305,
-53.0503311157227,
25.3127288818359,
47.3001823425293,
-9.89896202087402,
10.6509208679199,
60.1761360168457,
-10.5674438476563,
59.1221923828125,
16.8244380950928,
-15.0147876739502,
28.7494125366211,
-37.1655883789063,
44.6003570556641,
5.41577291488648,
-47.7167205810547,
11.7333507537842,
34.0819168090820,
-19.6998519897461,
23.5566959381104,
33.6477622985840,
-25.8316726684570,
45.4504547119141,
18.2540225982666,
37.7342567443848,
-4.63550472259522,
-5.24872827529907,
30.8258323669434,
-31.5118923187256,
1.78628206253052,
9.73937034606934,
21.2492980957031,
-3.52434849739075,
-10.5273818969727,
47.6376914978027,
31.2034034729004,
-10.5397033691406,
-16.1096935272217,
-9.46252632141113,
23.0041561126709,
16.9564990997314,
9.40167617797852,
68.2154998779297,
18.1917438507080,
-43.5075798034668,
-7.41991424560547,
45.2285690307617,
49.0664901733398,
13.2054100036621,
0.114472866058350,
-33.9748420715332,
16.7678184509277,
5.34593057632446,
-26.9271450042725,
47.5266189575195,
43.2022171020508,
11.5154762268066,
-35.9345474243164,
4.17036485671997,
26.5197391510010,
-24.7012348175049,
30.2692375183105,
26.3282318115234,
5.92150831222534,
49.4578323364258,
9.98258686065674,
-43.2343215942383,
60.6823196411133,
35.2076530456543,
-60.7069702148438,
35.9991035461426,
2.71769380569458,
1.56110143661499,
7.53889989852905,
-19.4558849334717,
15.2923259735107,
-35.4668807983398,
-4.69094562530518,
54.4329032897949,
36.0376052856445,
-51.2420310974121,
-44.9558258056641,
33.6296844482422,
34.9021759033203,
-32.9430618286133,
-13.5421047210693,
37.0364990234375,
-38.7727699279785,
14.1167602539063,
55.9397926330566,
-8.77398109436035,
17.4438323974609,
25.7808876037598,
23.6786117553711,
46.7577590942383,
7.06227493286133,
14.0988655090332,
64.8570556640625,
5.12862396240234,
-23.8351840972900,
75.3082733154297,
5.85481882095337,
-46.7173271179199,
67.4647827148438,
-23.6155090332031,
-38.2464790344238,
48.2499084472656,
50.4263992309570,
10.3998155593872,
-48.1909446716309,
-24.7377128601074,
-9.51818656921387,
39.1378135681152,
-23.2739562988281,
-52.6404151916504,
50.9647064208984,
1.50051021575928,
-39.3800811767578,
27.0970191955566,
-4.40380620956421,
-29.3895816802979,
26.6166000366211,
18.9000778198242,
18.7092189788818,
-34.2313880920410,
-20.3114624023438,
33.5479164123535,
0.306282520294189,
24.7868080139160,
40.4336814880371,
12.7526779174805,
-15.9530372619629,
9.72197341918945,
4.80179691314697,
41.8675842285156,
59.5322570800781,
-6.24251365661621,
50.2907409667969,
25.3031768798828,
5.26008272171021,
-24.0293273925781,
-14.2398471832275,
50.8514747619629,
-14.9703025817871,
32.4199943542481,
-23.6456031799316,
-6.78447055816650,
51.5698127746582,
-29.0934104919434,
12.7205886840820,
35.9825363159180,
60.2122039794922,
-21.5277938842773,
-32.3963775634766,
12.5171985626221,
-25.8302001953125,
17.0017051696777,
-29.8092651367188,
-31.9674911499023,
23.3874626159668,
12.2388858795166,
-36.2111701965332,
-48.4040565490723,
-12.4595680236816,
20.2689552307129,
4.39797306060791,
-7.66259241104126,
60.1073379516602,
6.06513071060181,
-11.0360889434814,
-20.9776039123535,
14.8060016632080,
80.3777313232422,
-18.9436912536621,
-7.69954395294189,
20.3994560241699,
-1.88869571685791,
24.7407951354980,
8.59977531433106,
-27.4582519531250,
40.0053825378418,
17.2756576538086,
-39.0602111816406,
-5.61927223205566,
-55.0636482238770,
-19.4380455017090,
-26.2065067291260,
-25.6210479736328,
45.1412353515625,
-10.3432483673096,
-3.47525978088379,
1.12128496170044,
15.6611127853394,
-12.5236072540283,
-51.2677345275879,
9.44502830505371,
18.2951984405518,
24.3606910705566,
-45.6778335571289,
11.6301059722900,
44.5796737670898,
-52.4210510253906,
17.2820529937744,
10.8280372619629,
26.6907272338867,
1.40242099761963,
-35.9725952148438,
49.6680030822754,
-58.0736274719238,
-25.1340293884277,
33.7762527465820,
-54.4978904724121,
-12.0683584213257,
-11.3062267303467,
12.7009048461914,
41.0709877014160,
41.3743934631348,
-22.6533298492432,
-25.3998126983643,
7.42424154281616,
-40.1047363281250,
26.9912242889404,
-37.9832305908203,
-58.3229827880859,
44.6782112121582,
32.3998718261719,
-3.98142671585083,
3.31740570068359,
40.5401268005371,
39.6782035827637,
1.32826566696167,
-29.9287128448486,
-13.3292207717896,
24.6149177551270,
-6.53544569015503,
-48.7806053161621,
44.4906387329102,
20.2218246459961,
-22.4500732421875,
-3.43884849548340,
-22.3742065429688,
-12.5867061614990,
-44.8675270080566,
-2.92459869384766,
-36.4582061767578,
-21.2821712493897,
45.8256187438965,
-14.8952808380127,
14.8785266876221,
24.7640514373779,
-17.4385452270508,
-10.6513423919678,
-4.51867103576660,
-22.3279323577881,
-21.0854701995850,
1.45525884628296,
-39.2731246948242,
-24.5203094482422,
40.3468093872070,
26.1523036956787,
-2.17440986633301,
-57.0237693786621,
21.1921291351318,
20.2491149902344,
-54.2987403869629,
64.9168853759766,
6.83251714706421,
-62.0270309448242,
7.33571100234985,
10.1191444396973,
-30.4102096557617,
-27.5177898406982,
-6.08029270172119,
-25.9384994506836,
29.2586269378662,
13.0220832824707,
-37.1918411254883,
-11.8935184478760,
-24.5644340515137,
-21.8181610107422,
-21.2756881713867,
-39.6231002807617,
-29.6497459411621,
-6.67402982711792,
-18.6304264068604,
-9.79003906250000,
-2.76857280731201,
-23.8219051361084,
-12.9184608459473,
-32.1314201354981,
-7.93708324432373,
1.52200508117676,
-30.6018924713135,
-35.5666656494141,
-34.6269302368164,
36.8103637695313,
-17.6897468566895,
-56.2437667846680,
48.4058265686035,
17.0830059051514,
-5.42598772048950,
14.7103881835938,
-29.1184349060059,
-22.8304996490479,
-1.54669618606567,
-61.5249099731445,
-24.7109928131104,
39.2357254028320,
17.9102058410645,
16.1914196014404,
-19.1244277954102,
4.98280620574951,
-10.2371406555176,
-34.4021606445313,
-7.63918209075928,
3.29615783691406,
-21.3216838836670,
-59.0639572143555,
-14.4584102630615,
15.1002235412598,
28.8203468322754,
23.3395595550537,
47.7016601562500,
-6.60561418533325,
-32.1816787719727,
1.33650159835815,
-33.2814407348633,
6.53605318069458,
44.6103134155273,
5.03424596786499,
-2.83738136291504,
61.7556343078613,
-34.2969589233398,
-24.6533317565918,
51.3456916809082,
-1.85156393051147,
13.7455091476440,
-9.19905090332031,
-31.2492103576660,
-15.9925603866577,
-10.6447753906250,
-31.4289932250977,
6.88136529922485,
46.7334709167481,
-41.7887382507324,
-29.4366683959961,
68.8814163208008,
-9.69806861877441,
-42.4166526794434,
58.6526107788086,
-31.8309612274170,
-39.0302391052246,
52.5531463623047,
3.26943683624268,
27.3107376098633,
-16.3996829986572,
-32.2299499511719,
21.9001121520996,
27.2806701660156,
19.8917846679688,
-10.5002231597900,
31.3686599731445,
9.33357143402100,
6.89742851257324,
18.3817176818848,
39.2022438049316,
48.1795425415039,
-39.7484970092773,
25.8912658691406,
9.76290893554688,
-54.7727775573731,
-24.6609191894531,
-20.1480140686035,
-24.4780235290527,
-0.381937503814697,
22.0766181945801,
4.61723804473877,
35.2612762451172,
-20.9094219207764,
21.7839508056641,
9.58888244628906,
-4.97079706192017,
24.4683055877686,
-47.8698196411133,
43.7867965698242,
9.19955825805664,
16.6573848724365,
61.0752334594727,
-9.28165435791016,
-32.1894378662109,
-34.5238265991211,
12.6710605621338,
24.4594821929932,
19.8377952575684,
-8.72449684143066,
-30.0744819641113,
22.7485084533691,
30.1614265441895,
39.1990203857422,
34.9983558654785,
-24.4066314697266,
-23.4123325347900,
-4.76666069030762,
66.9770202636719,
-5.41577053070068,
-18.0112571716309,
55.9204254150391,
-54.5554618835449,
-28.6222705841064,
-20.0032196044922,
-23.6710109710693,
2.47992086410522,
-46.3803482055664,
-45.3258514404297,
-8.38037014007568,
-34.3518753051758,
-37.4733924865723,
12.1968336105347,
-18.3622817993164,
8.29237365722656,
1.69834852218628,
8.13263416290283,
29.7019405364990,
17.8297824859619,
20.9609031677246,
-40.8824729919434,
0.185520172119141,
-6.99424791336060,
-37.2783164978027,
5.76281118392944,
-50.1348800659180,
27.7933464050293,
52.9258842468262,
-48.7271499633789,
50.6308288574219,
0.837258338928223,
-58.8101005554199,
-12.5868330001831,
-39.4494590759277,
16.4241580963135,
-32.2664718627930,
25.1618156433105,
61.3748283386231,
-39.1277046203613,
14.7435493469238,
-25.2561836242676,
-19.3613090515137,
29.8852806091309,
-2.28423070907593,
10.3639192581177,
3.97831821441650,
-24.9047183990479,
-8.74718284606934,
35.5866394042969,
12.9686126708984,
27.1703910827637,
4.49760723114014,
23.3766403198242,
49.8461837768555,
-40.2798004150391,
-18.0031051635742,
48.0227851867676,
19.1882514953613,
-3.59050226211548,
49.4799079895020,
-3.99603176116943,
-1.19150447845459,
50.9748535156250,
15.4636459350586,
7.89292812347412,
10.9432334899902,
-8.38905906677246,
-27.0640563964844,
1.51669788360596,
13.3372087478638,
34.7860260009766,
24.3886604309082,
48.3614768981934,
-2.16307115554810,
-53.7028465270996,
64.6255187988281,
-6.61669111251831,
-38.2056884765625,
68.9505310058594,
22.7159767150879,
-43.5664863586426,
-14.8243370056152,
10.0265903472900,
-13.6338291168213,
-5.90135478973389,
-12.1802206039429,
43.1082153320313,
20.3526115417480,
7.84412050247192,
18.4250679016113,
-39.6058006286621,
46.6289825439453,
-38.5267944335938,
-8.86999511718750,
61.8519210815430,
-43.2968597412109,
-2.16153764724731,
19.0798740386963,
27.2998466491699,
-29.4764232635498,
25.5365219116211,
30.7814102172852,
-60.4366416931152,
13.4405841827393,
-24.8942375183105,
11.8905429840088,
31.4191799163818,
19.5310363769531,
72.9411849975586,
4.02274370193481,
-41.4594154357910,
3.28608512878418,
16.0925979614258,
-55.5050354003906,
4.96966791152954,
29.1856079101563,
-45.5744895935059,
-46.1986656188965,
-6.00174570083618,
-12.6463479995728,
-5.16794633865356,
22.1437644958496,
-1.92335891723633,
5.01855278015137,
-2.02635574340820,
50.0506134033203,
27.0798645019531,
23.9355926513672,
61.2527999877930,
15.0567808151245,
60.1340789794922,
23.7884941101074,
8.55494308471680,
47.9445037841797,
-26.0486869812012,
35.3997268676758,
58.4014129638672,
-50.1005630493164,
-20.0026569366455,
13.9603271484375,
-4.40931892395020,
4.54914855957031,
49.4317207336426,
23.6887702941895,
-10.6147193908691,
10.2847719192505,
14.9680538177490,
3.41373538970947,
-41.4396095275879,
20.1096191406250,
5.78665304183960,
-52.2771186828613,
56.2298698425293,
15.6693058013916,
-44.0303039550781,
46.8205223083496,
47.7529373168945,
21.3059921264648,
25.4318256378174,
-11.2378187179565,
42.3772659301758,
68.7385101318359,
-15.2603683471680,
-30.0233802795410,
-22.7930202484131,
-10.4331464767456,
-1.76078748703003,
-24.8485240936279,
-35.5260162353516,
-14.3129968643188,
-45.9287338256836,
-57.0741310119629,
49.2749099731445,
1.36548662185669,
-51.8887596130371,
15.3586635589600,
-33.0144653320313,
-18.9801025390625,
26.5289783477783,
2.65281534194946,
9.93250465393066,
25.4833431243897,
-8.67187118530273,
-5.95359563827515,
44.0370330810547,
-11.1633472442627,
7.91110754013062,
-15.1236715316772,
-30.6818561553955,
16.8135089874268,
-25.7368602752686,
-1.07037019729614,
-27.6052093505859,
7.73984479904175,
24.2824134826660,
-38.4119720458984,
-23.5791454315186,
10.2814426422119,
-3.07750058174133,
-1.34043598175049,
40.0045204162598,
35.2342185974121,
-12.3349361419678,
-21.3355178833008,
64.4983596801758,
-8.41127014160156,
12.6916179656982,
38.2461967468262,
-4.54088401794434,
38.4349861145020,
-14.1413078308105,
1.60019540786743,
-23.4048118591309,
39.3420410156250,
11.7637119293213,
-56.2582969665527,
41.7586860656738,
-10.7362079620361,
-16.4042148590088,
18.9550724029541,
39.4283409118652,
31.6881065368652,
-33.3586196899414,
15.3503417968750,
35.8232269287109,
1.19039678573608,
-18.4501552581787,
-29.9493312835693,
45.3147888183594,
1.38241529464722,
-70.1900177001953,
3.90069818496704,
51.9618072509766,
18.6741065979004,
19.0017337799072,
2.59359550476074,
-34.6701316833496,
29.7488269805908,
-17.6790695190430,
-17.5266036987305,
-2.65011429786682,
-65.1567459106445,
-16.1877727508545,
34.6518325805664,
24.5628814697266,
15.8010845184326,
32.2744789123535,
-48.1024551391602,
7.48382186889648,
81.1162338256836,
-19.4572830200195,
-44.3809471130371,
-10.9739446640015,
22.3029861450195,
-7.49676609039307,
-2.06964445114136,
21.5027122497559,
-13.8925476074219,
-48.9203720092773,
-44.0125236511231,
8.36602401733398,
20.6892910003662,
51.9471893310547,
0.342499256134033,
-42.1915512084961,
-11.4184761047363,
1.90410566329956,
4.09291696548462,
-4.69747734069824,
50.3577003479004,
24.6937408447266,
-4.78286552429199,
-16.1402339935303,
38.6648597717285,
11.5767726898193,
-15.6324367523193,
32.3399925231934,
-39.8878059387207,
39.7762985229492,
3.85514211654663,
-30.9772434234619,
-13.5273132324219,
-34.1361389160156,
52.7106742858887,
3.16452360153198,
1.91624593734741,
26.4321765899658,
-26.7817173004150,
-15.0954732894897,
10.2103252410889,
-24.2703399658203,
8.07615089416504,
9.04712390899658,
-56.6321945190430,
27.2459869384766,
-21.2628440856934,
-27.0722885131836,
41.5225105285645,
-75.9350585937500,
-19.1110382080078,
30.4771804809570,
-47.3823242187500,
-23.8106384277344,
-0.825186729431152,
1.11892223358154,
14.2797956466675,
-22.7141304016113,
-53.2961082458496,
-9.38124465942383,
-6.81815671920776,
-56.1252555847168,
31.3178825378418,
43.5415611267090,
-49.5114364624023,
30.6907501220703,
33.9975814819336,
25.0662937164307,
-5.85100317001343,
-38.1983795166016,
33.7448883056641,
-12.4360065460205,
55.4438972473145,
20.6879081726074,
-59.1322135925293,
18.7912178039551,
26.5280418395996,
-9.88844394683838,
-66.8519897460938,
39.1351928710938,
-14.7439117431641,
-51.9271316528320,
18.0444335937500,
-10.6758012771606,
20.4016094207764,
-13.5107402801514,
23.1684112548828,
-26.9263839721680,
-40.5872955322266,
-31.3577346801758,
18.2259941101074,
18.7399597167969,
-21.6137390136719,
43.4034996032715,
-31.4266643524170,
38.7894363403320,
24.8308181762695,
-17.6715488433838,
-19.5694503784180,
-39.5857009887695,
-32.3921508789063,
-19.1259536743164,
20.3143730163574,
-11.8694534301758,
17.7252998352051,
-47.3498001098633,
24.0132560729980,
61.2275009155273,
-25.1115779876709,
17.6764526367188,
18.1090335845947,
63.1351318359375,
-8.13861083984375,
-5.98097419738770,
63.0070877075195,
-20.5989990234375,
-53.3276863098145,
-27.4376258850098,
24.3970832824707,
-1.15742015838623,
12.1573677062988,
-9.74278640747070,
-7.10439777374268,
14.9662055969238,
-87.2063674926758,
24.3565826416016,
39.7942695617676,
-61.8549118041992,
-25.0582675933838,
2.45244312286377,
11.7839183807373,
-36.5539512634277,
34.6401214599609,
49.8074378967285,
3.01390933990479,
40.5945205688477,
-47.7149543762207,
31.6919746398926,
36.2184867858887,
-53.2389411926270,
14.5347795486450,
-21.0491447448730,
-2.64758348464966,
-37.5594253540039,
-15.5404644012451,
6.60662794113159,
-46.7907257080078,
-42.9699134826660,
-34.0779647827148,
15.0307416915894,
-44.0835952758789,
-28.2649688720703,
33.8666687011719,
40.6133041381836,
-31.6294059753418,
-2.35357427597046,
71.4649734497070,
-0.954368591308594,
-7.61533546447754,
-26.9985733032227,
-9.14769554138184,
55.2492446899414,
27.0257740020752,
-47.9072380065918,
7.32093763351440,
21.1033802032471,
-50.3957901000977,
-24.6525878906250,
28.5370960235596,
27.5203495025635,
-6.44980573654175,
-44.5827713012695,
-8.97042846679688,
59.7869110107422,
-10.1504201889038,
8.89976692199707,
1.68845987319946,
-31.9963417053223,
-21.1848831176758,
-37.4375686645508,
55.2497062683106,
12.7860527038574,
-21.8642082214355,
12.0435295104980,
18.9425716400147,
48.0180130004883,
0.534009456634522,
34.8786659240723,
-6.99900627136231,
-43.0532341003418,
41.9356269836426,
-22.3969631195068,
-10.6044397354126,
-8.08014869689941,
-51.0541572570801,
-7.48463106155396,
7.53682804107666,
42.4224624633789,
3.05381107330322,
21.1613349914551,
54.0286560058594,
21.0326824188232,
50.8441848754883,
44.5948524475098,
-33.7747421264648,
-1.27149057388306,
49.8910408020020,
-23.8883514404297,
10.6435642242432,
-26.8886642456055,
-3.29004478454590,
51.9999732971191,
-7.14716768264771,
-14.8438262939453,
-22.7004795074463,
28.9774551391602,
-9.71323490142822,
39.0456390380859,
51.3099212646484,
-9.61339473724365,
35.3505249023438,
-6.37988138198853,
34.6727371215820,
11.0245523452759,
-5.52026462554932,
49.5606918334961,
-31.4677276611328,
-40.1279678344727,
-8.70352172851563,
28.4636497497559,
-35.5024490356445,
-65.5941543579102,
31.2390003204346,
-43.6613998413086,
-18.5010814666748,
57.6946716308594,
-13.2039394378662,
23.0274620056152,
11.0469636917114,
-20.6455116271973,
-16.6197681427002,
-13.3792476654053,
53.4682540893555,
-36.3185997009277,
9.55046844482422,
22.4593505859375,
-48.5047111511231,
4.35383844375610,
-39.1687927246094,
-2.93638944625855,
31.0452041625977,
16.8985233306885,
-10.0341281890869,
-7.86785697937012,
-21.6431503295898,
30.2654800415039,
9.50450897216797,
-59.1024398803711,
-3.11155891418457,
-41.2602081298828,
20.0770492553711,
-26.2627048492432,
-24.2096939086914,
55.9247512817383,
-43.6657943725586,
-1.97161483764648,
26.7026710510254,
15.6310501098633,
26.5092678070068,
-29.9103889465332,
9.23042201995850,
56.5932044982910,
-18.9893302917480,
-2.49667263031006,
-10.7973880767822,
-31.2795867919922,
64.6301269531250,
-17.0195369720459,
-24.4146480560303,
38.6961517333984,
-23.6461982727051,
-4.15070724487305,
-9.22033882141113,
-29.9199676513672,
-31.0382614135742,
-33.2185745239258,
-43.8961639404297,
-31.2592391967773,
-37.1753616333008,
-17.7589950561523,
15.5895767211914,
-24.2431297302246,
-37.3986358642578,
-21.4300594329834,
35.0175971984863,
21.8800487518311,
8.82989692687988,
10.9392223358154,
-12.6811485290527,
13.0202465057373,
63.5125160217285,
4.61319684982300,
0.523465633392334,
52.7969894409180,
-39.7617607116699,
-4.87716817855835,
-17.3950309753418,
12.3725357055664,
45.8277473449707,
-38.0008773803711,
23.8855762481689,
22.1446418762207,
-34.5705947875977,
-22.2039756774902,
-9.44107341766357,
8.65969657897949,
29.8028469085693,
-29.8952941894531,
-22.1599159240723,
11.6085548400879,
-18.6783580780029,
-25.4769363403320,
5.05584383010864,
29.9085407257080,
-46.1193122863770,
-22.9799537658691,
11.2237224578857,
-13.2371330261230,
27.4216461181641,
-32.8647994995117,
-45.2022323608398,
3.56384134292603,
-23.5955123901367,
14.8088512420654,
-2.15087604522705,
-26.4706096649170,
10.3796129226685,
8.46541404724121,
32.4625091552734,
16.7875175476074,
-8.45784759521484,
13.1831340789795,
22.3181419372559,
-30.5844173431397,
1.14708185195923,
69.9268417358398,
-21.7081756591797,
-21.9047832489014,
27.2229385375977,
-27.2559432983398,
-6.16680669784546,
34.8495826721191,
-0.0470294952392578,
0.292368888854980,
57.2552680969238,
-15.3677692413330,
-37.6024703979492,
44.7155494689941,
19.0288314819336,
-15.7655620574951,
3.76507186889648,
42.8199768066406,
32.0399055480957,
43.4344100952148,
33.7236366271973,
47.3742408752441,
24.3839340209961,
-28.8146610260010,
-3.92350983619690,
-2.89049863815308,
53.0628852844238,
13.2981338500977,
4.40221405029297,
9.27739143371582,
-34.2233848571777,
13.3898792266846,
-20.6979560852051,
24.2327537536621,
5.82744121551514,
-25.8225650787354,
65.7671203613281,
38.2577285766602,
-11.4907855987549,
-32.6776199340820,
28.5972518920898,
21.4075679779053,
24.5589752197266,
51.3628005981445,
16.1997756958008,
48.6401939392090,
24.3335227966309,
-24.1711025238037,
-20.4998893737793,
42.2012214660645,
-6.25543308258057,
-51.1882514953613,
27.0099849700928,
32.8556442260742,
-9.33837413787842,
-13.1758308410645,
0.805379867553711,
-41.2084960937500,
-4.15886831283569,
33.0975685119629,
-43.2309608459473,
-45.0604438781738,
46.8256645202637,
8.95709037780762,
-62.0552902221680,
12.8080949783325,
-18.2095413208008,
11.2708721160889,
11.1601371765137,
-21.9239273071289,
-3.77810621261597,
-36.5328216552734,
54.5058517456055,
13.8466491699219,
19.2088813781738,
26.3752670288086,
15.5796146392822,
0.0679888725280762,
-34.0281791687012,
-0.314066886901855,
-34.1231155395508,
38.7987518310547,
28.2628173828125,
-14.2488107681274,
-33.6980857849121,
-6.14732503890991,
-35.8085098266602,
-4.20417213439941,
38.1292724609375,
-46.2824516296387,
61.5024185180664,
6.73408317565918,
12.7546501159668,
59.7215614318848,
4.26753759384155,
54.2625007629395,
3.42396020889282,
39.8398513793945,
65.7809143066406,
25.5717544555664,
38.8469085693359,
20.9368705749512,
-19.3817253112793,
-21.9028472900391,
-8.77578926086426,
-45.9875259399414,
18.5657749176025,
-17.8055057525635,
-73.7924041748047,
4.70524644851685,
-14.8700942993164,
-13.3381700515747,
-20.6083583831787,
46.7550926208496,
30.9140167236328,
-62.8532028198242,
29.5271644592285,
18.1186389923096,
9.86339187622070,
26.8461570739746,
38.9621658325195,
36.6249198913574,
7.88479089736939,
29.5786399841309,
15.8591709136963,
56.3017501831055,
21.9300575256348,
-20.8545780181885,
15.2188110351563,
16.1052780151367,
-38.9250221252441,
-11.7561826705933,
61.2561416625977,
-28.7618961334229,
-34.4801902770996,
7.39750576019287,
-25.2972183227539,
22.1223163604736,
23.4046802520752,
-47.0649833679199,
-10.0262126922607,
23.2801990509033,
-9.89751911163330,
9.24390697479248,
-21.2311363220215,
-29.5388908386230,
33.7722396850586,
31.0546417236328,
31.2849826812744,
-19.8207569122314,
-49.2542953491211,
13.1771240234375,
43.9225959777832,
18.3301658630371,
-5.15068054199219,
21.6396121978760,
16.4076423645020,
16.2440872192383,
37.5250358581543,
52.2700805664063,
10.2126464843750,
19.6988639831543,
51.3362998962402,
-24.5219497680664,
7.94507980346680,
49.0618820190430,
14.0151176452637,
-76.1333007812500,
-1.98897886276245,
42.6271209716797,
-52.6775360107422,
45.8235054016113,
-6.40202045440674,
11.4800643920898,
42.3016815185547,
9.09166622161865,
62.0827636718750,
11.9554023742676,
-39.1740646362305,
4.70302772521973,
39.3484191894531,
-50.2016143798828,
38.2790336608887,
46.4401168823242,
-19.7903861999512,
17.3950004577637,
61.5444526672363,
-6.46375036239624,
-32.1341133117676,
15.3001708984375,
-34.0783081054688,
48.9490737915039,
-48.2209281921387,
-31.0624771118164,
40.2488555908203,
-56.8356399536133,
-8.12390613555908,
6.16263484954834,
12.0480127334595,
3.80852413177490,
-32.5181465148926,
13.0853500366211,
-0.925311088562012,
-13.6812982559204,
37.5094070434570,
34.5597114562988,
46.3128776550293,
14.7790842056274,
14.4409122467041,
-47.1732101440430,
11.1927165985107,
46.7532348632813,
-52.9229698181152,
20.5108871459961,
1.34605598449707,
32.5775451660156,
-19.7996120452881,
-17.4512634277344,
15.5607280731201,
-43.0647544860840,
-10.4250192642212,
-37.4140853881836,
75.9018249511719,
14.6226902008057,
-47.0540161132813,
35.7398757934570,
-17.9762229919434,
-15.9345378875732,
-38.9021301269531,
-14.1559123992920,
-8.04369735717773,
-13.1925668716431,
48.6198120117188,
-9.50834083557129,
47.9465675354004,
39.7995300292969,
-38.2754440307617,
52.1286048889160,
21.3213195800781,
-10.1888103485107,
-33.2182044982910,
-5.04824352264404,
45.1144027709961,
29.2063941955566,
26.1960830688477,
-51.3884162902832,
-13.2330017089844,
27.0253410339355,
-14.2386531829834,
-28.1694717407227,
-35.5251464843750,
-34.2136764526367,
-21.3734703063965,
47.4935111999512,
-5.15523004531860,
-41.7225799560547,
39.4843864440918,
-16.5238227844238,
13.2541046142578,
54.2719993591309,
-40.6313781738281,
11.1623497009277,
64.7198715209961,
5.47206020355225,
-17.4175491333008,
12.0618915557861,
54.3176574707031,
1.62423133850098,
20.1930999755859,
64.5548858642578,
-16.4021911621094,
-19.8337764739990,
-29.3266429901123,
-2.73618507385254,
-11.4717302322388,
-20.6098461151123,
4.58509969711304,
22.5231723785400,
12.4695930480957,
-44.9797668457031,
18.7574863433838,
6.68022155761719,
36.5414047241211,
-19.2220630645752,
-30.0326995849609,
41.4063415527344,
-51.2424507141113,
27.4157924652100,
42.8966941833496,
11.2559833526611,
12.0947847366333,
-6.37993288040161,
48.4624252319336,
47.2663345336914,
15.6517963409424,
-35.3465843200684,
-16.8320007324219,
-17.3662471771240,
-38.0841522216797,
-12.6479091644287,
43.3766784667969,
28.4736480712891,
-47.6688537597656,
46.3197593688965,
-0.185464859008789,
-39.4209594726563,
59.5301628112793,
10.7363338470459,
-50.7121696472168,
41.2884292602539,
35.7016525268555,
-1.04582118988037,
39.2520561218262,
-8.08052158355713,
31.0021305084229,
-15.2419862747192,
11.0243015289307,
64.5144042968750,
37.2941284179688,
-11.8427238464355,
-16.0925941467285,
59.6080245971680,
-56.8361663818359,
-16.4963645935059,
29.3742923736572,
-6.11082077026367,
17.4148178100586,
-20.0273704528809,
-4.98755693435669,
21.4134292602539,
-16.3227252960205,
-41.3342056274414,
3.04554176330566,
-39.9227676391602,
1.98008489608765,
48.0355606079102,
2.07586908340454,
40.0643157958984,
-22.7130832672119,
-32.1034164428711,
16.6387481689453,
-14.4323453903198,
-41.7625198364258,
-19.9926109313965,
49.0287170410156,
-51.5661277770996,
-49.6603355407715,
69.6712493896484,
-17.1182060241699,
-29.6363658905029,
-1.81742858886719,
21.7975044250488,
5.42721080780029,
-57.3092460632324,
71.8614425659180,
28.2176742553711,
-58.1630249023438,
-10.6046895980835,
-41.7563934326172,
15.2837982177734,
6.14728355407715,
-30.9884033203125,
-25.0880165100098,
1.42479419708252,
-24.6040191650391,
-16.5609874725342,
40.5819358825684,
-19.6263084411621,
19.5878620147705,
-43.0681610107422,
11.7174301147461,
98.5818634033203,
-47.5026168823242,
-6.37164211273193,
29.7026901245117,
-53.3760185241699,
-31.6592617034912,
-8.67560195922852,
-53.1568565368652,
-6.95529079437256,
-0.299249649047852,
-18.0214958190918,
35.1793365478516,
22.5949325561523,
-12.4754219055176,
2.71886396408081,
-10.0811347961426,
-21.6976280212402,
-21.6008453369141,
-40.0724067687988,
-7.18496990203857,
-29.1534538269043,
-5.54240369796753,
33.7320671081543,
-15.2133865356445,
24.9740104675293,
41.5305290222168,
-29.8197116851807,
-6.06472206115723,
-20.1015663146973,
-14.6315059661865,
14.1961345672607,
-49.4801025390625,
16.7249832153320,
-7.81098079681397,
-7.62964916229248,
5.71773624420166,
-58.1804656982422,
-35.9108390808106,
-10.3277282714844,
48.0643234252930,
-7.95264148712158,
-37.1985206604004,
-6.86313915252686,
-24.9611167907715,
-13.9361400604248,
35.4310951232910,
3.09795904159546,
-12.1414394378662,
33.4026451110840,
9.67759704589844,
-20.1346340179443,
-18.6021270751953,
-8.40657711029053,
-27.5967445373535,
18.0679740905762,
-14.4968357086182,
-36.3455162048340,
-40.4999389648438,
-35.5268478393555,
-26.7935924530029,
-25.8787117004395,
15.5870323181152,
-30.8959941864014,
5.13877630233765,
-24.9544372558594,
4.84076595306397,
57.4897575378418,
6.92822360992432,
-35.8723945617676,
-12.7640380859375,
17.5401554107666,
-56.9007949829102,
-27.3299751281738,
9.36224269866943,
33.3498077392578,
23.3061046600342,
-8.79641246795654,
-32.3880577087402,
27.8073444366455,
24.9176120758057,
11.8508615493774,
16.8760375976563,
-24.2799930572510,
50.8650436401367,
-47.1147232055664,
-44.3409156799316,
18.6212158203125,
6.95335531234741,
19.1573104858398,
-0.554143428802490,
67.7060089111328,
11.2506237030029,
-36.4883613586426,
44.8388404846191,
-2.62719678878784,
-48.4691696166992,
55.3773689270020,
-0.465684890747070,
-63.2390632629395,
56.2335090637207,
13.1968221664429,
-48.1610221862793,
10.5023078918457,
29.9513320922852,
-38.4358482360840,
-15.2277927398682,
53.4018478393555,
-58.1630477905273,
-27.1899757385254,
52.7633247375488,
-2.02761411666870,
-31.1198368072510,
-53.9704322814941,
14.1745147705078,
27.0824050903320,
-87.6445999145508,
-20.1082534790039,
15.8860950469971,
-23.7336139678955,
30.4557456970215,
-21.4020748138428,
4.27138090133667,
11.0449371337891,
7.48690891265869,
32.2911949157715,
32.0082588195801,
40.4130859375000,
-37.7635269165039,
45.0663528442383,
61.1664581298828,
-1.51521015167236,
-0.733207702636719,
-17.2326393127441,
-1.64041709899902,
-6.19749546051025,
39.8694953918457,
13.0881271362305,
0.935502529144287,
33.7979431152344,
-36.1881675720215,
-7.94766569137573,
60.4669837951660,
39.5116310119629,
5.90334224700928,
-18.5674705505371,
37.5641021728516,
37.8538436889648,
-27.1323585510254,
11.7905921936035,
-29.0037231445313,
-34.5386848449707,
36.7678184509277,
22.5185203552246,
-14.1968698501587,
-20.4893589019775,
43.1969604492188,
-21.9002609252930,
-28.7991523742676,
86.5288925170898,
18.2467842102051,
-42.0897216796875,
3.42907905578613,
40.8832702636719,
3.97583580017090,
12.0353775024414,
58.7305145263672,
35.2298965454102,
11.4085826873779,
2.39553499221802,
-24.2529182434082,
-38.3829727172852,
-12.3168344497681,
14.0837469100952,
27.0594444274902,
-23.9830493927002,
17.6190090179443,
21.2975540161133,
-53.7950820922852,
-18.5301227569580,
9.36347579956055,
61.7363166809082,
9.36477565765381,
-35.8069839477539,
32.3986091613770,
-22.0739974975586,
25.2779197692871,
71.0324554443359,
-14.5295257568359,
24.5056877136230,
6.75228691101074,
11.8852081298828,
17.1704273223877,
-17.6391563415527,
29.9453430175781,
-35.8778114318848,
-25.4124794006348,
40.4077453613281,
43.0718460083008,
-17.8149414062500,
-57.8639488220215,
15.5047531127930,
-18.5603561401367,
-13.9526481628418,
-22.3085994720459,
-38.3584747314453,
-26.0882911682129,
-19.4522590637207,
46.5340080261231,
-25.4378890991211,
23.8155574798584,
21.9226303100586,
-41.7904090881348,
23.3151721954346,
30.8244018554688,
18.5868644714355,
-54.3829345703125,
-0.268142700195313,
-15.4126272201538,
-54.0251502990723,
14.2065925598145,
-2.48958063125610,
15.2062005996704,
-23.5371780395508,
-34.9936141967773,
-14.6371507644653,
-15.6867637634277,
20.9150581359863,
-1.20597028732300,
-21.1087131500244,
-9.41563987731934,
24.4520435333252,
17.9328956604004,
31.0535964965820,
46.5030479431152,
-10.1802597045898,
26.9565868377686,
56.9288024902344,
7.01039791107178,
-38.2901802062988,
37.6625175476074,
41.8768501281738,
-59.7248687744141,
38.8080368041992,
25.1950187683105,
-36.9318771362305,
30.8263359069824,
8.15415573120117,
33.7158050537109,
37.4935493469238,
32.4838104248047,
-14.3175582885742,
-45.2610740661621,
61.4221458435059,
38.2694168090820,
31.8451175689697,
-16.8869895935059,
-17.3679790496826,
48.2121963500977,
42.4556884765625,
36.4232864379883,
8.62324714660645,
26.3889617919922,
-39.5147933959961,
20.5107326507568,
40.5297622680664,
2.65827989578247,
36.4995040893555,
-57.8201446533203,
-5.11049079895020,
24.4703140258789,
-51.9682235717773,
36.6309928894043,
14.2963962554932,
-69.4177322387695,
44.7285728454590,
24.6999740600586,
10.0680332183838,
33.5717773437500,
-40.5286941528320,
13.4921789169312,
38.5093116760254,
13.3875389099121,
-16.3734207153320,
-23.1662216186523,
25.1623573303223,
47.3170242309570,
-21.3894386291504,
6.54060649871826,
53.8745346069336,
-36.8362197875977,
12.7225055694580,
65.6280136108398,
37.4972915649414,
21.6474075317383,
-28.6243515014648,
-10.9073333740234,
49.1508674621582,
16.9074134826660,
20.0117530822754,
58.2264709472656,
25.5497589111328,
-15.6868133544922,
-23.4777679443359,
65.0831832885742,
39.5472183227539,
-49.2849693298340,
51.6949462890625,
10.2834520339966,
-50.1686592102051,
49.5844192504883,
14.2328948974609,
-4.89376544952393,
4.28713035583496,
0.0187573432922363,
4.13229227066040,
-42.6221389770508,
-2.35123634338379,
17.6229782104492,
-40.5036125183106,
-33.7781639099121,
-8.93158245086670,
-25.2160949707031,
-31.0382232666016,
23.9017276763916,
25.1857452392578,
6.42375040054321,
26.2624092102051,
-39.9398612976074,
-34.1078033447266,
10.3548069000244,
27.4095954895020,
40.4275398254395,
-37.5361137390137,
-4.63256549835205,
40.6555252075195,
19.2487449645996,
43.3595008850098,
-23.2753829956055,
-16.4315090179443,
21.7610054016113,
-28.0595207214355,
10.6252460479736,
-2.54181241989136,
-45.8305931091309,
-33.5397567749023,
-25.2105865478516,
-31.5187397003174,
-44.0525093078613,
-31.1161918640137,
-27.8597335815430,
-44.5570220947266,
9.32817077636719,
51.9599418640137,
-40.0665626525879,
-0.382502079010010,
47.4631309509277,
10.8004322052002,
9.07928085327148,
27.3322696685791,
52.0558166503906,
11.0067119598389,
29.9321537017822,
2.92401075363159,
-17.9922084808350,
-14.6030235290527,
33.2173271179199,
10.4217271804810,
-69.4084014892578,
-14.2089385986328,
-23.1302413940430,
32.9645042419434,
13.8793106079102,
-10.9448013305664,
41.2799415588379,
-10.1431760787964,
-5.16372489929199,
44.1420249938965,
18.9818782806397,
-46.7173347473145,
-7.55927848815918,
63.9680328369141,
23.8078899383545,
-32.7065086364746,
17.2666835784912,
0.790376663208008,
-11.1952152252197,
20.6677398681641,
15.8340435028076,
48.7120323181152,
2.61817836761475,
-2.57426118850708,
34.4204597473145,
18.3252449035645,
23.0188274383545,
-11.4773731231689,
-28.1810913085938,
0.111776828765869,
24.7737960815430,
17.7411804199219,
2.28440809249878,
50.2607040405273,
6.43932914733887,
-53.0051383972168,
41.5905876159668,
53.2642135620117,
-46.6554756164551,
35.0754203796387,
16.4264526367188,
-58.0102462768555,
69.4769287109375,
-8.89085578918457,
-28.0989837646484,
76.4503631591797,
21.0516929626465,
-50.4165802001953,
21.5662899017334,
70.7067642211914,
-57.5607681274414,
19.2616767883301,
52.7086105346680,
-39.9799842834473,
-55.9226074218750,
0.889037609100342,
43.9595489501953,
-47.6338653564453,
19.0246047973633,
31.5060462951660,
-14.3852777481079,
7.28664922714233,
33.7678375244141,
25.8786544799805,
-55.3821716308594,
-5.75068426132202,
33.0670242309570,
4.62010765075684,
0.889649391174316,
18.6670589447022,
-11.5940132141113,
7.21441698074341,
13.3643875122070,
-9.20310211181641,
61.0193710327148,
-30.7879161834717,
-17.8397369384766,
64.5554504394531,
7.65601921081543,
-0.148579597473145,
9.81209754943848,
52.5660629272461,
-19.3865432739258,
-22.9547309875488,
53.4895935058594,
-25.1478691101074,
-72.8150024414063,
9.44235420227051,
29.3024406433105,
-14.1883258819580,
25.6283664703369,
-19.6187763214111,
-17.0905838012695,
23.9027462005615,
25.4267501831055,
47.1722412109375,
30.9783058166504,
45.9187545776367,
41.7287101745606,
16.0978775024414,
39.1703758239746,
32.9520759582520,
-45.6279525756836,
16.0575695037842,
59.3861122131348,
-38.0911178588867,
1.38741016387939,
13.2035560607910,
-45.6674194335938,
-23.0969200134277,
-10.6845140457153,
-25.6126289367676,
-20.2589569091797,
6.67855310440064,
32.0676307678223,
-17.1721210479736,
-50.7949485778809,
31.5125885009766,
-12.7577781677246,
-27.1216926574707,
11.5653476715088,
-37.4094772338867,
6.15434360504150,
57.1978416442871,
18.0011157989502,
-44.5034713745117,
6.97567462921143,
-13.8925151824951,
-31.0420494079590,
-6.03050518035889,
-65.9484634399414,
-5.65599966049194,
7.55092811584473,
-24.7936878204346,
12.5530529022217,
9.74153041839600,
16.3463211059570,
-7.64665174484253,
-30.1821556091309,
-4.22345542907715,
-49.8604431152344,
-1.23247861862183,
63.0297317504883,
6.08900880813599,
-23.2639541625977,
11.3337001800537,
6.87240219116211,
-43.2653274536133,
-2.70871019363403,
41.7168922424316,
43.5171813964844,
-22.0832290649414,
-40.9916419982910,
9.16827964782715,
32.6640548706055,
-24.8774871826172,
-29.3658676147461,
25.9687137603760,
-3.35489892959595,
19.0127372741699,
-35.5941848754883,
-13.7361640930176,
16.6530075073242,
5.44306516647339,
5.23279142379761,
-14.0247688293457,
57.8714408874512,
-7.99586772918701,
11.5271911621094,
21.2535533905029,
-6.45946168899536,
-9.40654850006104,
-28.2910652160645,
71.1025619506836,
-13.4208173751831,
0.891734123229981,
39.6784057617188,
-35.5287246704102,
21.0283374786377,
45.6380844116211,
44.4493255615234,
-18.3813209533691,
7.89864253997803,
13.0284957885742,
-65.2664184570313,
26.0130176544189,
69.5025939941406,
17.6702136993408,
-15.1407699584961,
-21.5672092437744,
-22.9528121948242,
3.90509700775147,
31.9335289001465,
16.4410552978516,
4.36264085769653,
4.76706981658936,
5.28293037414551,
-33.1047248840332,
-0.814669132232666,
33.1274795532227,
-15.8981904983521,
8.84728145599365,
51.5634613037109,
-14.4498767852783,
-28.4954071044922,
42.6048583984375,
-12.2585868835449,
-50.2406158447266,
24.9973716735840,
57.6032676696777,
6.46642589569092,
-55.8173065185547,
-10.0310811996460,
1.80885171890259,
12.7566051483154,
47.7276611328125,
-0.528759956359863,
26.2188663482666,
-22.0033435821533,
-34.0535850524902,
0.572644233703613,
-9.89624977111816,
58.4730529785156,
-27.2423133850098,
-37.2417831420898,
17.1226310729980,
-22.2167091369629,
37.8922042846680,
-8.32101726531982,
-59.0311317443848,
37.1724853515625,
18.7031497955322,
-57.4560928344727,
-21.8856239318848,
53.2534484863281,
-2.94888734817505,
-69.3637695312500,
20.3719215393066,
11.3077201843262,
-28.5197563171387,
32.5505599975586,
-12.7019462585449,
-52.3333740234375,
5.63363933563232,
-51.1950721740723,
-38.1461143493652,
26.7419147491455,
-30.1076831817627,
19.5709877014160,
13.7363624572754,
26.3275909423828,
15.5286273956299,
-60.3724403381348,
47.7726020812988,
0.434963226318359,
-29.9039077758789,
60.7501602172852,
10.6086683273315,
-37.6212234497070,
-39.2698669433594,
8.98032379150391,
40.5448989868164,
-0.718043327331543,
-41.1006126403809,
29.8223686218262,
16.9168262481689,
-44.6751899719238,
32.0636596679688,
45.3318557739258,
6.47424650192261,
-45.9895553588867,
3.47061586380005,
69.4831695556641,
21.7199134826660,
32.1373977661133,
15.9730281829834,
-53.3403015136719,
-19.1678543090820,
66.7883605957031,
-7.71991872787476,
-24.4416084289551,
37.2317581176758,
-34.6086845397949,
-39.5981025695801,
19.6344604492188,
56.5875587463379,
16.9836330413818,
-9.10451507568359,
22.0734157562256,
41.3001365661621,
42.4484405517578,
25.2868309020996,
-0.134395122528076,
-4.12115716934204,
23.2960948944092,
-37.0827445983887,
27.7588729858398,
2.67903137207031,
-21.9996089935303,
26.0690689086914,
-50.1342277526856,
33.1977767944336,
-25.0179424285889,
18.5997905731201,
74.9204711914063,
-7.31087350845337,
40.6671943664551,
-3.16035699844360,
-16.8841342926025,
3.79709386825562,
52.5767822265625,
-24.8553123474121,
-52.6002807617188,
3.11347103118897,
-43.0852584838867,
23.9502372741699,
16.3890151977539,
11.1214628219605,
14.4570598602295,
-37.2049293518066,
-30.3285942077637,
39.2926254272461,
35.9681587219238,
-62.5352935791016,
-16.7975120544434,
33.9239501953125,
51.9204635620117,
-3.02690362930298,
-19.6357479095459,
-4.88699054718018,
-22.0500640869141,
29.7257308959961,
-6.63202857971191,
50.3014602661133,
10.3213310241699,
-53.0289840698242,
21.7762069702148,
-26.8225631713867,
7.90130758285523,
63.1805686950684,
-0.613126754760742,
-28.4556846618652,
-17.6557006835938,
4.06397438049316,
17.6508674621582,
-46.6198806762695,
-32.3979644775391,
13.1545867919922,
14.6827907562256,
44.4145431518555,
-13.7439842224121,
-4.73622846603394,
-12.7531251907349,
-35.6082611083984,
44.4732627868652,
-36.2458190917969,
-30.8932228088379,
43.8026428222656,
-21.4330844879150,
0.527321815490723,
25.0436935424805,
-4.94273805618286,
-32.3107490539551,
-24.4701805114746,
-6.74746227264404,
11.4457578659058,
37.2914619445801,
5.06773853302002,
29.6539306640625,
28.6393241882324,
-38.5433158874512,
-20.1011962890625,
30.6804313659668,
41.0505409240723,
4.71977329254150,
-22.4622955322266,
2.09246349334717,
27.6484298706055,
17.6184959411621,
-0.599109649658203,
10.9837770462036,
-6.33096694946289,
-50.3346939086914,
-10.1081638336182,
51.8954849243164,
0.393292427062988,
-53.0770263671875,
47.6105384826660,
9.79182147979736,
-54.5974578857422,
45.8387069702148,
-9.01051139831543,
0.314754486083984,
22.3408241271973,
-24.0396423339844,
14.0418653488159,
-20.2675590515137,
-34.3817749023438,
-9.52806091308594,
-38.0233154296875,
-53.1007499694824,
-41.9425773620606,
-51.5772094726563,
-24.6863594055176,
-12.4997920989990,
18.1761360168457,
-15.7569599151611,
-30.3770179748535,
59.0762100219727,
-1.95362329483032,
12.1461286544800,
53.8360023498535,
-19.1121902465820,
25.3345298767090,
78.1813964843750,
-8.68816471099854,
18.4366989135742,
55.7998733520508,
-29.1034622192383,
-27.1940555572510,
15.6831636428833,
4.22820568084717,
-52.9396057128906,
2.32575893402100,
4.88258171081543,
-27.8775329589844,
13.9908323287964,
-38.1021270751953,
-1.59970569610596,
6.67403221130371,
-36.1678237915039,
19.8677597045898,
5.10957813262939,
2.81553745269775,
46.0057220458984,
43.0113945007324,
29.3274841308594,
-7.91737604141235,
-57.9612579345703,
15.9173240661621,
33.2495307922363,
-58.6374359130859,
-33.9560852050781,
4.64674568176270,
-4.87698078155518,
32.7082672119141,
15.0211172103882,
-51.0415382385254,
31.1813812255859,
35.6212768554688,
29.0994300842285,
-4.53178787231445,
-23.7060737609863,
24.1422042846680,
-39.9645004272461,
24.3035297393799,
10.2997579574585,
-50.9996185302734,
-42.3297195434570,
17.3177528381348,
-6.62361049652100,
-35.8988113403320,
26.7267684936523,
-3.10516405105591,
-10.5314683914185,
-42.8422470092773,
-13.3842983245850,
-25.8144683837891,
7.15357875823975,
8.49670219421387,
-42.6158943176270,
2.86555194854736,
-39.1716117858887,
20.4356155395508,
39.8243255615234,
9.36943054199219,
8.15540981292725,
31.4118766784668,
46.2276611328125,
-28.6577167510986,
-18.2912025451660,
-13.2638988494873,
0.926767349243164,
-39.3979339599609,
-7.76006698608398,
23.0129356384277,
-62.6327095031738,
-18.0163230895996,
-14.1817684173584,
-55.0494537353516,
-31.7796401977539,
44.2515335083008,
7.83386993408203,
38.6922950744629,
1.84531879425049,
-19.1069927215576,
15.6475229263306,
-40.1683692932129,
36.1143455505371,
-22.9476280212402,
19.5470352172852,
-23.0276584625244,
-13.7916669845581,
28.8677749633789,
-34.9343795776367,
50.4072570800781,
12.1672077178955,
-12.5367689132690,
-47.8373641967773,
1.02100944519043,
26.5472412109375,
-1.35364294052124,
35.5105438232422,
37.6878814697266,
-29.7177391052246,
-10.3586263656616,
85.8095245361328,
-8.84174346923828,
-7.17669677734375,
62.3398818969727,
40.7859954833984,
15.8140182495117,
-4.38379287719727,
-25.4682712554932,
7.09659385681152,
19.5698013305664,
-16.0871505737305,
28.9989967346191,
31.2003040313721,
1.59824466705322,
-42.7152976989746,
-3.73124504089355,
31.4076900482178,
-44.0461883544922,
19.2929458618164,
13.7013177871704,
-48.7571754455566,
-16.8505592346191,
25.0774726867676,
10.2678775787354,
-49.6767196655273,
20.5321102142334,
52.9887619018555,
11.3449783325195,
-22.0455741882324,
15.4275751113892,
35.9905319213867,
7.21602153778076,
60.6409034729004,
17.5708084106445,
-27.0071620941162,
37.2602233886719,
40.1949729919434,
-40.2481651306152,
-22.7841892242432,
50.8070602416992,
29.5699443817139,
7.15863132476807,
30.2467269897461,
10.3595151901245,
-14.8774566650391,
-9.37944507598877,
3.63921260833740,
14.7619667053223,
-35.5970611572266,
-30.1395416259766,
36.2892684936523,
-2.01956701278687,
-5.42858123779297,
-4.35179805755615,
-17.4436397552490,
76.4575500488281,
-13.8718585968018,
-35.0080299377441,
47.6843605041504,
-55.0430564880371,
-47.8252258300781,
-25.9992980957031,
7.77806377410889,
30.9599685668945,
-49.4242057800293,
-36.5157432556152,
7.11898994445801,
-5.12187290191650,
-33.7061119079590,
-37.8315925598145,
3.52166652679443,
16.5498046875000,
-43.6307716369629,
-30.0463256835938,
2.21140289306641,
21.4442443847656,
7.14500904083252,
-45.6797294616699,
37.9668159484863,
39.7523002624512,
26.1178302764893,
14.9276990890503,
-0.0664672851562500,
42.8892860412598,
-39.9386253356934,
22.9583759307861,
19.7583923339844,
-53.7526245117188,
-17.3297004699707,
-59.2186813354492,
-35.5208015441895,
28.3047485351563,
33.0926895141602,
6.19728851318359,
25.5239391326904,
20.6941986083984,
13.8667106628418,
27.5855865478516,
30.1739997863770,
-23.3332481384277,
-25.2949142456055,
77.5649108886719,
39.5103225708008,
21.2854423522949,
5.42291831970215,
-38.1621360778809,
41.7908515930176,
32.7397994995117,
-49.3375205993652,
29.2792472839355,
36.5759201049805,
-24.6490058898926,
3.43366622924805,
-23.3127403259277,
-9.63962745666504,
-32.6450271606445,
3.30448722839355,
12.1698398590088,
-61.6507644653320,
31.4954013824463,
-12.2418165206909,
-37.3400001525879,
40.3891639709473,
-37.3311462402344,
-47.4054145812988,
-44.7967910766602,
-45.0838088989258,
26.2434539794922,
34.4711303710938,
8.36512756347656,
-36.8932418823242,
-31.3670959472656,
3.58864974975586,
12.4079990386963,
-0.00235176086425781,
50.5739288330078,
-3.21143627166748,
-45.4262008666992,
54.4252548217773,
-21.6774101257324,
20.5735511779785,
48.4429931640625,
23.4926452636719,
17.0288028717041,
-20.7027473449707,
38.0639762878418,
3.14247798919678,
-54.1596832275391,
-32.8895072937012,
46.1307029724121,
-48.3927650451660,
-15.8106384277344,
24.5508079528809,
-34.4511108398438,
63.5393676757813,
-41.0726470947266,
18.3177566528320,
23.9000720977783,
-45.1086273193359,
22.7697334289551,
-49.2460365295410,
31.1227645874023,
29.5631847381592,
10.6710920333862,
-5.70492696762085,
-23.4652938842773,
27.1884078979492,
-33.5705261230469,
13.2920904159546,
3.39516353607178,
-19.5062217712402,
-33.9505538940430,
-25.4606647491455,
-17.6230812072754,
-45.3745994567871,
25.6210403442383,
-40.1834983825684,
-44.3781051635742,
-34.1953964233398,
-41.4518852233887,
-20.4195671081543,
-5.60594558715820,
22.2880516052246,
-45.4873504638672,
31.3795127868652,
1.84367942810059,
8.82327365875244,
8.97566795349121,
-37.6297912597656,
32.6458587646484,
-41.3040428161621,
44.1148223876953,
49.9395027160645,
-16.7749176025391,
-13.3138656616211,
15.9543638229370,
11.8812036514282,
-71.7293624877930,
35.0151557922363,
36.0002326965332,
-59.5526771545410,
-20.9621181488037,
-39.2174224853516,
-20.2970542907715,
37.1383972167969,
-38.1201896667481,
-15.2169733047485,
-24.8987579345703,
-6.22688388824463,
14.7325716018677,
-22.5979652404785,
43.5670967102051,
-25.5383491516113,
-2.08205986022949,
25.1279544830322,
-37.6061859130859,
-11.6153297424316,
-23.3018074035645,
-25.1210918426514,
30.0294570922852,
-5.43180370330811,
-52.2542572021484,
18.1028671264648,
-1.89351177215576,
-30.0784244537354,
28.4667816162109,
-2.86203098297119,
-4.42583847045898,
47.1893005371094,
-5.73298835754395,
8.19828510284424,
2.20740985870361,
-31.8525199890137,
14.5245122909546,
-34.3624801635742,
-5.98976993560791,
13.4552488327026,
-24.7502937316895,
28.8865203857422,
44.9040908813477,
14.8135194778442,
-4.86441469192505,
32.9962692260742,
3.44103240966797,
-30.8009681701660,
-6.52193069458008,
-34.2255401611328,
-15.4640665054321,
-39.8454322814941,
-37.3208389282227,
51.1349182128906,
-14.9393424987793,
-46.9390602111816,
41.3695449829102,
-14.0181694030762,
-43.7618675231934,
41.3705520629883,
26.8855590820313,
23.4849834442139,
7.82206344604492,
0.557456016540527,
44.5947189331055,
-18.0102157592773,
-25.3455848693848,
7.78180313110352,
1.58815574645996,
12.9981555938721,
-24.3483276367188,
-13.1838989257813,
-20.8834762573242,
-54.4084892272949,
-36.0280227661133,
-19.3213481903076,
21.3501319885254,
-53.7352371215820,
-12.7078046798706,
27.7555389404297,
-66.0839080810547,
-7.01119899749756,
7.67252063751221,
17.8898010253906,
39.8224487304688,
21.7671585083008,
-10.5728864669800,
-1.63913106918335,
9.17467975616455,
-25.1784362792969,
35.4863624572754,
34.8848838806152,
-53.9636230468750,
16.6759262084961,
36.7802391052246,
-44.1612358093262,
20.2362937927246,
-17.7083034515381,
-20.9708213806152,
-18.1482200622559,
-21.0450420379639,
29.0929145812988,
10.4812364578247,
15.3771753311157,
-30.2703781127930,
34.0851135253906,
30.5482616424561,
-8.39389991760254,
-20.8508014678955,
-43.3118438720703,
14.6373777389526,
-33.9190368652344,
-36.8115005493164,
32.9774627685547,
23.4549922943115,
-40.0305976867676,
-35.6268043518066,
18.5129127502441,
44.0875625610352,
-13.3014059066772,
-9.42436790466309,
57.1164093017578,
0.583876609802246,
-0.874776840209961,
-47.6739730834961,
-2.72324943542480,
28.0859107971191,
-65.5466156005859,
26.6366157531738,
-24.4875354766846,
-21.8366088867188,
25.4455318450928,
-31.7437438964844,
13.7701807022095,
22.6568603515625,
20.7590141296387,
-2.55112648010254,
-31.8050079345703,
-29.6893959045410,
31.4081459045410,
-6.07334089279175,
-48.9857025146484,
7.28969669342041,
-7.06457471847534,
-5.73938655853272,
8.82710075378418,
-10.0515794754028,
-38.2047462463379,
-45.1479682922363,
-42.5935707092285,
25.3185920715332,
0.568349838256836,
-18.9240264892578,
75.2787017822266,
-30.6939659118652,
-32.1293792724609,
44.8505401611328,
-59.6641769409180,
-19.3779029846191,
38.9187774658203,
2.67584133148193,
26.7968044281006,
-8.17900657653809,
-50.0745239257813,
-6.99319314956665,
-3.46232128143311,
-5.48198890686035,
58.6285858154297,
13.4154815673828,
-13.1576366424561,
61.1516838073731,
8.70227718353272,
-18.4900341033936,
6.21275520324707,
7.21029758453369,
34.9256668090820,
-26.0670604705811,
-33.9415969848633,
47.6660957336426,
-2.47305870056152,
-35.2575531005859,
-18.8305721282959,
-13.5888614654541,
-5.67921829223633,
-41.3709526062012,
-8.77954673767090,
43.5260124206543,
-24.4682979583740,
-58.9299240112305,
56.7248344421387,
7.73849391937256,
-40.7853965759277,
33.4562072753906,
24.3174743652344,
14.3363447189331,
-18.8102760314941,
31.4437637329102,
38.6302719116211,
46.0174751281738,
-10.4997320175171,
-24.0933189392090,
26.8924541473389,
-43.7503128051758,
0.289740562438965,
-15.1420125961304,
34.6220550537109,
28.3111267089844,
-6.15793561935425,
13.9007635116577,
10.7168560028076,
34.4284896850586,
-13.8300418853760,
12.6839885711670,
11.8348274230957,
10.4363489151001,
-17.7574825286865,
42.5878181457520,
36.7710342407227,
-29.3900718688965,
49.0789375305176,
-2.55816316604614,
2.62481021881104,
-7.46742820739746,
10.4460878372192,
1.96980953216553,
-42.7617568969727,
35.7672233581543,
-11.1236934661865,
25.0143108367920,
-14.8535985946655,
-46.3467178344727,
-0.0652608871459961,
-35.1393852233887,
-11.9227371215820,
-21.2763977050781,
-21.8331604003906,
-3.03396558761597,
-0.648702621459961,
-56.0302963256836,
25.9614639282227,
63.6347236633301,
-25.8577861785889,
-55.1608161926270,
32.8352127075195,
33.3918876647949,
-30.1653938293457,
51.8122444152832,
-18.6186332702637,
-52.4429855346680,
-17.1930122375488,
32.5638961791992,
-25.2638893127441,
-26.8526763916016,
30.3320198059082,
-60.0643768310547,
-3.95502567291260,
10.6301012039185,
16.6616878509522,
19.1403427124023,
-16.1843299865723,
38.9515724182129,
40.7080192565918,
-3.16908168792725,
45.7612915039063,
24.7247886657715,
-31.8438072204590,
55.1734046936035,
8.16859531402588,
-22.3113746643066,
61.9913902282715,
14.5520830154419,
30.6274795532227,
42.8487739562988,
5.16195201873779,
46.9987716674805,
37.8163909912109,
-15.6578683853149,
-18.2125778198242,
45.4884490966797,
12.7172880172730,
13.2423686981201,
28.4201736450195,
-27.8668766021729,
26.3005409240723,
-25.6406116485596,
-0.521545410156250,
64.8110046386719,
24.4816856384277,
36.8108978271484,
-3.32914733886719,
0.336448669433594,
24.3209609985352,
-3.92130851745605,
-46.9674949645996,
28.7362594604492,
45.3379898071289,
-37.7684097290039,
-23.9729499816895,
-18.6957015991211,
-25.1831398010254,
-7.51177406311035,
25.3536415100098,
-23.3194160461426,
2.37340545654297,
6.24056339263916,
-56.6779594421387,
17.6190662384033,
-1.79388999938965,
-19.8117065429688,
-1.51960372924805,
2.14553356170654,
30.1391906738281,
-6.33867073059082,
-21.0619125366211,
-37.0273437500000,
-10.8474969863892,
-0.439159393310547,
4.63956928253174,
42.5816574096680,
17.2392082214355,
-31.7381973266602,
-31.5859069824219,
-9.45219612121582,
-11.1977767944336,
42.2179565429688,
42.0447158813477,
34.9050254821777,
-2.77889919281006,
-44.7130355834961,
16.3914413452148,
26.1722507476807,
8.21035480499268,
27.5483016967773,
39.7444305419922,
-1.99260377883911,
30.6605148315430,
44.1692619323731,
-42.1230316162109,
13.6224002838135,
25.1508502960205,
-51.6127090454102,
-7.10364341735840,
15.6023626327515,
59.1105384826660,
0.983683586120606,
-15.1172485351563,
33.7599716186523,
-35.1715354919434,
46.0340080261231,
16.5778121948242,
-8.66639232635498,
31.4137821197510,
-48.9792709350586,
-12.7953872680664,
21.0451469421387,
-24.4467830657959,
-13.4377346038818,
30.2234210968018,
-10.2701501846313,
24.0262336730957,
50.8203735351563,
-14.6506099700928,
26.7830810546875,
3.70615768432617,
-14.1037120819092,
32.3080139160156,
46.7581558227539,
7.48720073699951,
38.6268768310547,
36.7356300354004,
-27.4799671173096,
44.0762863159180,
-8.72252845764160,
18.8089828491211,
26.3994560241699,
14.3198299407959,
24.6658134460449,
-57.2233428955078,
13.2194375991821,
-19.0330734252930,
26.5025138854980,
-9.17392539978027,
-62.9906082153320,
58.6933670043945,
-9.17961120605469,
-42.9167404174805,
-36.2308731079102,
1.68600749969482,
-24.8795242309570,
-55.4952888488770,
-6.36824226379395,
14.4466638565063,
38.0781860351563,
-36.3420219421387,
5.34763908386231,
-13.2061080932617,
-9.56915569305420,
70.5565948486328,
-0.421130180358887,
12.3071594238281,
39.3329467773438,
38.4197959899902,
-12.7271471023560,
22.0183563232422,
29.9673652648926,
-37.9457893371582,
24.5029525756836,
1.01455879211426,
2.72262191772461,
15.1703567504883,
1.23862648010254,
-10.7004528045654,
-49.2151718139648,
-35.2033233642578,
-43.7144355773926,
25.5538406372070,
42.8042716979981,
-26.9586296081543,
-21.5355758666992,
-14.4108219146729,
-45.5426940917969,
-16.7255020141602,
17.1735248565674,
-37.2415695190430,
-42.2974624633789,
24.8548126220703,
44.3339271545410,
-18.1081848144531,
34.4567184448242,
0.164848327636719,
-45.5737152099609,
30.2368278503418,
26.4719886779785,
37.6404914855957,
-15.3659839630127,
-31.6535034179688,
-7.29747962951660,
30.5147514343262,
37.3973922729492,
-3.53191232681274,
-18.8254261016846,
-46.3852920532227,
-42.8567390441895,
-44.4928817749023,
-7.98199081420898,
35.3731842041016,
0.274625778198242,
-31.0947837829590,
-2.59812355041504,
21.7522563934326,
25.5522384643555,
12.5081348419189,
-1.08811330795288,
2.77249622344971,
37.5451087951660,
25.5616149902344,
11.5600938796997,
58.4596710205078,
-19.1494750976563,
-7.62979125976563,
50.8547363281250,
16.2161560058594,
14.8620853424072,
-13.8915205001831,
36.8840217590332,
25.3863334655762,
-3.40341377258301,
56.4957275390625,
49.9637374877930,
-20.7447662353516,
-36.8607406616211,
36.6673660278320,
-20.9887161254883,
-13.6414060592651,
34.9880065917969,
3.82325172424316,
-19.2299461364746,
-36.5286026000977,
51.2526245117188,
-11.7504072189331,
-15.6658496856689,
69.9248275756836,
-24.4425277709961,
-50.5020675659180,
18.2431831359863,
60.4270401000977,
21.3500785827637,
31.6650581359863,
12.4033775329590,
-43.8915710449219,
45.3304061889648,
20.7986888885498,
-24.9619483947754,
60.4184265136719,
-7.88487243652344,
-7.14164495468140,
39.6752586364746,
-4.83380126953125,
51.2341270446777,
-23.9411964416504,
-50.1441993713379,
48.1479339599609,
-27.2450733184814,
-13.8886823654175,
3.04708099365234,
-43.9675254821777,
58.6133384704590,
0.343638420104980,
-23.5658569335938,
13.9587240219116,
-44.9987716674805,
22.5873527526855,
-8.01752281188965,
17.9360218048096,
8.50144958496094,
-73.8174972534180,
27.3061180114746,
27.3422546386719,
43.5398483276367,
4.56367206573486,
-15.3063907623291,
-2.04090881347656,
-15.0675592422485,
60.1676826477051,
-15.9793157577515,
-37.0404968261719,
-10.1013545989990,
44.4717559814453,
-2.71599578857422,
19.4241294860840,
24.2035007476807,
-47.0970344543457,
50.0265197753906,
-48.1356353759766,
22.7938919067383,
18.8795719146729,
-61.7786979675293,
35.6308670043945,
7.78584575653076,
-34.3945617675781,
-12.5875520706177,
38.7324485778809,
-0.675968170166016,
-31.1247749328613,
-36.5592575073242,
15.3778371810913,
-13.6942443847656,
-35.9696960449219,
26.0500049591064,
-23.0176429748535,
18.9923133850098,
-24.7085914611816,
-30.9720764160156,
65.6989822387695,
0.961318969726563,
11.8182373046875,
40.6806907653809,
-21.8489532470703,
-36.3353309631348,
36.9951362609863,
24.2960205078125,
-12.1568622589111,
7.39813995361328,
8.57263946533203,
-4.95482778549194,
1.05753135681152,
40.3817024230957,
-8.90615272521973,
28.0889930725098,
7.67555713653564,
-60.0778007507324,
14.8685865402222,
43.6219406127930,
15.7358064651489,
-68.1606674194336,
8.34476661682129,
54.7945976257324,
-51.9468460083008,
2.43195343017578,
-16.2461700439453,
-61.7318801879883,
0.352561950683594,
-22.9408092498779,
-12.5101404190063,
53.6768798828125,
7.80387496948242,
15.8801822662354,
26.6984214782715,
-17.2682285308838,
34.5646896362305,
10.5153770446777,
30.1766433715820,
1.01848793029785,
-57.7777175903320,
4.02415084838867,
-37.5088272094727,
-2.83111143112183,
-15.1777591705322,
-45.0400466918945,
-34.8579483032227,
-58.5942726135254,
31.2783527374268,
11.3942995071411,
28.9729843139648,
-6.06468057632446,
-54.8324813842773,
49.8494262695313,
-20.8660087585449,
-32.4770507812500,
21.2454662322998,
-12.9740190505981,
-22.3398380279541,
-7.05019092559814,
33.1430969238281,
13.5625200271606,
-42.1340675354004,
-14.0841417312622,
-9.83323383331299,
-60.2017860412598,
-6.55519485473633,
-7.66947746276856,
-48.2357292175293,
4.45952987670898,
7.73934650421143,
-35.3931846618652,
-37.8660278320313,
34.1525840759277,
34.3004760742188,
-11.5039119720459,
-10.5996189117432,
-41.7301101684570,
-4.70984649658203,
42.5228958129883,
37.6723289489746,
6.43043708801270,
-25.6762485504150,
-29.3837547302246,
-14.2460279464722,
34.9354324340820,
32.6208381652832,
-0.504737854003906,
-13.8752832412720,
14.8085460662842,
-7.08901500701904,
-32.5441741943359,
52.0082473754883,
-6.66420030593872,
-71.8984527587891,
20.8032054901123,
37.5477828979492,
22.4145507812500,
5.66228389739990,
39.0144653320313,
34.0990982055664,
-57.6908874511719,
29.2497100830078,
70.6228866577148,
-0.530673980712891,
-5.57864093780518,
-31.5810317993164,
-36.3377838134766,
1.83148956298828,
19.4665431976318,
-6.97975063323975,
-51.2000694274902,
-43.1820678710938,
-27.6370773315430,
28.7441978454590,
24.6850166320801,
-54.4932479858398,
-12.4436950683594,
-9.23493003845215,
14.5637998580933,
7.92442989349365,
-13.8511819839478,
26.2786369323730,
-31.8219985961914,
37.4489517211914,
40.2477035522461,
9.68693161010742,
48.3072853088379,
-17.6858863830566,
16.5284118652344,
13.0336790084839,
1.63429069519043,
2.15350055694580,
-37.0905380249023,
55.9693679809570,
35.2502136230469,
-57.0393104553223,
38.2271499633789,
39.4276771545410,
-32.8852043151856,
29.3984813690186,
56.3360748291016,
26.2204780578613,
-9.53415679931641,
-6.19009113311768,
-0.983605861663818,
-19.7871246337891,
34.7864151000977,
40.4578399658203,
-18.0154953002930,
-25.3430328369141,
-28.9316482543945,
-12.9153966903687,
-8.61533927917481,
8.70738410949707,
25.8019008636475,
4.06507205963135,
-16.9152812957764,
-11.6865863800049,
20.0657691955566,
-25.3170852661133,
24.2045478820801,
35.9492874145508,
0.552556037902832,
60.4511184692383,
-6.90703582763672,
19.8802375793457,
25.2586021423340,
18.4809303283691,
21.8383712768555,
-43.8487396240234,
53.3614730834961,
15.0142850875855,
18.9880867004395,
3.15947818756104,
-29.3232955932617,
18.4776287078857,
-5.36711454391480,
-8.47276020050049,
-27.4814338684082,
14.2536249160767,
-48.4421386718750,
25.7082195281982,
13.2382392883301,
-4.94609737396240,
34.8442649841309,
-25.3596611022949,
24.4704551696777,
-41.5330200195313,
15.2480192184448,
42.8470306396484,
37.1976661682129,
-26.5725021362305,
-28.5023059844971,
31.4995384216309,
-36.3631057739258,
59.6300430297852,
-12.1339807510376,
-41.9852600097656,
32.9950981140137,
-34.9303092956543,
-30.4311027526855,
-11.9460639953613,
-10.2171115875244,
-57.2740173339844,
-8.16584300994873,
68.3169860839844,
10.7463340759277,
26.2165546417236,
3.35473728179932,
5.75441741943359,
36.3600463867188,
-16.0493583679199,
-34.9759368896484,
7.51416683197022,
60.6847534179688,
-32.2357940673828,
-4.75513648986816,
68.1842651367188,
-13.1278114318848,
-26.2726402282715,
40.9634017944336,
46.4249038696289,
-3.35895442962647,
18.4539070129395,
11.4164934158325,
37.2404479980469,
5.28204917907715,
5.41221714019775,
27.0966529846191,
12.6602268218994,
37.1820144653320,
-41.4457015991211,
12.8651456832886,
-3.72294139862061,
14.7204504013062,
67.7978515625000,
-48.1794471740723,
9.27816677093506,
53.8969612121582,
17.5041007995605,
29.5933246612549,
57.4479637145996,
36.1054763793945,
-51.8839797973633,
-14.6513719558716,
57.3982162475586,
11.1698293685913,
15.0144987106323,
1.16787242889404,
-66.4895248413086,
33.0804901123047,
17.0324821472168,
-34.9911727905273,
14.7276477813721,
-55.2735710144043,
-9.92436981201172,
25.0707397460938,
-9.73265457153320,
10.1624956130981,
40.8050918579102,
-18.4374122619629,
-16.0511970520020,
26.2316589355469,
-55.2805595397949,
21.5038166046143,
48.5982780456543,
13.7631206512451,
7.09618663787842,
-41.4777717590332,
-30.5462512969971,
-39.4886550903320,
-21.7180728912354,
21.6944236755371,
-5.33813381195068,
-4.21774196624756,
23.8705253601074,
-36.2428131103516,
-13.4607620239258,
44.6926383972168,
2.52301216125488,
9.90717220306397,
17.2824954986572,
37.7084350585938,
38.5859260559082,
10.6032476425171,
11.9327116012573,
-38.4167022705078,
37.0547943115234,
39.7659683227539,
-32.2334518432617,
16.8818969726563,
-18.3028202056885,
7.49399280548096,
12.5161952972412,
-10.8319215774536,
68.8200836181641,
13.8303632736206,
-28.9435920715332,
20.4992389678955,
-5.16117382049561,
-20.5355319976807,
4.28515338897705,
-10.2252397537231,
-13.4329147338867,
53.8317871093750,
-7.05709648132324,
-50.5579414367676,
64.9351806640625,
6.77117156982422,
-31.4688034057617,
51.0752029418945,
0.207150459289551,
6.35376453399658,
7.88368701934814,
-44.8830184936523,
26.2076377868652,
45.2292976379395,
9.78832817077637,
16.4437904357910,
-23.5480175018311,
-25.0256443023682,
27.1968898773193,
-21.0584487915039,
-39.6501770019531,
20.0504913330078,
-2.04431915283203,
-25.2543220520020,
17.0986366271973,
56.1972999572754,
21.8948097229004,
-15.9640445709229,
35.6490974426270,
56.8961868286133,
-19.9813022613525,
-23.5688896179199,
45.6707992553711,
-17.7091636657715,
-11.3330698013306,
32.6254692077637,
-9.27552318572998,
-39.8051910400391,
-26.7683448791504,
38.9471664428711,
-34.0850334167481,
-47.2135696411133,
-12.6518011093140,
-42.0378570556641,
-2.51907634735107,
-7.68499517440796,
-18.6995124816895,
7.41659259796143,
-26.4777755737305,
-29.8932991027832,
3.61269474029541,
-25.1488742828369,
-21.8198165893555,
9.78521347045898,
23.3353691101074,
-12.4340982437134,
15.3462715148926,
26.1692276000977,
-47.3954315185547,
-46.3154067993164,
2.91148853302002,
29.9325637817383,
-12.8883466720581,
20.3633460998535,
47.4563484191895,
7.35697460174561,
13.1349143981934,
34.7943649291992,
53.0433120727539,
0.322620391845703,
-51.8706016540527,
-1.43606090545654,
14.1664400100708,
10.3907670974731,
11.5894632339478,
-37.8420982360840,
17.6406974792480,
9.09536933898926,
-37.5579719543457,
39.8455657958984,
41.0232925415039,
9.57559776306152,
-30.2502307891846,
-0.911377906799316,
51.1301422119141,
-41.9238967895508,
-55.1079025268555,
11.6711015701294,
16.5579414367676,
18.4167995452881,
6.10878181457520,
41.3134384155273,
37.5872459411621,
-31.3575992584229,
-11.6987609863281,
-17.8451881408691,
-6.49991273880005,
-9.07980823516846,
-57.6958427429199,
8.43241596221924,
18.9648780822754,
-4.60720872879028,
24.3823471069336,
-16.5259017944336,
55.0003814697266,
32.8328247070313,
-64.1810531616211,
56.7091064453125,
25.1206455230713,
14.5590620040894,
44.7710609436035,
-46.4370384216309,
-9.30367279052734,
-24.7330093383789,
-43.0589485168457,
2.81798171997070,
-46.2541618347168,
-52.7495384216309,
8.82168579101563,
-35.6443939208984,
-64.1369781494141,
10.4932680130005,
14.9357776641846,
12.8615427017212,
-3.95335006713867,
-23.6198768615723,
-1.97395086288452,
16.7961254119873,
18.3600883483887,
-41.5782203674316,
26.5100021362305,
29.2749481201172,
-59.2466278076172,
-27.7191047668457,
-22.5177516937256,
-11.7515163421631,
-43.2840728759766,
-0.00784206390380859,
20.6346588134766,
-24.5103416442871,
1.87738800048828,
-1.56352329254150,
38.8716354370117,
-31.8615016937256,
12.3790302276611,
36.9699554443359,
-23.4339866638184,
64.8818283081055,
-6.02566719055176,
-11.3714160919189,
-31.4772434234619,
-57.8794403076172,
39.2410888671875,
39.9564132690430,
-16.9676532745361,
11.9379978179932,
43.5558738708496,
-18.5553932189941,
52.2154388427734,
37.1670036315918,
-21.7039947509766,
43.1599693298340,
0.354120254516602,
-32.9749565124512,
-0.941255092620850,
27.0709419250488,
46.0402679443359,
16.8890686035156,
-7.45341014862061,
9.35290145874023,
3.37125873565674,
-5.60563564300537,
-26.4626502990723,
-38.9597396850586,
-18.0466728210449,
-54.3430099487305,
-13.2541713714600,
-7.23255491256714,
-22.9612579345703,
34.2743263244629,
-0.594098091125488,
44.1909484863281,
32.3213653564453,
-27.1047897338867,
-21.5531692504883,
-26.5030975341797,
-7.07186460494995,
-41.4485397338867,
-29.4778251647949,
24.6309318542480,
36.1782608032227,
-14.4360656738281,
-32.8074226379395,
4.46827793121338,
16.2313346862793,
27.7068691253662,
-28.8472900390625,
-4.57368946075439,
29.5147819519043,
2.07722377777100,
11.8021812438965,
-2.63564300537109,
-0.236956596374512,
-1.81041431427002,
43.4867248535156,
-17.5271434783936,
-31.6881389617920,
66.9013977050781,
-28.3182926177979,
-10.6595411300659,
13.6600484848022,
-68.2465515136719,
-0.309565544128418,
-11.6696653366089,
-42.1086349487305,
34.9179534912109,
27.0775299072266,
-3.21547412872314,
11.7933082580566,
19.7873210906982,
-16.3654747009277,
-52.6863594055176,
-24.3422966003418,
9.28808593750000,
21.7759265899658,
-29.5757503509522,
0.249155044555664,
46.2358703613281,
-10.8143262863159,
28.4380722045898,
25.2523803710938,
28.6406135559082,
10.9124364852905,
25.8823661804199,
30.3750648498535,
-29.8440437316895,
51.0786437988281,
20.5083751678467,
-31.7157382965088,
-2.06492471694946,
38.1859970092773,
12.7936992645264,
-21.1262283325195,
-34.0290222167969,
-23.3178844451904,
-41.9092636108398,
-23.9901466369629,
44.5480346679688,
-38.8602523803711,
17.3070411682129,
-36.5418205261231,
-8.92037105560303,
63.6932106018066,
-76.4543304443359,
23.6335945129395,
27.2224674224854,
2.90034198760986,
33.6113281250000,
-27.4259681701660,
45.5017280578613,
34.6416511535645,
-10.8523120880127,
48.9821815490723,
56.0025024414063,
16.9033279418945,
14.7259082794189,
27.5708007812500,
2.50553798675537,
31.2699966430664,
46.2023849487305,
39.2321815490723,
6.65431118011475,
-27.2822380065918,
-6.12881851196289,
-42.3791084289551,
13.0707931518555,
72.0370788574219,
2.21053314208984,
-1.38177299499512,
12.0942802429199,
-18.3541908264160,
34.5587615966797,
51.5144271850586,
19.2620658874512,
41.7227401733398,
-15.5009508132935,
17.9787921905518,
22.1128978729248,
-1.15262842178345,
39.8558959960938,
-42.4653854370117,
-21.1690864562988,
8.41056823730469,
37.7694015502930,
38.4052276611328,
-50.7322616577148,
-11.0425338745117,
51.0279121398926,
6.10852050781250,
-40.8294792175293,
-23.5439529418945,
-16.2629184722900,
-29.3246688842773,
-2.65511989593506,
-17.4677238464355,
-30.8054351806641,
1.16891288757324,
-25.8865356445313,
18.5046749114990,
-33.2903404235840,
-16.2770996093750,
45.6498146057129,
-34.2747535705566,
-2.05323123931885,
-3.35795736312866,
14.2395381927490,
25.9007263183594,
20.9381141662598,
28.8785400390625,
24.6374378204346,
45.3626403808594,
36.4035034179688,
31.4277515411377,
42.3536300659180,
31.9184265136719,
-33.0712661743164,
1.86664390563965,
2.42016696929932,
-24.0605506896973,
-14.1775398254395,
-58.4299850463867,
13.5282192230225,
-17.3606758117676,
-48.1682739257813,
24.4776191711426,
22.6511058807373,
2.86329460144043,
-5.02070283889771,
48.7755966186523,
16.2522888183594,
-1.22093439102173,
-19.4292316436768,
-16.9232864379883,
38.3511657714844,
18.5298309326172,
10.8790569305420,
5.36988830566406,
-2.80389308929443,
21.2117424011230,
36.3650817871094,
-43.6669006347656,
7.74608516693115,
47.2990379333496,
-26.6261863708496,
1.30793094635010,
11.6975135803223,
-15.9805679321289,
-16.6263065338135,
53.3251419067383,
36.0455894470215,
-22.6480827331543,
36.0718917846680,
10.6274900436401,
-37.6140594482422,
26.0106048583984,
39.5084075927734,
22.8120326995850,
21.6313934326172,
40.1588287353516,
40.2309455871582,
-34.7818069458008,
11.4438438415527,
38.7056655883789,
-2.88537740707397,
19.3197631835938,
0.499788284301758,
9.06908321380615,
22.5829734802246,
-15.1046361923218,
-22.4155139923096,
-37.2614669799805,
-26.7190246582031,
10.9156360626221,
-47.7989196777344,
-25.3972129821777,
28.9561500549316,
24.5384864807129,
25.5804328918457,
-15.4210662841797,
-22.8023986816406,
26.8956680297852,
43.4175148010254,
28.4097023010254,
39.2549362182617,
-9.98569679260254,
23.4025573730469,
56.6161499023438,
-26.8320922851563,
0.480150222778320,
56.0972709655762,
-10.6285486221313,
9.73720073699951,
51.6232604980469,
-31.8985214233398,
-42.8404006958008,
10.3378009796143,
47.0719528198242,
2.35323810577393,
0.666980743408203,
-20.0593357086182,
10.9448604583740,
31.3984947204590,
-8.14929389953613,
3.18445968627930,
-35.2481155395508,
35.1827545166016,
-10.7932977676392,
0.516477584838867,
4.57238674163818,
-16.8471946716309,
53.4401664733887,
-33.3121490478516,
-0.880241394042969,
26.6801528930664,
29.2797088623047,
-15.0149192810059,
-8.14612102508545,
55.6282424926758,
-12.6749143600464,
-31.0244064331055,
-19.6227855682373,
60.2630996704102,
-1.22481441497803,
-55.4029464721680,
28.2105827331543,
-50.7984809875488,
-54.9804611206055,
-27.0725631713867,
-5.14926719665527,
15.5465049743652,
2.34801197052002,
39.7750396728516,
-65.7635421752930,
11.1781215667725,
42.5543098449707,
-62.4409561157227,
-0.0718107223510742,
-31.7868690490723,
27.3397483825684,
-25.5902233123779,
-81.6838989257813,
39.3286743164063,
36.1348037719727,
-12.0107011795044,
-10.3222084045410,
39.9163360595703,
-7.18134784698486,
-34.8235969543457,
50.9517707824707,
54.6347732543945,
-5.69074344635010,
-0.0636529922485352,
-21.4414634704590,
-8.62534999847412,
62.3487052917481,
-0.248663902282715,
-56.7728157043457,
37.6095275878906,
36.4064750671387,
-32.5124359130859,
51.5753746032715,
-1.32183551788330,
-58.4753799438477,
14.6727085113525,
-5.83342266082764,
-8.29753017425537,
-20.8320083618164,
-26.2887496948242,
-21.2145957946777,
-53.8489570617676,
-27.0745162963867,
25.6512451171875,
32.7762107849121,
11.0415630340576,
43.2455291748047,
10.9078330993652,
-27.6657257080078,
45.4202384948731,
-10.2700099945068,
-25.3457641601563,
25.4999866485596,
28.0753479003906,
25.4792213439941,
-45.2428741455078,
3.57058620452881,
28.6992435455322,
15.3311214447021,
19.1873798370361,
40.8587951660156,
29.6693878173828,
4.14662361145020,
46.2627639770508,
5.91911888122559,
7.83404731750488,
-24.5082454681397,
-10.1035432815552,
3.99192810058594,
2.99063014984131,
-8.07098770141602,
13.4123067855835,
32.7036056518555,
-40.4490661621094,
-22.0449829101563,
-33.4350357055664,
13.2269773483276,
-33.1864318847656,
5.49059772491455,
48.3018493652344,
-24.1206340789795,
39.2248764038086,
43.9486732482910,
-14.9218540191650,
-31.9727249145508,
36.4812431335449,
-32.8815841674805,
-28.7641010284424,
55.4124984741211,
-9.53606224060059,
-8.10219383239746,
7.77841567993164,
18.0537147521973,
45.8475265502930,
28.7834663391113,
32.1174545288086,
7.28819084167481,
-7.29757976531982,
58.5115318298340,
3.48663425445557,
-29.7731590270996,
-0.382974624633789,
-36.0012664794922,
-6.06684017181397,
25.2088222503662,
37.9409408569336,
-4.56588172912598,
-16.2383995056152,
18.7839164733887,
-38.0361862182617,
9.64838123321533,
55.6824645996094,
-21.7249183654785,
-35.1577262878418,
4.72038841247559,
19.0296840667725,
25.7417259216309,
34.1675262451172,
23.2064514160156,
-36.0188903808594,
-19.4032592773438,
5.03656291961670,
-38.8219451904297,
31.6662845611572,
-22.4817619323730,
-39.0851173400879,
30.5895309448242,
-21.3383331298828,
-8.52800750732422,
-7.35954284667969,
-19.9410057067871,
-15.8391523361206,
41.6668205261231,
6.73886680603027,
13.4643774032593,
49.5210342407227,
-45.2698745727539,
-2.27182006835938,
46.0457229614258,
10.1328258514404,
-35.0362968444824,
5.22019958496094,
11.0908155441284,
-40.9655532836914,
-19.3847713470459,
-13.3384408950806,
-8.15238857269287,
-28.2910938262939,
-40.0296592712402,
-0.439016342163086,
15.3437547683716,
38.1031799316406,
26.3362026214600,
15.5146579742432,
50.7769393920898,
-21.8386230468750,
-45.1124992370606,
-22.8485717773438,
-27.2224884033203,
-13.2482872009277,
9.15311241149902,
7.68868064880371,
-53.8017234802246,
-30.4748573303223,
-31.1961135864258,
12.2109966278076,
55.8926391601563,
-49.4245758056641,
-29.3605022430420,
54.2621231079102,
33.4303894042969,
26.2604274749756,
16.5156097412109,
27.0323715209961,
49.5678482055664,
-11.2315654754639,
38.1814422607422,
21.7407245635986,
-66.9232788085938,
22.8540840148926,
39.1693153381348,
25.5446701049805,
21.9450607299805,
-10.9207258224487,
19.3160419464111,
-46.2862472534180,
-28.3894252777100,
10.7415466308594,
-51.7849349975586,
22.1611366271973,
-9.31571483612061,
-38.2113113403320,
-39.1773529052734,
-21.7402935028076,
42.0898590087891,
-43.2524719238281,
-14.0305404663086,
21.8824310302734,
14.9670906066895,
-29.7380561828613,
-52.0574798583984,
-21.1910018920898,
-14.3846950531006,
51.3724746704102,
12.9095535278320,
-44.2752342224121,
-17.4390468597412,
47.8037185668945,
-6.80410766601563,
-15.7632198333740,
51.0556564331055,
-34.8050994873047,
-33.5256042480469,
-13.6772985458374,
3.54104804992676,
39.5639877319336,
-45.7119293212891,
8.20059204101563,
52.1826324462891,
-22.1894149780273,
22.6267356872559,
50.5455017089844,
5.33722114562988,
-62.8483428955078,
18.7283401489258,
40.7441558837891,
-49.0478897094727,
4.01936340332031,
-14.5266761779785,
-53.7186660766602,
5.08670234680176,
41.8669967651367,
-32.5679321289063,
-52.6376724243164,
-25.3077812194824,
0.763422012329102,
-4.30904340744019,
-10.7537870407105,
22.3485183715820,
-26.5477371215820,
-10.1969184875488,
-9.79669761657715,
-5.00348281860352,
36.4789657592773,
-15.7644844055176,
-73.4656066894531,
19.3410377502441,
23.6995506286621,
-40.1337623596191,
33.8946304321289,
19.6361713409424,
27.5401191711426,
-42.0807228088379,
8.08186244964600,
80.7796478271484,
-3.38924360275269,
36.1733398437500,
-16.1644325256348,
0.803613662719727,
0.396718025207520,
-18.1332511901855,
53.6792564392090,
26.1817417144775,
16.6228027343750,
-20.6920394897461,
-24.2319374084473,
-5.45829868316650,
4.75737571716309,
12.9669513702393,
-24.0756130218506,
10.9545879364014,
11.1697711944580,
5.23867034912109,
16.7104835510254,
20.4759902954102,
23.1164054870605,
3.70996189117432,
41.1611785888672,
6.38632202148438,
-33.1040840148926,
-18.1600685119629,
-27.1647186279297,
1.48858451843262,
25.3111572265625,
26.7527122497559,
-16.8731384277344,
4.29966545104981,
46.1579818725586,
-59.0901222229004,
8.01870822906494,
50.9156837463379,
-36.7229690551758,
-15.2096338272095,
27.3777961730957,
43.9002838134766,
15.1738624572754,
40.9618797302246,
15.4400730133057,
18.8395862579346,
13.8478736877441,
-28.4075584411621,
-1.30118942260742,
38.4906654357910,
15.4179115295410,
-13.3621978759766,
38.8212432861328,
-20.2200012207031,
-26.8072528839111,
12.1897983551025,
17.8554763793945,
-8.95465373992920,
-30.8722801208496,
-9.88676643371582,
-37.9451293945313,
18.2099075317383,
33.8754310607910,
-40.3116645812988,
-51.5018959045410,
22.5376625061035,
0.900742530822754,
-61.8302078247070,
-10.0314273834229,
-10.4644088745117,
-16.1843891143799,
-26.4661178588867,
-0.854402542114258,
43.7472381591797,
13.1572542190552,
-2.63486337661743,
-31.3492088317871,
29.8146209716797,
62.0232772827148,
-36.0012054443359,
-31.1044445037842,
4.33037090301514,
-44.4323272705078,
-51.1526603698731,
4.01962280273438,
-9.31385326385498,
4.14359855651856,
30.5759220123291,
-19.5719203948975,
-50.4771881103516,
-7.88850498199463,
32.5891418457031,
-19.9475307464600,
55.0453338623047,
25.4965667724609,
-58.8878936767578,
3.85136890411377,
17.0716705322266,
46.7133140563965,
-0.0185117721557617,
23.2485466003418,
-14.6468133926392,
-8.72491836547852,
18.5992851257324,
-29.2934570312500,
20.6006603240967,
-14.4225530624390,
-14.4853096008301,
-30.2589626312256,
17.4583034515381,
6.47240734100342,
-4.76215600967407,
41.3522644042969,
-9.56470394134522,
-19.7635421752930,
6.50266170501709,
48.0576248168945,
-21.9083404541016,
-26.8522300720215,
-18.8730850219727,
-50.5988159179688,
-20.8173255920410,
8.70933532714844,
13.0621347427368,
-36.0651931762695,
32.4653549194336,
0.846976280212402,
-59.4038352966309,
30.4836997985840,
15.8934803009033,
21.7528686523438,
-6.98691797256470,
-38.2946434020996,
22.8495273590088,
15.0128726959229,
-2.32112789154053,
-8.88741874694824,
-18.6704597473145,
-19.2403373718262,
-21.8190422058105,
-15.8518943786621,
37.4299468994141,
-12.8459587097168,
-74.1006088256836,
8.79864215850830,
38.5417747497559,
5.58788871765137,
-49.4583625793457,
14.6781558990479,
-10.1522283554077,
-25.6557655334473,
57.7701110839844,
-9.06204605102539,
18.9798355102539,
-26.8361492156982,
17.3819828033447,
37.3240661621094,
-13.8146476745605,
16.5651741027832,
-61.8900985717773,
35.3667526245117,
39.6072158813477,
1.23317623138428,
47.5840682983398,
42.7085113525391,
30.3960762023926,
-44.1329345703125,
11.7338314056396,
74.8365249633789,
-9.88038635253906,
-54.4002647399902,
30.0072536468506,
-12.1082248687744,
-28.9369544982910,
58.5054969787598,
-4.33112716674805,
35.4900817871094,
-0.587321281433106,
-18.5140686035156,
47.0737915039063,
7.74600124359131,
4.37928009033203,
-56.6450042724609,
-30.6002464294434,
-34.0146865844727,
5.91359519958496,
50.9692840576172,
-15.4690036773682,
42.4692993164063,
-7.66698503494263,
-6.81778717041016,
51.9360809326172,
16.5685596466064,
33.8813362121582,
-27.1087570190430,
55.5053787231445,
39.3911209106445,
-54.1813430786133,
41.8668937683106,
-4.45425891876221,
35.0938339233398,
-13.5612239837646,
-6.79545211791992,
34.1921463012695,
-30.4796981811523,
48.9468269348145,
-22.0695438385010,
17.9747352600098,
7.78060531616211,
-13.6440372467041,
58.6626968383789,
-23.6154365539551,
-39.3439636230469,
-23.1566619873047,
56.8732681274414,
16.4877681732178,
-35.6086654663086,
-27.6694431304932,
-35.3275337219238,
-9.46992778778076,
-38.7632827758789,
36.3185882568359,
-18.2992954254150,
-69.6600723266602,
-31.1680469512939,
-11.2864809036255,
30.2864551544189,
13.4909143447876,
-7.64843082427979,
-54.4427375793457,
46.1210937500000,
37.2191696166992,
16.6241149902344,
35.0123405456543,
-53.6856918334961,
29.2215671539307,
-4.08881664276123,
-47.3333053588867,
-11.6275072097778,
-46.3888092041016,
-40.1638946533203,
3.89910888671875,
42.3585281372070,
-22.5716094970703,
-63.5862731933594,
-6.40914249420166,
14.4765548706055,
4.33120155334473,
-29.2285556793213,
-1.59223556518555,
35.3814659118652,
-13.5554981231689,
-25.8379974365234,
3.15562152862549,
15.6030950546265,
-34.6250228881836,
-29.8240089416504,
-15.4273061752319,
24.6691436767578,
21.2310676574707,
-37.0656814575195,
-2.85182762145996,
9.44624710083008,
41.6537055969238,
-33.3009834289551,
-56.6458511352539,
-3.35047149658203,
-11.8885354995728,
-14.3792352676392,
5.04067325592041,
24.3057785034180,
-46.4066429138184,
-31.2913017272949,
-11.9056682586670,
-20.9445381164551,
-28.7343635559082,
-0.406874656677246,
-6.19651174545288,
-41.8321037292481,
11.6914348602295,
-31.5293540954590,
2.85592174530029,
-8.77295684814453,
-42.1274185180664,
27.1093597412109,
-36.9167785644531,
0.459632873535156,
22.7794837951660,
-21.9275760650635,
7.37865161895752,
26.1507358551025,
12.3674526214600,
-10.4534683227539,
26.3112030029297,
-26.8649940490723,
-15.8408927917480,
51.9290771484375,
17.5199623107910,
15.4789361953735,
16.7931499481201,
-0.0378952026367188,
12.6402711868286,
16.5309066772461,
16.6088294982910,
3.64285373687744,
13.1769723892212,
17.5041465759277,
-43.1045455932617,
-5.95051860809326,
-6.11347675323486,
-1.27002620697021,
-6.02175903320313,
-17.6797447204590,
63.9980773925781,
3.49474906921387,
-12.3618631362915,
7.13413619995117,
-42.5031585693359,
-30.3859348297119,
-0.713194847106934,
-9.65219020843506,
-30.7563247680664,
11.5469350814819,
36.4260406494141,
-13.3002748489380,
-35.7313919067383,
14.4836606979370,
-3.15761089324951,
-4.34343910217285,
-27.1672916412354,
-65.1261901855469,
43.3868331909180,
-20.5700511932373,
-21.6701850891113,
19.4346733093262,
-11.0272493362427,
38.9410171508789,
-60.5610160827637,
1.66993141174316,
27.2289981842041,
-51.1924171447754,
1.13556766510010,
-9.85755634307861,
8.91477489471436,
-21.3339271545410,
-5.29113292694092,
7.61320781707764,
-35.4947166442871,
26.7993392944336,
14.6502408981323,
-14.4980983734131,
15.2369794845581,
-13.3581285476685,
-51.6512222290039,
8.26034259796143,
16.4357223510742,
13.3327016830444,
13.1196584701538,
-9.58450317382813,
27.7733173370361,
26.3103561401367,
35.9296531677246,
-17.0475273132324,
-46.6679687500000,
12.4261131286621,
41.8103408813477,
-21.5601081848145,
-18.6787147521973,
30.2619686126709,
-22.7358417510986,
17.0873565673828,
-24.9501647949219,
-13.1139240264893,
60.0698547363281,
-55.1954841613770,
4.05856323242188,
81.4800872802734,
-3.70182704925537,
9.82660198211670,
7.58929538726807,
-1.27992773056030,
-2.06888103485107,
11.5453586578369,
10.3416776657105,
-35.1999588012695,
31.4635620117188,
9.84915637969971,
-1.39034795761108,
-22.9710884094238,
-16.7811985015869,
50.9690818786621,
-76.6979675292969,
1.79446125030518,
45.5197372436523,
-44.9070243835449,
42.1151847839356,
31.4409255981445,
12.2710638046265,
15.4476823806763,
17.8392906188965,
10.6680269241333,
-61.6376457214356,
3.92396163940430,
40.2717361450195,
-63.7728347778320,
-32.0871086120606,
44.6410140991211,
6.68932628631592,
-47.0487594604492,
2.52102756500244,
52.8450393676758,
18.3561401367188,
24.5513458251953,
4.03223800659180,
15.8311033248901,
-12.3421850204468,
-43.9900665283203,
54.7963333129883,
12.2905073165894,
-0.918706893920898,
2.53529834747314,
-6.48536205291748,
38.4680938720703,
29.5078773498535,
13.3080282211304,
-29.2877235412598,
41.5330505371094,
30.4188194274902,
-52.8506126403809,
8.74308204650879,
35.4963836669922,
-11.0753135681152,
-16.0338096618652,
-22.6466445922852,
-5.97179794311523,
29.0315799713135,
-28.8016357421875,
-12.7769136428833,
18.5589218139648,
-38.1060562133789,
-24.0779857635498,
41.1743927001953,
15.2825202941895,
12.6238727569580,
33.3699111938477,
-30.5911483764648,
-35.1334152221680,
-26.3964729309082,
5.38689613342285,
-25.0653877258301,
-49.4202041625977,
27.3084945678711,
-50.0879211425781,
-20.7570934295654,
27.1178970336914,
-36.0472793579102,
-64.9968414306641,
-14.4532909393311,
28.8595809936523,
-61.8237800598145,
16.6486301422119,
3.98077583312988,
-59.4886245727539,
0.996520996093750,
11.9767980575562,
45.3432464599609,
24.1603507995605,
4.11392116546631,
-5.74277639389038,
-6.66566705703735,
29.8292922973633,
14.7855615615845,
-18.9003868103027,
-26.2367134094238,
-51.5056343078613,
-4.33772468566895,
6.72626972198486,
-14.0376930236816,
0.740103721618652,
25.3843803405762,
33.0112419128418,
-55.0764732360840,
-22.5839099884033,
-17.7536354064941,
-63.9449768066406,
-28.8099288940430,
21.9431114196777,
35.0337524414063,
8.73263835906982,
50.8314781188965,
0.0208120346069336,
-42.1403236389160,
59.3162002563477,
11.6246480941772,
-30.4495277404785,
51.9310417175293,
-15.6178159713745,
-3.23823976516724,
29.2003021240234,
-23.7316131591797,
4.17606258392334,
-12.9490680694580,
-23.0032291412354,
3.48379516601563,
26.2072753906250,
8.68957042694092,
-38.4664535522461,
16.1072006225586,
76.6407470703125,
-48.9064407348633,
-9.26861572265625,
48.6127815246582,
-69.1127014160156,
17.2914810180664,
31.0248069763184,
-23.0506706237793,
-40.6576843261719,
6.50833511352539,
46.1520652770996,
-29.5705146789551,
28.0417385101318,
-1.00662517547607,
-42.6491012573242,
-0.544690132141113,
10.6225919723511,
49.3991546630859,
8.72807407379150,
-10.9577970504761,
25.2439231872559,
4.88362789154053,
-20.5447425842285,
6.73822307586670,
7.10500717163086,
25.4761962890625,
17.7942848205566,
-22.7423057556152,
58.1352005004883,
33.8819580078125,
22.1344413757324,
26.6963119506836,
-26.5845451354980,
16.2898826599121,
-2.81073379516602,
10.3773279190063,
-3.13911533355713,
-34.0697402954102,
18.8884086608887,
8.93252468109131,
-55.6886787414551,
-20.3696861267090,
47.1400527954102,
-13.8125114440918,
22.4292678833008,
24.8052215576172,
-31.4588050842285,
47.9201850891113,
25.9744205474854,
-24.1271705627441,
45.2451019287109,
47.6313858032227,
23.4768791198730,
2.75160026550293,
-45.1625862121582,
11.5192785263062,
-14.6884622573853,
7.98596477508545,
-4.40595722198486,
-22.8817329406738,
27.1428909301758,
-51.2005386352539,
38.0851936340332,
-28.9007434844971,
0.976807594299316,
75.8478698730469,
-63.3579521179199,
20.2903289794922,
46.4973640441895,
-5.04094791412354,
-44.5125389099121,
-11.5012016296387,
46.1517257690430,
21.2136993408203,
-47.2553710937500,
3.19038009643555,
66.6528701782227,
-50.6793594360352,
29.7376613616943,
13.8978958129883,
-43.2863922119141,
71.8272552490234,
34.2110137939453,
35.6784172058106,
-27.9953689575195,
-52.8274688720703,
48.1581192016602,
41.7745475769043,
-2.81796550750732,
-2.93131923675537,
16.9490013122559,
35.9988174438477,
20.2455310821533,
-28.8597888946533,
64.5998916625977,
-11.5276584625244,
-6.44353199005127,
85.8670806884766,
-37.5106430053711,
42.0952796936035,
-1.00656318664551,
-24.2068805694580,
1.17984104156494,
-14.2344017028809,
23.5127754211426,
-56.3043441772461,
30.7185859680176,
-27.0133686065674,
-25.7779121398926,
31.4988803863525,
-8.06641292572022,
56.5606307983398,
-21.7838478088379,
-18.3154220581055,
-35.9456481933594,
7.43547248840332,
-9.11378479003906,
-50.8844985961914,
41.0908317565918,
-27.1905822753906,
28.6128311157227,
1.99673938751221,
-15.2071838378906,
5.36625099182129,
-16.4381771087647,
37.0478363037109,
0.498617172241211,
21.1450481414795,
-29.0221748352051,
27.2433109283447,
40.6196327209473,
-58.2784423828125,
-20.5123310089111,
-17.8341407775879,
5.84580326080322,
11.4818935394287,
31.9875144958496,
7.25023460388184,
-28.7486381530762,
12.9437007904053,
9.75467395782471,
-26.6314907073975,
14.1638898849487,
18.7943916320801,
-60.1656990051270,
41.3808898925781,
10.3014726638794,
-46.6297988891602,
52.6462478637695,
9.19704151153565,
24.2584838867188,
27.1704292297363,
22.7888469696045,
40.7326469421387,
-9.08494663238525,
12.9511270523071,
36.9910583496094,
-6.27328681945801,
3.85306644439697,
9.72337913513184,
-32.2730407714844,
11.6748619079590,
-6.19482040405273,
-52.2593078613281,
-48.2461853027344,
20.0615520477295,
37.0387458801270,
-40.4102935791016,
-14.8021707534790,
-11.0948009490967,
6.31124877929688,
1.50563526153564,
-39.5030136108398,
-29.7730331420898,
-22.2705421447754,
-13.3573122024536,
-31.9519672393799,
5.72734165191650,
21.7204475402832,
-40.3904190063477,
-30.7857112884522,
24.4649810791016,
-25.0230674743652,
-56.3308067321777,
22.8304405212402,
30.9306297302246,
5.19972896575928,
1.68220901489258,
-8.04994773864746,
-43.8336906433106,
-0.371047019958496,
31.6752223968506,
-34.0102424621582,
5.85769748687744,
9.66152858734131,
6.35611438751221,
-12.5578165054321,
5.49696540832520,
73.6356124877930,
-20.3022518157959,
-25.6252174377441,
-24.3494606018066,
-33.2574386596680,
-15.2552413940430,
-20.3094139099121,
-18.2742958068848,
-42.6003570556641,
2.52972888946533,
-2.28381347656250,
-1.63020944595337,
-24.8269805908203,
39.9865875244141,
-1.69212627410889,
-48.0422554016113,
37.7954750061035,
-30.6494331359863,
5.58441638946533,
-3.54761695861816,
29.6092567443848,
11.2170934677124,
12.3890628814697,
8.63981151580811,
-19.3532409667969,
31.2139854431152,
-57.4551086425781,
-42.7163276672363,
-5.37245941162109,
35.4353332519531,
-49.0540847778320,
-6.38066387176514,
74.9852447509766,
-11.6510534286499,
-40.9309844970703,
16.5553550720215,
61.9475669860840,
19.4927215576172,
40.4258155822754,
-27.2295112609863,
-23.4861621856689,
-14.7949485778809,
-47.0494461059570,
-29.4689903259277,
-21.7218265533447,
-58.8233184814453,
-23.6898975372314,
23.4834117889404,
1.47416400909424,
44.6780853271484,
-6.62759780883789,
-47.1866073608398,
-36.2615547180176,
30.6720924377441,
17.6475372314453,
-13.9884080886841,
-22.9238395690918,
-46.8521842956543,
-35.5558891296387,
-20.1222553253174,
12.5653047561646,
-39.1433944702148,
15.5266447067261,
28.1789436340332,
4.31846046447754,
-7.13327980041504,
-5.71068954467773,
9.73062038421631,
-50.7509040832520,
16.5831375122070,
18.5519046783447,
14.1437120437622,
-22.1604671478272,
-46.9837417602539,
-18.5419845581055,
-67.8891067504883,
38.7398490905762,
-2.08826780319214,
-18.9634895324707,
58.5011215209961,
14.9496879577637,
17.1988983154297,
-19.8241539001465,
-5.86375856399536,
-30.3001327514648,
-17.2519416809082,
-25.3409938812256,
-40.4795875549316,
27.3799896240234,
-36.4208412170410,
-31.4964466094971,
-14.3273744583130,
13.8953819274902,
34.2987785339356,
-62.6847801208496,
2.87193393707275,
50.3324699401856,
-52.3416366577148,
19.0281524658203,
60.1040344238281,
-30.7289657592773,
-22.9450721740723,
-26.0411567687988,
10.7347335815430,
11.6398906707764,
-53.9433250427246,
-21.5265121459961,
-32.1215286254883,
-57.3029022216797,
-42.6898269653320,
-15.4218883514404,
-0.728341102600098,
-42.6470031738281,
-59.2910690307617,
2.01591014862061,
1.78288269042969,
-62.8470039367676,
-8.20286655426025,
32.2009849548340,
-12.8765878677368,
-28.8204154968262,
-15.7630958557129,
-23.9315986633301,
14.5308494567871,
30.9086380004883,
-6.98649787902832,
9.79574203491211,
-16.1657791137695,
-26.0676422119141,
27.7816467285156,
58.6733322143555,
-34.4105987548828,
-18.8170948028564,
35.0781974792481,
-66.8234710693359,
0.0298080444335938,
31.1248893737793,
1.51918029785156,
33.4815521240234,
-26.0445289611816,
29.1905708312988,
30.3537769317627,
-53.4846687316895,
25.6989135742188,
0.308885574340820,
-45.2773513793945,
32.9687538146973,
38.0405235290527,
3.24303817749023,
48.2187156677246,
51.1247711181641,
-40.9419136047363,
17.3023662567139,
31.9041671752930,
-15.1978979110718,
2.48088932037354,
-1.10051870346069,
-13.9771442413330,
-46.1057090759277,
31.8682632446289,
-12.6189432144165,
-65.5909271240234,
47.5959281921387,
11.2909307479858,
-21.1990776062012,
33.5836830139160,
-22.3347778320313,
-13.3451251983643,
39.4919204711914,
-36.8485870361328,
12.7237129211426,
51.2100753784180,
18.4190750122070,
37.0225982666016,
-28.7786827087402,
28.9621448516846,
27.1956787109375,
-16.3290004730225,
27.7853050231934,
-53.4422378540039,
-11.8230562210083,
31.0881805419922,
20.7066497802734,
36.5505676269531,
-5.40333461761475,
26.7826213836670,
39.7743911743164,
15.0344200134277,
1.08512115478516,
14.3899841308594,
52.8055648803711,
-43.9051818847656,
-25.3964576721191,
70.6180877685547,
-10.9709272384644,
-18.0965805053711,
24.8387451171875,
0.461510658264160,
-44.9883651733398,
7.85619735717773,
10.5253934860230,
-31.8528327941895,
-6.66588592529297,
-40.2801284790039,
34.0265312194824,
-10.4879207611084,
-39.4738883972168,
46.3923416137695,
-48.4874954223633,
23.8971347808838,
17.4081497192383,
-58.7304496765137,
44.0199012756348,
21.6752986907959,
-9.75959014892578,
25.5688629150391,
44.6487998962402,
3.79644203186035,
-24.8880996704102,
-36.6224098205566,
19.0761299133301,
55.5912399291992,
-46.9934349060059,
-29.8509864807129,
32.9706077575684,
4.05496215820313,
-58.7760581970215,
-8.44545173645020,
62.0294647216797,
-37.2836799621582,
-22.2827186584473,
12.4863061904907,
-40.5650711059570,
5.59274005889893,
-8.95928192138672,
6.74482250213623,
7.69710731506348,
-50.4150161743164,
-14.2486200332642,
27.6345882415772,
46.3629417419434,
-16.5632572174072,
-4.07975769042969,
42.1256599426270,
24.9930820465088,
4.76487350463867,
9.10338211059570,
55.5495300292969,
-8.17615509033203,
-50.5943336486816,
-27.0105075836182,
-7.53538322448731,
-6.85150814056397,
-19.6524543762207,
-48.8782234191895,
-17.3121032714844,
63.0845451354981,
12.2044210433960,
5.71281719207764,
5.90199947357178,
20.9513130187988,
21.6785068511963,
-22.8770332336426,
32.4259185791016,
0.123525619506836,
19.7375907897949,
29.6075134277344,
-33.4032363891602,
-9.89587593078613,
-37.1175498962402,
-1.55353450775146,
-31.2508277893066,
-57.5372695922852,
1.64321899414063,
-23.3812217712402,
36.5070610046387,
-0.816022872924805,
-23.6290206909180,
-0.880874633789063,
-14.4456377029419,
19.4586105346680,
20.1149711608887,
53.7956695556641,
-31.1794967651367,
-38.1543884277344,
-7.60791397094727,
6.92040634155273,
36.4965972900391,
-49.1568641662598,
2.71070003509522,
-27.2073745727539,
-42.9360046386719,
41.9834938049316,
-46.0905876159668,
-57.0463867187500,
-2.33272457122803,
6.27471065521240,
-21.9090461730957,
-31.2102088928223,
42.1947593688965,
-7.85899448394775,
-14.7226610183716,
8.92553043365479,
6.78477859497070,
45.6868438720703,
-26.8729953765869,
-33.0121765136719,
-6.04981040954590,
23.4592094421387,
4.78470611572266,
16.5539588928223,
33.3730239868164,
-41.7006187438965,
29.6532154083252,
28.2825279235840,
-3.17247724533081,
-27.5522651672363,
-36.4229240417481,
40.0291290283203,
-23.9338493347168,
-61.1332588195801,
13.5403957366943,
-5.90407848358154,
-54.5383148193359,
19.9665756225586,
11.0213289260864,
-8.71481132507324,
-11.6086502075195,
-15.4501428604126,
65.4468841552734,
-25.5557441711426,
-9.61374759674072,
2.92062282562256,
-23.5763969421387,
55.1474075317383,
-30.2816009521484,
-43.9617538452148,
-15.5538311004639,
-29.5327873229980,
-39.8705635070801,
12.1353206634521,
-12.4318914413452,
-78.0723724365234,
-2.90606594085693,
18.8579940795898,
-20.9161262512207,
-44.4365196228027,
-10.1493759155273,
-14.5918292999268,
25.0641441345215,
21.6134872436523,
-32.3402404785156,
1.99641418457031,
12.8097944259644,
37.7832565307617,
14.3227529525757,
-7.48408603668213,
-20.2031211853027,
-24.4080715179443,
-5.15594291687012,
-15.9115152359009,
-27.2472648620605,
-31.3671245574951,
14.9206237792969,
-21.2627677917480,
-6.55288887023926,
60.1053466796875,
13.1953296661377,
37.7679443359375,
8.89146041870117,
-2.49093580245972,
12.7247314453125,
-14.6232414245605,
31.4015007019043,
-16.3197860717773,
-36.7646217346191,
6.58144855499268,
10.6596784591675,
7.97129058837891,
-12.7720499038696,
-31.2231025695801,
-10.3231010437012,
45.2066268920898,
-13.9519414901733,
-51.0609817504883,
30.1287097930908,
19.0452156066895,
-25.8529891967773,
11.4735946655273,
50.1473770141602,
10.1615829467773,
1.33251571655273,
-32.2635154724121,
-41.2033576965332,
42.2407226562500,
-21.6481533050537,
-54.7504844665527,
-35.1263275146484,
-2.74495315551758,
24.1314849853516,
-4.55689048767090,
26.3844909667969,
-31.6759433746338,
2.41124916076660,
32.5436248779297,
-36.1541061401367,
0.503047943115234,
-12.7348918914795,
-0.530218124389648,
13.1492691040039,
0.528887748718262,
-8.11006832122803,
-1.04983329772949,
30.2455253601074,
24.8249626159668,
31.3622703552246,
-2.23982620239258,
9.34848117828369,
3.37858772277832,
-28.8264427185059,
-19.2053184509277,
-20.8314552307129,
-41.1642494201660,
-50.7591514587402,
-13.5631008148193,
-34.3639221191406,
-30.1258964538574,
-16.3568763732910,
-9.52567195892334,
4.98232555389404,
26.7344894409180,
-20.0345878601074,
-39.2171401977539,
35.8039627075195,
-62.4640350341797,
-32.0422325134277,
48.0111846923828,
14.6279687881470,
34.4583129882813,
7.31968975067139,
43.5782623291016,
20.9584541320801,
4.87401390075684,
22.8619461059570,
12.8883533477783,
29.8087940216064,
17.8948364257813,
42.8793792724609,
16.7198085784912,
42.5032043457031,
15.8319416046143,
-30.4468059539795,
6.10447502136231,
32.1590118408203,
3.82578468322754,
-57.1827468872070,
-12.0756120681763,
-4.80479764938355,
29.1022396087647,
41.3867950439453,
12.0662689208984,
20.0769844055176,
13.1709442138672,
21.6622047424316,
22.1150474548340,
6.90410900115967,
9.32903385162354,
0.0907974243164063,
-15.3105154037476,
29.2414932250977,
-2.50089550018311,
20.5202102661133,
52.5976943969727,
-45.2408370971680,
1.87011432647705,
50.1142349243164,
-7.84436893463135,
-41.3853759765625,
36.1731185913086,
45.4373741149902,
-15.0247478485107,
20.6808185577393,
-23.6609382629395,
21.5516204833984,
24.6247863769531,
7.67131423950195,
29.1193199157715,
-14.2429676055908,
43.3346519470215,
50.1366653442383,
36.1266326904297,
32.7284660339356,
-10.8953275680542,
-26.3922958374023,
36.5397300720215,
3.74295425415039,
-40.2449531555176,
63.0459594726563,
2.39188194274902,
-54.6571159362793,
-0.804627418518066,
-17.2518882751465,
4.26871490478516,
-1.72891902923584,
4.61855125427246,
16.6168556213379,
-19.7754688262939,
22.1780433654785,
39.9212074279785,
14.1388664245605,
47.1489944458008,
49.9245452880859,
15.3691425323486,
10.0070457458496,
60.6495971679688,
34.8924713134766,
-38.8207054138184,
-1.70119285583496,
-23.8204460144043,
12.3367824554443,
-6.52261161804199,
-19.3260631561279,
47.1272048950195,
-51.6178932189941,
-0.944289207458496,
22.7677307128906,
-52.6872253417969,
1.94346332550049,
21.4406013488770,
-30.6635742187500,
-7.10663604736328,
7.53863048553467,
-1.75176382064819,
20.5094413757324,
-52.7088279724121,
-38.8073806762695,
-26.0527420043945,
-5.02600860595703,
42.7070884704590,
-8.20325660705566,
20.2202415466309,
10.1371545791626,
-11.9127187728882,
-18.4185123443604,
32.5014953613281,
44.8679885864258,
-23.9222335815430,
-1.86473989486694,
13.9383163452148,
59.2796745300293,
-4.80560493469238,
11.7427339553833,
55.2481536865234,
-13.9368677139282,
-2.23849582672119,
-23.0507545471191,
23.9188346862793,
-42.2959823608398,
-65.4997100830078,
-0.606432914733887,
-42.5942344665527,
0.446158409118652,
-13.6076755523682,
8.04448318481445,
11.1849765777588,
-63.4570236206055,
-29.3209400177002,
36.8784370422363,
41.3860015869141,
-1.07998371124268,
-10.0302381515503,
-24.2500648498535,
-33.9831695556641,
-35.1128120422363,
39.8942375183106,
21.1338958740234,
-70.5517501831055,
8.10389995574951,
18.6767787933350,
-30.9711189270020,
29.2322959899902,
46.5329055786133,
-51.0302162170410,
-6.22970199584961,
44.4058494567871,
36.3994903564453,
-4.78289222717285,
-25.5453834533691,
64.2893829345703,
-22.7016010284424,
-18.7929840087891,
48.8670234680176,
17.0549335479736,
-35.5149688720703,
-25.1176357269287,
42.9220809936523,
-26.1310768127441,
29.7332077026367,
16.7686100006104,
-34.3807220458984,
28.9929485321045,
-49.7020606994629,
-37.3259658813477,
-1.32156801223755,
-1.19631052017212,
35.2614440917969,
4.43530845642090,
7.93348121643066,
-3.79176521301270,
-33.8461074829102,
15.1335926055908,
47.8173217773438,
-31.1600399017334,
-44.3890914916992,
-15.2310447692871,
-20.6156272888184,
4.87797927856445,
-36.4526634216309,
25.3705749511719,
-5.97419834136963,
-51.3890075683594,
14.6851968765259,
-44.4748229980469,
19.6593246459961,
47.5404129028320,
-23.9724311828613,
-33.5614242553711,
4.48028945922852,
-26.1355056762695,
-52.2520103454590,
-19.4972114562988,
-8.71822547912598,
4.03319835662842,
-56.0236625671387,
-44.3028526306152,
-1.91682958602905,
30.9004440307617,
-10.5918855667114,
-50.5454292297363,
-18.0428009033203,
-2.65392971038818,
-2.98665714263916,
-39.8536682128906,
-34.9237709045410,
-42.4439735412598,
-7.28667068481445,
-33.2856750488281,
-56.8116111755371,
-28.7104911804199,
-14.9977064132690,
26.2971210479736,
-53.7308883666992,
-40.3999671936035,
50.0845108032227,
9.56385040283203,
-6.75491237640381,
49.0321960449219,
2.01604175567627,
-62.6561927795410,
37.0797805786133,
8.16158866882324,
-4.05303192138672,
56.1167449951172,
-19.7851314544678,
1.05219554901123,
-7.57212877273560,
22.5501956939697,
2.74555110931397,
-60.9237937927246,
51.5289077758789,
-3.49240398406982,
6.74407100677490,
11.4495887756348,
-26.1098594665527,
64.2650222778320,
13.6137781143188,
31.5789222717285,
-17.8373336791992,
-28.0043907165527,
28.9314842224121,
-38.9838027954102,
32.7619361877441,
-2.24790573120117,
-3.08295154571533,
32.3495521545410,
-36.5438461303711,
27.2396507263184,
-14.4042253494263,
-52.0112457275391,
24.8652267456055,
20.0006752014160,
-26.4899559020996,
-35.6472244262695,
21.5198879241943,
25.4948425292969,
-70.5546112060547,
-9.15803813934326,
38.6563186645508,
-24.2900619506836,
43.9794921875000,
39.1342430114746,
35.4289932250977,
-21.0949020385742,
-61.9123382568359,
-2.03108072280884,
-21.7271308898926,
19.6060352325439,
-53.5712471008301,
-17.9434623718262,
29.8950195312500,
-38.4685630798340,
45.4563255310059,
-24.4511489868164,
8.02609252929688,
6.03716850280762,
-56.6898994445801,
80.7143249511719,
-4.29349708557129,
-31.9870681762695,
39.6347274780273,
0.504595756530762,
4.92128562927246,
4.02736091613770,
12.1759204864502,
33.4960098266602,
-27.0274543762207,
-1.42677211761475,
76.3101501464844,
-24.3154563903809,
3.40428733825684,
56.9963684082031,
-27.3326110839844,
-14.3192758560181,
34.7465591430664,
44.4402580261231,
-28.4803237915039,
-8.86743259429932,
50.4126777648926,
13.9268465042114,
11.4971513748169,
-16.0082912445068,
31.4001655578613,
14.7094392776489,
-30.2494659423828,
21.5074729919434,
8.96322536468506,
-0.197267532348633,
-17.7002544403076,
38.7257919311523,
11.0160303115845,
-52.6465682983398,
-18.6258163452148,
-20.8776397705078,
-24.4147319793701,
-49.2530441284180,
46.9397811889648,
39.7229690551758,
-64.2645339965820,
33.2033538818359,
21.0891380310059,
-12.5654497146606,
49.5120506286621,
21.7542495727539,
9.95328998565674,
41.4137802124023,
53.1824378967285,
9.14665508270264,
-48.0921096801758,
36.6041831970215,
53.6881980895996,
-32.7743415832520,
52.9124832153320,
22.7289772033691,
-71.5595550537109,
-21.2680721282959,
29.4022216796875,
33.1203994750977,
-31.9627532958984,
-0.622879981994629,
22.5535697937012,
-31.1449623107910,
17.7606201171875,
37.9301071166992,
-21.8027992248535,
16.3499412536621,
18.8593254089355,
-35.9336814880371,
-5.50060749053955,
-11.9364662170410,
-19.9628524780273,
-6.03977012634277,
-20.2296276092529,
-48.4677963256836,
-22.8161010742188,
3.43155479431152,
-0.615508079528809,
5.76334857940674,
46.1414794921875,
31.8061447143555,
-54.7700996398926,
49.5206985473633,
57.1279907226563,
-63.8137130737305,
7.91172695159912,
24.9666633605957,
-87.3505096435547,
1.80147933959961,
27.2389373779297,
-29.2295646667480,
21.1274452209473,
-25.4320030212402,
25.9637680053711,
-25.1994152069092,
-17.5892333984375,
58.6633529663086,
0.979346275329590,
-1.50913572311401,
0.548758506774902,
5.82970333099365,
12.0397100448608,
49.9318504333496,
16.1608963012695,
2.40319252014160,
-8.34657669067383,
18.8100585937500,
33.0326232910156,
-1.95733833312988,
-8.56176853179932,
-50.4435997009277,
-6.03763484954834,
-0.722732543945313,
-11.8508052825928,
34.6017494201660,
-13.6665039062500,
-64.2784118652344,
28.1414031982422,
7.70023345947266,
-20.5602416992188,
69.3316345214844,
-24.1718406677246,
-38.3617858886719,
52.5937232971191,
32.9864654541016,
-36.7933883666992,
-50.4432601928711,
56.6589126586914,
-14.8181381225586,
-82.5391845703125,
42.8700103759766,
48.8222045898438,
-2.96915721893311,
-23.2328338623047,
-1.73190832138062,
-3.66417264938355,
9.23748779296875,
26.1709270477295,
-44.2681427001953,
1.42143249511719,
59.5271148681641,
-10.6819381713867,
-65.0926132202148,
4.52362823486328,
-28.6602363586426,
-51.2736854553223,
-20.9703216552734,
-47.3977203369141,
43.6658325195313,
-16.8137664794922,
-19.4864578247070,
1.42643928527832,
-47.8328781127930,
-34.4174804687500,
-29.3555908203125,
43.0761604309082,
5.28135204315186,
-44.9957847595215,
-39.5317802429199,
-8.07061004638672,
2.56335639953613,
3.25698757171631,
-8.69911861419678,
-6.11599540710449,
0.935259819030762,
-40.9688491821289,
-22.1256599426270,
12.0591917037964,
37.1666679382324,
-55.2296409606934,
-47.4748077392578,
30.1329994201660,
-29.2427768707275,
-58.5559043884277,
-21.1384582519531,
40.6256141662598,
24.3117904663086,
6.62584018707275,
-14.0680990219116,
-32.0767898559570,
22.6582031250000,
-30.5496635437012,
-51.1664733886719,
-5.28446483612061,
-55.4729537963867,
-24.5314903259277,
4.35133171081543,
1.85322952270508,
-10.8394336700439,
0.405196189880371,
21.4582824707031,
8.87906742095947,
52.1808471679688,
3.09282016754150,
16.2711524963379,
-13.8511343002319,
-36.4055328369141,
24.2398643493652,
9.60283946990967,
9.25253200531006,
-52.6878356933594,
21.5558300018311,
50.1377029418945,
-1.03972625732422,
39.6628150939941,
10.6178054809570,
0.582652091979981,
4.74025726318359,
-18.9214305877686,
-24.7003688812256,
21.4933471679688,
-27.6994647979736,
-47.0303306579590,
-25.3900966644287,
-30.0823364257813,
13.2048549652100,
-43.5190696716309,
15.8300409317017,
-5.01746940612793,
-52.1192054748535,
38.9153366088867,
24.0593109130859,
18.8884620666504,
-31.8857841491699,
-1.34429454803467,
-19.1941795349121,
4.75358295440674,
49.8900337219238,
-31.5008850097656,
22.2117996215820,
-15.8663215637207,
6.57893276214600,
13.4281682968140,
-17.4799289703369,
37.2973327636719,
-34.5850677490234,
-8.38240337371826,
30.0821475982666,
19.9949073791504,
14.7018718719482,
-26.5699157714844,
7.70063018798828,
15.4899549484253,
4.14202308654785,
48.1772918701172,
31.2619647979736,
-21.9352226257324,
-2.25742673873901,
-15.1139106750488,
-38.6552734375000,
4.75715160369873,
30.3710670471191,
10.4950857162476,
-25.4817657470703,
-31.1392364501953,
-24.2182960510254,
-14.5739345550537,
15.0002317428589,
8.79539585113525,
-36.8314132690430,
-21.2310752868652,
-1.46774768829346,
22.5383605957031,
23.0914039611816,
26.7295455932617,
34.7157669067383,
-31.7397193908691,
21.2681617736816,
63.9782257080078,
-25.7723236083984,
-37.2255973815918,
-5.25285863876343,
-21.6945152282715,
-25.9720191955566,
-54.6580047607422,
-5.08728885650635,
-9.69953536987305,
-25.8177146911621,
36.6834640502930,
-28.6153450012207,
37.0605621337891,
7.43020534515381,
-31.6313476562500,
44.0389099121094,
-27.9479103088379,
-34.5977134704590,
-43.2410507202148,
-7.11612033843994,
35.9647598266602,
16.6731224060059,
-23.9113502502441,
-29.7380332946777,
50.8741035461426,
-21.9674396514893,
-29.7147102355957,
41.8355903625488,
37.5470008850098,
15.6526956558228,
2.31824970245361,
13.3972873687744,
-34.7089271545410,
29.0352840423584,
27.1959686279297,
-1.89276361465454,
-2.64830207824707,
-2.03220939636230,
74.6531677246094,
-55.3443908691406,
2.35837650299072,
46.8401336669922,
-46.0591468811035,
44.8108482360840,
-16.7095069885254,
29.5025501251221,
75.3149871826172,
-45.5080795288086,
-27.4095153808594,
0.404209136962891,
-23.0601005554199,
20.3813476562500,
-28.9369487762451,
-42.3889923095703,
43.1545219421387,
-44.9546508789063,
-40.7438583374023,
-15.3787612915039,
21.8747367858887,
16.5489044189453,
-22.1799354553223,
69.6073913574219,
-7.28081321716309,
-38.0987129211426,
-16.6197834014893,
47.6273574829102,
11.3368167877197,
-69.4535217285156,
14.9312915802002,
-21.3966903686523,
31.6172542572022,
-28.3517646789551,
-19.4428348541260,
30.8986778259277,
-47.0286560058594,
49.4434089660645,
9.60916900634766,
-38.2916259765625,
-20.5000457763672,
27.0066490173340,
-17.2554969787598,
10.9543924331665,
25.7931213378906,
-21.0751953125000,
33.6217498779297,
-44.1523590087891,
55.3927879333496,
16.9016380310059,
-26.3578720092773,
19.9829177856445,
-11.2714557647705,
57.0637245178223,
-35.7932624816895,
3.79723167419434,
7.82279872894287,
-24.6035728454590,
46.8649978637695,
12.3618669509888,
-21.1854114532471,
-32.5767707824707,
-14.0509891510010,
-31.8600120544434,
41.9290390014648,
-11.7235975265503,
-18.5875606536865,
7.26004695892334,
-51.0363922119141,
16.5210838317871,
-34.1193923950195,
21.3670768737793,
38.2111892700195,
15.3784952163696,
-24.9152297973633,
-51.9006462097168,
4.51434707641602,
-39.1645050048828,
-9.14229583740234,
5.29274940490723,
5.47301864624023,
43.7849197387695,
26.7567367553711,
-18.2910690307617,
12.4902820587158,
-6.08962535858154,
-7.54678535461426,
31.1626243591309,
22.5499362945557,
42.3681030273438,
-44.6886520385742,
-21.7159423828125,
33.2886085510254,
-11.6187152862549,
47.0920791625977,
-20.7581043243408,
-43.3895378112793,
34.6057281494141,
-7.06614398956299,
-20.7158699035645,
-12.6800756454468,
32.8179016113281,
8.71592330932617,
-46.4389801025391,
21.6133193969727,
35.4401855468750,
-40.0909271240234,
-58.2030258178711,
20.2319183349609,
26.2267227172852,
-49.4476928710938,
25.3149681091309,
38.3014945983887,
-16.8541870117188,
16.0275287628174,
8.63835334777832,
44.0339202880859,
15.0078029632568,
13.2499179840088,
63.2363815307617,
16.3159198760986,
19.7569789886475,
13.0965938568115,
2.53748130798340,
21.5254726409912,
4.90442466735840,
-1.56165695190430,
5.91134357452393,
30.5176219940186,
-8.73105907440186,
-40.2443847656250,
46.3529510498047,
8.49700736999512,
-32.5576210021973,
16.5839290618897,
-44.7024955749512,
-4.01000213623047,
10.8556051254272,
7.54916000366211,
42.2740859985352,
-40.6751327514648,
2.37806606292725,
-28.7967224121094,
-3.01479625701904,
67.2286911010742,
-4.53322124481201,
35.3041534423828,
53.0057411193848,
13.2226715087891,
-16.3517246246338,
-0.569202423095703,
-29.1539058685303,
-18.0226364135742,
-19.2318572998047,
-42.5393028259277,
17.5559310913086,
-50.9211311340332,
-12.2370395660400,
46.9645500183106,
-32.8128013610840,
-14.9870119094849,
21.1790790557861,
16.2445182800293,
-7.80365848541260,
15.4814453125000,
24.8601570129395,
20.9823055267334,
2.60403251647949,
-41.9979896545410,
56.1366386413574,
10.7994365692139,
-64.8327484130859,
-18.8806610107422,
-27.3088493347168,
50.3782882690430,
-28.2622489929199,
-11.2547206878662,
57.4946174621582,
-74.4725799560547,
-28.6529235839844,
-13.5290241241455,
-34.5420570373535,
8.14386749267578,
39.2273788452148,
42.8558769226074,
-17.2487106323242,
-43.5590438842773,
-6.90924263000488,
23.4447498321533,
3.90615463256836,
8.28482818603516,
39.8264999389648,
30.5136241912842,
-49.5839462280273,
-11.9612426757813,
23.4696922302246,
-55.3518142700195,
-17.1517219543457,
-5.38951396942139,
-3.02260637283325,
2.73245334625244,
-19.6065692901611,
-46.9770050048828,
-25.3036460876465,
49.0782928466797,
-21.2317428588867,
-30.5997085571289,
-25.7047901153564,
-29.2512702941895,
12.3841857910156,
19.7981109619141,
7.96827888488770,
-54.3753623962402,
3.52066326141357,
46.5581893920898,
-21.3162117004395,
-6.08390283584595,
57.3568191528320,
-35.4982490539551,
-42.5055999755859,
36.6090087890625,
-42.4182891845703,
-31.6210060119629,
11.7284221649170,
-11.5040044784546,
-17.7971076965332,
42.9488983154297,
-1.04897880554199,
-57.4004669189453,
54.9446182250977,
5.55272674560547,
-20.4872245788574,
40.4039993286133,
6.10621929168701,
27.5253047943115,
8.00085830688477,
-28.6116428375244,
17.7376918792725,
45.2463455200195,
0.599331855773926,
-16.2123241424561,
-29.7055320739746,
9.25785636901856,
45.2801475524902,
-33.9665985107422,
32.2900657653809,
-17.6415939331055,
-47.1583328247070,
47.7035942077637,
-45.0545463562012,
11.5457801818848,
14.9665288925171,
-53.2726058959961,
35.5754318237305,
38.9318389892578,
-34.2977371215820,
-31.5301780700684,
-10.9422101974487,
1.37564086914063,
3.46327400207520,
-42.7362556457520,
36.1667098999023,
-5.70917415618897,
-32.1701354980469,
33.9414253234863,
-42.3246650695801,
-8.29255580902100,
-10.3580455780029,
12.0025930404663,
14.9074449539185,
-10.4503469467163,
1.83579730987549,
-45.2334289550781,
24.8799629211426,
43.4090232849121,
32.4460754394531,
13.5153951644897,
46.7707710266113,
26.1346931457520,
-39.0300483703613,
32.4746818542481,
7.64878654479981,
1.40600967407227,
-27.9153938293457,
13.1298227310181,
-9.59276390075684,
-43.6999015808106,
29.2427444458008,
-32.8251457214356,
-21.3701267242432,
-45.8926620483398,
-30.1732482910156,
34.4911766052246,
9.13564109802246,
-12.0074472427368,
-28.4075889587402,
-8.66782093048096,
55.3301391601563,
-9.10259532928467,
-14.5113258361816,
14.8000259399414,
-41.8778343200684,
41.2473640441895,
13.4172801971436,
10.8000583648682,
-14.5561809539795,
-70.4556274414063,
6.94230461120606,
-10.8605566024780,
-22.2658100128174,
29.1576652526855,
-21.7678527832031,
8.95550346374512,
32.9665031433106,
-35.8621978759766,
54.0456619262695,
-8.04878234863281,
-15.9325618743896,
26.8672904968262,
1.63405799865723,
26.0339183807373,
12.5212392807007,
39.6678504943848,
46.6117897033691,
12.4970664978027,
-6.53961658477783,
55.9069633483887,
-8.39666557312012,
7.56650352478027,
39.4651794433594,
-45.1274490356445,
-23.0087642669678,
-4.28463125228882,
8.61612606048584,
-32.7095680236816,
-31.3922615051270,
4.61315345764160,
17.3665008544922,
-3.33962106704712,
-14.3742904663086,
41.0185317993164,
14.8190135955811,
-15.6392545700073,
11.5090694427490,
24.1720314025879,
-7.50154829025269,
24.1282882690430,
12.5782585144043,
-25.7379016876221,
52.3108749389648,
1.44271564483643,
-41.7301330566406,
24.0589141845703,
43.1971282958984,
23.6405754089355,
-10.4054384231567,
19.0907001495361,
27.5220699310303,
-36.5261344909668,
-40.5960197448731,
-2.90691757202148,
-25.5891380310059,
4.25349330902100,
-3.95526027679443,
-44.7756614685059,
-1.17618179321289,
-20.3605861663818,
-8.23593521118164,
-18.6384887695313,
-36.7938995361328,
-3.73406887054443,
-37.6535720825195,
-14.5376663208008,
-17.6703872680664,
-11.9394254684448,
75.8779907226563,
-11.2002267837524,
-46.6072235107422,
44.0690383911133,
-3.37451171875000,
18.9043693542480,
7.33411979675293,
-46.0840148925781,
-28.1244621276855,
-50.2324829101563,
-16.3871231079102,
-42.1205825805664,
29.0177898406982,
7.12009811401367,
-41.4714202880859,
39.0241622924805,
-44.4501266479492,
38.3139114379883,
5.94644737243652,
-35.1320953369141,
67.4346923828125,
4.73217582702637,
17.9033565521240,
19.1213684082031,
27.4400291442871,
45.1725234985352,
6.96690368652344,
33.8617744445801,
34.0863265991211,
-11.2754096984863,
28.6810207366943,
45.7195587158203,
43.9587593078613,
2.72826862335205,
-30.0870094299316,
37.3760108947754,
21.5766944885254,
11.1141786575317,
-2.02172183990479,
-6.09511756896973,
37.6551132202148,
51.3106498718262,
-1.49286651611328,
-42.9707794189453,
-28.4300498962402,
-12.4799098968506,
34.8211212158203,
34.8469390869141,
-12.8721351623535,
-32.0132179260254,
24.3344211578369,
-3.12440586090088,
-41.0493927001953,
6.29690551757813,
-6.83233976364136,
8.62227249145508,
1.61040878295898,
-20.6918964385986,
-20.8329200744629,
13.0022201538086,
33.9408187866211,
-41.0026435852051,
-8.60965347290039,
29.8768920898438,
6.47022438049316,
-31.0941696166992,
-9.16976451873779,
17.7596893310547,
-49.4072685241699,
6.57541751861572,
58.1243515014648,
35.3098258972168,
-45.9373550415039,
-54.5989341735840,
5.25326061248779,
6.68533897399902,
57.9424057006836,
14.8036756515503,
-27.8136749267578,
-25.2296791076660,
2.52388191223145,
0.682999610900879,
-45.5728912353516,
30.9047889709473,
-31.7912292480469,
-55.1307029724121,
18.1120605468750,
-52.3415794372559,
-17.8899745941162,
-2.88299655914307,
-66.4832839965820,
-29.7825813293457,
-27.9539184570313,
-39.1745452880859,
9.08874225616455,
-10.6754560470581,
-25.3879852294922,
13.5984506607056,
6.12447834014893,
-28.7581329345703,
-22.3636131286621,
3.18235874176025,
10.4986696243286,
30.5249595642090,
-4.50912380218506,
-31.6478481292725,
29.2106895446777,
-0.789901733398438,
-49.7121963500977,
-14.5129671096802,
-17.0736656188965,
53.5104370117188,
9.42566967010498,
-50.4574432373047,
64.1914443969727,
25.1100349426270,
23.2435226440430,
17.4263420104980,
-29.9006614685059,
4.21105957031250,
-8.16520023345947,
-31.7250118255615,
-17.1614990234375,
-14.5912914276123,
-56.6092033386231,
-45.9156188964844,
14.5969438552856,
30.0141029357910,
-20.7167186737061,
-16.1429672241211,
29.0024108886719,
57.9155693054199,
1.90220928192139,
0.696218490600586,
34.0516281127930,
-40.0968856811523,
29.2564125061035,
42.3780860900879,
9.39699077606201,
-23.2470664978027,
-5.38403415679932,
90.0916366577148,
-30.1408576965332,
-14.1821022033691,
1.60690593719482,
-51.9259757995606,
11.7493953704834,
4.15504360198975,
12.9369068145752,
-17.1810245513916,
-13.3863887786865,
-9.12208843231201,
-31.6097164154053,
-26.1507186889648,
-13.1459922790527,
2.39908885955811,
-0.992967605590820,
49.2937545776367,
15.5522174835205,
-48.1739501953125,
-7.05142736434937,
26.1500892639160,
18.1174030303955,
51.2147636413574,
9.93970680236816,
-30.1227607727051,
-44.1949539184570,
-7.57058525085449,
53.6967849731445,
8.59675025939941,
30.8735332489014,
-35.8973350524902,
-54.2721939086914,
-15.4821529388428,
1.85044765472412,
-1.67731809616089,
-55.2922973632813,
8.66478919982910,
44.9730758666992,
30.1442661285400,
16.6490669250488,
45.6765365600586,
-9.70387268066406,
-30.7514286041260,
19.5552501678467,
-23.8916416168213,
-32.4590988159180,
-11.3603916168213,
-12.4355211257935,
-70.0099639892578,
-40.4972305297852,
-1.45367622375488,
-16.6929588317871,
-24.4286918640137,
-12.0208950042725,
18.6737213134766,
-44.1066436767578,
8.13790225982666,
8.31687736511231,
-15.5829753875732,
-13.9671669006348,
-42.6125793457031,
46.5686645507813,
25.5394783020020,
18.6313896179199,
34.7618141174316,
51.0700149536133,
-19.4642715454102,
6.26441860198975,
33.8177032470703,
-38.6567916870117,
-2.12357521057129,
-28.2978096008301,
33.4472427368164,
-33.8867416381836,
-29.1745071411133,
46.7276802062988,
-19.2278442382813,
-45.5541076660156,
-24.0140476226807,
8.60157108306885,
-35.7981300354004,
-1.59801626205444,
-15.5690441131592,
-26.6169433593750,
-40.4251136779785,
-34.4986915588379,
40.6900749206543,
-4.79272699356079,
-1.60709524154663,
-4.51782035827637,
3.20107841491699,
29.0166740417480,
-9.31745433807373,
16.2012290954590,
-4.17468500137329,
-29.2112197875977,
5.39573287963867,
1.22178840637207,
-17.5156116485596,
23.1505775451660,
8.29955291748047,
-47.8140335083008,
19.2766914367676,
-17.3212223052979,
-31.4655494689941,
35.2278747558594,
-56.9865875244141,
13.8743028640747,
27.7449951171875,
-78.6889801025391,
26.7605895996094,
18.4510631561279,
9.41619491577148,
-38.0353622436523,
13.5201740264893,
39.5016632080078,
-57.9303016662598,
43.0782318115234,
-28.8993740081787,
8.61482620239258,
5.51746559143066,
-43.4339561462402,
-31.0445556640625,
-21.9250183105469,
25.4219055175781,
-23.2379016876221,
-17.4123344421387,
-42.1596221923828,
30.0879783630371,
-33.9533691406250,
4.41810321807861,
6.89998054504395,
-63.0787391662598,
77.7221832275391,
-3.25252532958984,
34.5500106811523,
22.4032936096191,
-34.2860870361328,
16.6033821105957,
1.50121021270752,
15.4671907424927,
-26.2195587158203,
19.3989410400391,
24.0273647308350,
13.7626829147339,
25.5464935302734,
-0.630661964416504,
36.7789611816406,
-2.42940235137939,
-35.7252197265625,
8.26539516448975,
43.7863502502441,
18.4266433715820,
-16.6607589721680,
-12.8222494125366,
32.6274642944336,
20.6902732849121,
-6.59288311004639,
25.5891647338867,
-37.4663696289063,
-30.4745979309082,
54.3599739074707,
36.4308090209961,
-13.7141857147217,
-30.9452209472656,
10.7450284957886,
43.4574699401856,
-33.6776733398438,
0.486940383911133,
52.5120124816895,
-53.3236351013184,
9.67542934417725,
3.03512287139893,
-20.1098098754883,
8.59507751464844,
-69.6465225219727,
26.4310703277588,
-6.19122219085693,
-35.1473464965820,
2.16240310668945,
-9.45628929138184,
43.3820343017578,
-41.6424674987793,
29.6868667602539,
62.1105575561523,
-14.8828163146973,
1.87575721740723,
-31.3753509521484,
34.7989807128906,
16.5535583496094,
22.9872741699219,
3.22160816192627,
-42.4458847045898,
46.8859939575195,
27.0339298248291,
-17.6561355590820,
4.19707012176514,
5.51325988769531,
-81.7417373657227,
31.4445476531982,
-2.01228332519531,
-11.7396869659424,
26.8482112884522,
-58.6395111083984,
27.6989994049072,
-43.5858917236328,
35.1586990356445,
-15.5788660049438,
-35.6090164184570,
16.0872001647949,
-13.9424991607666,
63.1968917846680,
3.35838222503662,
-14.0993442535400,
-1.92643356323242,
48.3385925292969,
-6.45772838592529,
3.62674331665039,
24.2166175842285,
33.3343811035156,
12.9386644363403,
-30.2228355407715,
9.73825359344482,
-21.2481002807617,
38.2497253417969,
-25.8359394073486,
-4.51923418045044,
22.6982402801514,
-64.0785827636719,
14.3547592163086,
43.1858940124512,
19.8729057312012,
-20.3813095092773,
-6.22602891921997,
-10.9041891098022,
-24.3232631683350,
19.5924415588379,
-18.4157238006592,
-9.03920936584473,
-39.7674293518066,
-19.0542106628418,
66.1420364379883,
8.70275020599365,
18.2501449584961,
-13.2072877883911,
-3.91477298736572,
44.0153045654297,
-14.7376613616943,
-21.5990867614746,
4.61390018463135,
-0.709488868713379,
-61.6411590576172,
10.5645360946655,
-2.47252368927002,
-47.8012390136719,
65.1596374511719,
-4.32791900634766,
-40.7159957885742,
3.82899856567383,
-2.27170801162720,
-28.1068782806397,
-19.3834381103516,
54.8910369873047,
0.556987762451172,
-42.1024055480957,
-30.1722412109375,
29.7762355804443,
14.0242204666138,
-49.9961013793945,
26.5510864257813,
-5.56898260116577,
-43.3029136657715,
25.5647430419922,
2.39887332916260,
-50.2309494018555,
33.8365173339844,
-11.6908054351807,
-9.02556037902832,
26.8736038208008,
-53.3202323913574,
68.3960113525391,
35.7227172851563,
-48.4534034729004,
2.59946441650391,
22.8756256103516,
17.9905128479004,
21.7637023925781,
-16.5377388000488,
-38.3180618286133,
-13.1247911453247,
-59.4967155456543,
-3.76460075378418,
39.6957092285156,
22.9399490356445,
6.61231231689453,
-3.50984764099121,
3.82229042053223,
9.16445446014404,
37.6911010742188,
-13.0176467895508,
-5.31886959075928,
12.7911863327026,
-37.3080291748047,
42.4653968811035,
46.1749153137207,
12.6563711166382,
12.0789890289307,
2.32400035858154,
36.2463607788086,
-55.2088165283203,
5.31974887847900,
18.1241340637207,
-42.4186248779297,
-2.06603813171387,
-44.6589889526367,
6.33082485198975,
-6.62455463409424,
24.6394729614258,
-0.620700836181641,
-34.3340148925781,
12.3109731674194,
-26.4328041076660,
51.3694686889648,
37.4249420166016,
12.3321943283081,
-12.2006826400757,
-44.8386192321777,
12.4207525253296,
45.7038612365723,
8.92001056671143,
-24.6454124450684,
52.3825035095215,
-12.6105356216431,
-26.2019081115723,
63.7943077087402,
34.0397872924805,
-54.6503410339356,
-37.1388969421387,
47.7052764892578,
-45.1593322753906,
1.76636600494385,
50.1829910278320,
-16.0122127532959,
-41.5962219238281,
-6.72889995574951,
61.9289703369141,
33.4103126525879,
31.6632785797119,
9.85755252838135,
38.3108901977539,
47.2308692932129,
45.7530288696289,
-12.7676916122437,
-14.2477302551270,
1.63489341735840,
-25.5710582733154,
34.9491233825684,
7.68301963806152,
44.1681785583496,
2.22232723236084,
30.8371715545654,
21.8115329742432,
-36.5447769165039,
-9.04117870330811,
-52.7215270996094,
-21.7816429138184,
-34.9059295654297,
73.4911499023438,
0.991043090820313,
-50.1650009155273,
68.3795547485352,
-28.2205276489258,
33.9759368896484,
-17.0022087097168,
-1.59089088439941,
46.9327087402344,
-1.61249971389771,
52.1656265258789,
-31.4908313751221,
20.4859371185303,
-19.3344593048096,
-53.8303680419922,
43.8501014709473,
23.2900810241699,
-22.7179374694824,
-27.4315299987793,
40.2463569641113,
50.7904052734375,
2.01850605010986,
18.0701332092285,
43.9423675537109,
-37.1683502197266,
-44.7510299682617,
3.39227962493897,
-3.35240936279297,
-22.7477645874023,
-9.81206321716309,
-1.94973897933960,
3.56924247741699,
-11.5337982177734,
-39.2623214721680,
-22.5848102569580,
-20.1068954467773,
22.6472702026367,
34.9426956176758,
29.7590484619141,
26.6171836853027,
36.6432762145996,
41.5251235961914,
-5.85767269134522,
1.61718082427979,
36.1751632690430,
-7.79551124572754,
0.459177970886230,
60.2537727355957,
17.8365402221680,
-3.42166137695313,
18.0107345581055,
3.86876392364502,
-68.5776062011719,
9.02267551422119,
15.4214696884155,
-59.4718780517578,
38.7410545349121,
-40.6015815734863,
-36.9202194213867,
46.5800743103027,
10.7431297302246,
-11.2047262191772,
-44.0922317504883,
-30.6801643371582,
-6.53836822509766,
37.5248260498047,
-37.2383651733398,
-27.8926811218262,
56.9386367797852,
14.8494119644165,
13.0711860656738,
-25.6083984375000,
5.77758121490479,
27.7496299743652,
7.28784370422363,
38.2105178833008,
-0.740814208984375,
-35.1501884460449,
-41.9159965515137,
4.53190422058106,
-24.6360778808594,
-47.7457847595215,
35.9245605468750,
37.2441940307617,
10.6412582397461,
19.6956634521484,
30.4910163879395,
-23.2589740753174,
-0.175482749938965,
10.3463382720947,
-5.89346599578857,
40.7074356079102,
-22.2618980407715,
29.8461189270020,
28.1973419189453,
-35.0753364562988,
47.3058395385742,
6.28031635284424,
-0.907672882080078,
1.76585388183594,
-46.9901390075684,
-21.5353279113770,
6.47223854064941,
27.4780445098877,
-1.19655942916870,
-45.4122428894043,
-9.54464817047119,
38.1888885498047,
-38.6323013305664,
32.5904731750488,
13.4935445785522,
-45.4481201171875,
33.8794326782227,
-29.9808597564697,
42.9909744262695,
-6.31382751464844,
-8.82243442535400,
27.2382392883301,
-34.3013610839844,
-15.4429702758789,
-5.84980106353760,
59.7695159912109,
-34.4461059570313,
-11.1656074523926,
61.0335235595703,
-24.8044662475586,
-22.9420185089111,
-21.4710388183594,
-48.4940567016602,
8.57062721252441,
1.84319972991943,
11.3068313598633,
38.1894874572754,
-47.5351409912109,
-26.7784900665283,
27.2660961151123,
34.3810729980469,
-8.15608406066895,
19.7416954040527,
19.8395004272461,
-39.5010643005371,
27.3355560302734,
24.8995914459229,
-3.97505760192871,
22.0337505340576,
-9.08551788330078,
-29.2629909515381,
44.0299835205078,
56.6328582763672,
-33.2937927246094,
-48.4544296264648,
27.3559455871582,
12.2460460662842,
14.6035413742065,
47.3591003417969,
29.3209266662598,
39.9166793823242,
26.0071563720703,
18.4831829071045,
-13.5148019790649,
18.4851646423340,
-19.0136413574219,
-19.9462051391602,
78.4414672851563,
-20.4130954742432,
-54.2919845581055,
-28.6139373779297,
-6.92281818389893,
15.1168346405029,
6.52690505981445,
-34.6268081665039,
-51.4013595581055,
-5.82968521118164,
-61.9561767578125,
33.1507339477539,
12.7689361572266,
-46.6279144287109,
54.9187316894531,
-14.4838485717773,
44.6000976562500,
56.1950683593750,
-29.0410213470459,
-12.4420127868652,
28.6801586151123,
-28.4017219543457,
-19.9148254394531,
41.4690284729004,
-41.9535255432129,
-6.01727294921875,
42.6372947692871,
10.9782180786133,
-14.3977842330933,
45.7345428466797,
12.2002687454224,
2.18750762939453,
14.8397417068481,
-68.3059158325195,
-5.63209819793701,
28.6684112548828,
-17.6762313842773,
-42.0213317871094,
-36.7767791748047,
-43.5513076782227,
25.5890541076660,
-21.3093376159668,
-46.0968933105469,
63.4064025878906,
3.00522899627686,
14.0316247940063,
47.0623054504395,
36.8185462951660,
37.4164733886719,
-43.4194602966309,
-37.8085289001465,
39.7561340332031,
4.93704509735107,
-8.02956485748291,
9.22165203094482,
-41.2868118286133,
-23.5662784576416,
-54.3506736755371,
-8.20001602172852,
45.2287483215332,
-62.1007041931152,
14.1856870651245,
12.0938730239868,
-7.53790283203125,
42.6287345886231,
-16.9533081054688,
-1.17705154418945,
-46.1977348327637,
-25.2539596557617,
14.3707389831543,
-7.95088529586792,
8.28972625732422,
-31.6506843566895,
17.8158245086670,
7.55907344818115,
-17.0292911529541,
43.2983551025391,
-3.96267127990723,
23.1630325317383,
-15.1157436370850,
-12.6136989593506,
58.9632034301758,
-2.83363199234009,
20.5193557739258,
-5.25998163223267,
-24.7167930603027,
-35.7178649902344,
-24.9726448059082,
37.6583061218262,
29.2064170837402,
18.2277679443359,
30.9314613342285,
40.6519737243652,
27.9346008300781,
5.06296253204346,
-14.6150665283203,
56.2733650207520,
-14.4121599197388,
-23.1762619018555,
43.1429252624512,
3.42117977142334,
22.0955581665039,
4.49708461761475,
33.0405502319336,
-20.6682891845703,
30.4864425659180,
47.5533638000488,
-5.02636480331421,
65.0126342773438,
-14.2954149246216,
-6.99744892120361,
24.5807952880859,
45.3775291442871,
24.3787193298340,
11.8779754638672,
0.187497138977051,
-34.9459686279297,
59.3622131347656,
-11.1944217681885,
12.9584875106812,
20.6890220642090,
-25.8771591186523,
1.66348075866699,
-53.4600715637207,
15.4427585601807,
35.8510131835938,
3.42396545410156,
-9.56034851074219,
6.55578327178955,
-1.63712024688721,
46.5483779907227,
-7.28752613067627,
-28.4756946563721,
43.5106391906738,
-48.5859451293945,
53.9851722717285,
39.8214187622070,
-16.9779186248779,
-9.23599720001221,
-35.2814331054688,
18.3820991516113,
-29.1800174713135,
-40.2905426025391,
-9.56729507446289,
-28.9919853210449,
-60.5621643066406,
-29.6766262054443,
-38.6157455444336,
-21.8184223175049,
42.7265853881836,
-28.4476318359375,
-1.75871276855469,
58.6846160888672,
-22.6140232086182,
-32.1102867126465,
26.5182723999023,
-23.8291873931885,
-40.5376052856445,
14.1903562545776,
-22.5163650512695,
36.1411819458008,
-8.28532791137695,
-72.7583389282227,
30.4072132110596,
-41.4743423461914,
-38.8770904541016,
4.53615474700928,
1.25883674621582,
7.47502994537354,
-1.08102416992188,
35.5418815612793,
-36.2434158325195,
-24.1198215484619,
-0.287873268127441,
22.0055313110352,
27.1957874298096,
-41.7691268920898,
38.7830390930176,
26.0784187316895,
43.1671905517578,
44.9947471618652,
-12.1285390853882,
44.9815139770508,
3.02838134765625,
-19.6636314392090,
-15.3414773941040,
-29.4549922943115,
-39.9713783264160,
40.1133003234863,
1.06633377075195,
-53.7623252868652,
-15.9376239776611,
-34.1146926879883,
42.2982902526856,
-53.4711837768555,
18.7406940460205,
22.1566123962402,
-31.7273120880127,
52.9226570129395,
-68.4504776000977,
37.0920944213867,
4.04044055938721,
-60.8791465759277,
44.2373199462891,
8.36837387084961,
22.8088531494141,
35.2860870361328,
-0.715048789978027,
-4.45706224441528,
52.3964729309082,
21.5432281494141,
-52.7461166381836,
-8.60115146636963,
28.5933914184570,
1.31934928894043,
-51.3516654968262,
-34.7108612060547,
30.4304313659668,
-29.4994468688965,
-28.6729316711426,
55.7148017883301,
-22.4058151245117,
-38.1965065002441,
48.7657356262207,
13.0615158081055,
23.4417495727539,
53.9825286865234,
28.8053283691406,
42.2039985656738,
19.4462947845459,
61.8218612670898,
0.371049880981445,
-28.1254043579102,
81.5022811889648,
34.2612304687500,
33.6747436523438,
-9.93873786926270,
-32.9813766479492,
9.34424209594727,
10.0676898956299,
53.7797088623047,
11.2941341400146,
26.1205863952637,
-27.7192840576172,
-18.6048164367676,
65.7172012329102,
-40.3333587646484,
24.9801006317139,
51.0248298645020,
-39.0702056884766,
-27.2863216400147,
-18.1400699615479,
-41.8653259277344,
-33.5795898437500,
-14.0175647735596,
38.6472854614258,
-15.8291072845459,
-55.1103973388672,
39.8225822448731,
-35.6630325317383,
-5.99183130264282,
-23.7611694335938,
-3.06693553924561,
32.1117210388184,
-22.6519279479980,
12.8222713470459,
-51.6236915588379,
-6.45807933807373,
36.2313919067383,
19.8234329223633,
-13.6246013641357,
12.3718662261963,
52.3983612060547,
8.69899559020996,
-26.0191917419434,
26.8410148620605,
17.3341445922852,
-47.8001785278320,
49.7999496459961,
-24.4319915771484,
-43.7649917602539,
34.0894317626953,
-40.4437408447266,
-16.2826461791992,
-3.53426647186279,
-41.9432449340820,
9.77446365356445,
-16.6101646423340,
-32.5408020019531,
24.9714717864990,
-37.9923019409180,
-40.9065475463867,
22.8919677734375,
32.1536865234375,
-26.5312862396240,
-65.5832901000977,
0.731035232543945,
30.9096851348877,
-11.2964057922363,
-53.4443511962891,
5.77630519866943,
-22.9911899566650,
-44.1261215209961,
42.8795318603516,
-22.6874122619629,
8.50687503814697,
3.61595153808594,
-29.6052818298340,
44.1928634643555,
17.7002525329590,
44.6835861206055,
-19.4463901519775,
-46.6155281066895,
-11.2338628768921,
2.93699455261230,
18.3464431762695,
-61.2076339721680,
14.0554742813110,
29.2498264312744,
29.5663833618164,
14.1693267822266,
-53.5700340270996,
0.923803329467773,
7.55640316009522,
24.3363075256348,
5.29692554473877,
12.9777050018311,
-32.3380317687988,
-9.35435199737549,
9.37623691558838,
-62.5729446411133,
-5.48653888702393,
-39.3147697448731,
-9.62610721588135,
-11.8922214508057,
-1.84142351150513,
57.7135658264160,
-50.2193298339844,
-60.1024932861328,
7.48806476593018,
41.0847969055176,
5.95315074920654,
39.2227783203125,
17.5659904479980,
-22.6617126464844,
49.1503753662109,
7.33032321929932,
19.6840553283691,
-3.63964796066284,
-21.4747505187988,
23.8773689270020,
24.7716979980469,
-39.2884292602539,
-9.27665901184082,
47.8830566406250,
-58.8804168701172,
26.2713966369629,
43.2026138305664,
-36.3365402221680,
-31.1335391998291,
-25.4845924377441,
43.6778182983398,
39.7523231506348,
0.581974983215332,
-5.62273788452148,
26.0596771240234,
44.3652801513672,
11.1023674011230,
-40.1505088806152,
-41.7622070312500,
29.0715942382813,
-15.9127140045166,
-47.0232696533203,
29.3819046020508,
-20.5632019042969,
-53.5974807739258,
-51.4798545837402,
-17.5858879089355,
29.3016319274902,
-50.9605407714844,
20.7595653533936,
65.4158554077148,
-2.02705574035645,
18.1690769195557,
15.4707527160645,
51.6832733154297,
12.5504970550537,
33.6985435485840,
9.31345748901367,
-34.0147743225098,
57.8901405334473,
13.6299438476563,
39.4765205383301,
-0.608372688293457,
6.66536521911621,
50.5313644409180,
-21.2473354339600,
3.35695934295654,
-7.69392967224121,
-10.5290422439575,
-52.9881477355957,
-3.28936767578125,
44.7174377441406,
-6.56208133697510,
7.47761440277100,
-16.1150856018066,
-14.3197774887085,
-28.8008823394775,
10.7216348648071,
51.5591888427734,
-32.2720184326172,
-34.8180160522461,
29.5669898986816,
24.0795726776123,
-45.9300460815430,
-43.9616279602051,
51.7054023742676,
0.939262390136719,
-54.3265304565430,
34.5131072998047,
-9.33864974975586,
7.77240371704102,
39.5084037780762,
-27.8787441253662,
31.4653892517090,
26.0155353546143,
24.6775932312012,
-4.42583560943604,
-9.60989475250244,
65.8522491455078,
-9.12950706481934,
40.7471237182617,
27.8163452148438,
-31.0647659301758,
45.3501663208008,
-39.0717620849609,
-55.0515251159668,
-25.2266445159912,
-39.0785980224609,
-41.2358245849609,
-43.1354675292969,
30.8248081207275,
13.7033004760742,
-0.657544136047363,
4.01394176483154,
-30.6752433776855,
-2.04908084869385,
4.92608451843262,
7.01679992675781,
-36.8047485351563,
-12.7631378173828,
67.2527618408203,
21.0533390045166,
20.1862468719482,
21.7702980041504,
-28.5115547180176,
18.0621719360352,
44.2079887390137,
-43.6626548767090,
-12.0272779464722,
57.0952835083008,
-6.70757198333740,
-68.5596618652344,
-2.70837306976318,
57.5962295532227,
-65.7624969482422,
-39.4269104003906,
31.2238426208496,
-55.5327377319336,
16.0547180175781,
67.8042449951172,
-22.4619827270508,
-46.2573165893555,
11.1070413589478,
47.3769149780273,
15.9234209060669,
34.6098403930664,
54.6487731933594,
2.12184047698975,
-19.7013492584229,
31.6250591278076,
45.5458679199219,
-20.9728870391846,
15.6092519760132,
50.1364212036133,
-36.6505393981934,
-1.51355361938477,
-11.9787626266480,
-43.6717681884766,
28.4099693298340,
-43.0738296508789,
-56.7174720764160,
-27.6357650756836,
-55.6793289184570,
-31.6902732849121,
25.7350540161133,
15.7576189041138,
22.1162567138672,
28.9592475891113,
-13.1134662628174,
4.31068897247314,
-32.1821823120117,
28.7870063781738,
13.4968576431274,
-13.1339750289917,
56.4785118103027,
-19.5249595642090,
-22.3359565734863,
42.3940582275391,
31.7707443237305,
-42.7916946411133,
-6.55007266998291,
-8.39825916290283,
-26.9035110473633,
5.56723213195801,
-51.3123893737793,
37.8182830810547,
1.65272235870361,
-52.6880950927734};
