shortreal in[32768] =
'{0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
-4.38911592937075e-06,4.38911592937075e-06,
0.000857615086715668,-0.000857615086715668,
-0.000130425411043689,1.70185739989392e-05,
-0.00294469785876572,0.00207644514739513,
0.000517314590979368,1.76012399606407e-05,
0.00888451281934977,-0.00483433110639453,
-0.00118979322724044,0.000103017773653846,
-0.0161311868578196,0.00776506913825870,
0.00295175332576036,2.91678588837385e-05,
0.0268595926463604,-0.0121033936738968,
-0.00542815960943699,-0.000286702532321215,
-0.0429344065487385,0.0182635802775621,
0.00903866346925497,0.00127281760796905,
0.0665498822927475,-0.0269927643239498,
-0.0118200145661831,-0.00539663946256042,
-0.102336540818214,0.0404747426509857,
-0.00669883098453283,0.0324266813695431,
0.102436713874340,-0.00545950885862112,
-0.0174739174544811,0.00462837843224406,
-0.116872042417526,0.0232486426830292,
0.0690425336360931,-0.0238357298076153,
0.144421368837357,-0.0498520135879517,
-0.297323763370514,0.0632123351097107,
-0.164491370320320,0.00982888787984848,
0.0569290779531002,0.0451888702809811,
0.410083800554276,-0.188530549407005,
-0.263645827770233,-0.163308382034302,
-0.392919868230820,0.294498562812805,
0.248755723237991,0.527588486671448,
0.539202868938446,-0.752772688865662,
-0.0791890770196915,-1.00755190849304,
-1.08938050270081,1.32884073257446,
-0.215780973434448,1.43418073654175,
1.63814187049866,-0.830794334411621,
0.647801756858826,-2.17863845825195,
-2.32431459426880,0.731393396854401,
-1.56910765171051,3.40720629692078,
3.05108094215393,-0.447411268949509,
3.71394872665405,-5.43856191635132,
-5.30884361267090,0.408017694950104,
-18.5073852539063,13.5823020935059,
-26.0687789916992,17.8305664062500,
-28.1438484191895,5.64882326126099,
-27.3125762939453,-3.57323980331421,
-20.3192501068115,9.07210254669190,
-3.06076955795288,28.3982944488525,
16.2501296997070,21.1651439666748,
21.8685855865479,-17.6394557952881,
8.75393104553223,-54.3817596435547,
-8.53807926177979,-55.1090316772461,
-11.0397119522095,-24.6573352813721,
1.02949464321136,4.37941741943359,
13.3652048110962,13.7510213851929,
13.9070215225220,3.96203231811523,
4.06555795669556,-19.4358692169189,
-4.13289737701416,-50.0434646606445,
2.87850165367126,-70.5329132080078,
27.5136985778809,-61.6138153076172,
47.3335075378418,-26.0172405242920,
40.0484199523926,2.96577715873718,
10.2771854400635,2.14516091346741,
-9.71932601928711,-15.2516822814941,
1.37613129615784,-14.6399679183960,
21.4920043945313,10.9131145477295,
15.6205263137817,32.8808593750000,
-15.7349863052368,21.8783817291260,
-35.0897102355957,-19.6480388641357,
-24.3956718444824,-51.8982734680176,
-6.97463178634644,-48.0531120300293,
-8.70646953582764,-18.2234382629395,
-12.2946414947510,3.50951695442200,
12.9963006973267,-2.89965510368347,
57.2841720581055,-22.2843322753906,
77.2303085327148,-24.6693058013916,
50.2490196228027,0.0566104650497437,
2.92156696319580,33.6583976745606,
-23.9154262542725,47.3199920654297,
-20.0616226196289,46.7733306884766,
-5.97481489181519,49.2110786437988,
2.03339838981628,50.7554435729981,
2.69306135177612,30.5889549255371,
-0.108316153287888,-13.7981605529785,
1.29324328899384,-46.2840957641602,
18.7352943420410,-36.4782638549805,
47.7942390441895,-4.14428710937500,
53.8056297302246,7.31033372879028,
15.2749395370483,-2.31932544708252,
-36.8956527709961,4.34524011611939,
-47.5175819396973,29.9348716735840,
-12.7465744018555,27.3365516662598,
12.6147241592407,-25.0556068420410,
-8.91567230224609,-74.2345199584961,
-42.5316429138184,-51.9048118591309,
-26.5903263092041,19.5662117004395,
27.5510616302490,51.9542617797852,
53.4687347412109,9.22649192810059,
28.7906131744385,-52.0507659912109,
-3.69163370132446,-62.5675773620606,
-4.66626405715942,-34.5553359985352,
4.20142698287964,-20.3649253845215,
-6.33035755157471,-27.3562221527100,
-20.2456588745117,-11.4876937866211,
-8.33281803131104,35.9198532104492,
9.35693740844727,68.7326660156250,
-5.61313056945801,45.9990768432617,
-44.1722297668457,-12.0187349319458,
-48.9561843872070,-54.1802940368652,
-2.50499916076660,-59.5849685668945,
37.1852455139160,-42.8602180480957,
18.5480480194092,-26.3473911285400,
-27.9413852691650,-18.9945125579834,
-37.1573448181152,-18.3413562774658,
3.89629125595093,-21.1473903656006,
48.9551849365234,-19.7709445953369,
61.2755432128906,-5.79500436782837,
47.0730171203613,5.51590156555176,
27.8348236083984,-8.94002342224121,
10.5473279953003,-39.5007019042969,
-0.0273989457637072,-58.4990653991699,
7.40352487564087,-50.6911430358887,
32.2767868041992,-28.8785610198975,
48.4044609069824,-8.44538593292236,
34.6210441589356,8.60961151123047,
13.4867267608643,24.7781238555908,
16.8414020538330,31.9543399810791,
36.2639312744141,24.0462989807129,
35.3924751281738,15.9877138137817,
1.10429441928864,18.1870975494385,
-35.2256278991699,16.3131008148193,
-37.8775978088379,-12.1578168869019,
-7.13160467147827,-47.6587066650391,
22.7822074890137,-45.7200775146484,
26.9132480621338,2.92930936813355,
9.40071964263916,51.0101623535156,
-14.7207746505737,54.7210426330566,
-27.1417884826660,22.8161201477051,
-11.9297904968262,-4.77601051330566,
30.1665706634522,-15.3083324432373,
68.0091018676758,-20.0640735626221,
68.0992126464844,-19.4645061492920,
30.9273719787598,-1.86707949638367,
-12.3457040786743,22.0311546325684,
-31.5797119140625,18.0947341918945,
-31.8735599517822,-19.3171215057373,
-29.6625957489014,-43.1945037841797,
-26.9857959747314,-18.6163043975830,
-16.3895149230957,27.7248992919922,
-2.98618698120117,40.7750892639160,
-3.13201212882996,14.7924823760986,
-7.88606548309326,-9.57822418212891,
5.95898056030273,-2.50069618225098,
33.5983734130859,23.8106460571289,
37.3028793334961,41.4497756958008,
-4.82509994506836,42.6442375183106,
-55.0846748352051,33.4928550720215,
-57.6059913635254,9.79997539520264,
-6.49112510681152,-19.7549571990967,
46.0440597534180,-29.1352500915527,
52.9615516662598,-6.98758172988892,
23.3557434082031,18.7935123443604,
-11.7792081832886,21.0396003723145,
-40.8622283935547,13.4913539886475,
-66.6282501220703,21.1762237548828,
-77.6283721923828,26.2149868011475,
-55.9571075439453,-4.23179435729981,
-13.6485261917114,-55.9317855834961,
14.1716871261597,-69.4300155639648,
8.73586559295654,-19.5681648254395,
-9.53743839263916,34.8970184326172,
-18.7843208312988,29.2749195098877,
-25.4863910675049,-17.6775512695313,
-42.6562919616699,-38.4082832336426,
-59.3494606018066,-17.2154083251953,
-45.7973480224609,1.21346795558929,
-0.205030083656311,-8.48309516906738,
42.1709403991699,-21.9156017303467,
53.9113655090332,-17.3996562957764,
40.7770347595215,-11.5123949050903,
24.4410972595215,-23.9305152893066,
11.4643392562866,-33.9880142211914,
-4.19113779067993,-16.4085559844971,
-20.5017833709717,9.69088554382324,
-21.9217262268066,7.05931949615479,
1.00590634346008,-19.0483608245850,
28.7771987915039,-23.9460945129395,
34.2491950988770,3.18482971191406,
10.9558706283569,20.7789306640625,
-20.4599800109863,8.69445323944092,
-29.1962852478027,-1.99883651733398,
-3.00394177436829,20.2738456726074,
31.1015586853027,49.9884757995606,
29.4189205169678,43.1768264770508,
-11.4587583541870,-2.16996383666992,
-44.1469268798828,-44.0053939819336,
-20.7753486633301,-50.5594062805176,
47.2187042236328,-36.5870666503906,
92.9870529174805,-20.8913040161133,
77.8048019409180,-5.04611730575562,
32.6939392089844,6.95841598510742,
10.6222858428955,-5.17940568923950,
16.9489459991455,-39.2432556152344,
14.1535377502441,-55.1126899719238,
-9.41647148132324,-25.0282154083252,
-19.7329063415527,25.4618053436279,
1.11973285675049,53.9027900695801,
26.7054653167725,54.3557052612305,
18.1411037445068,50.8901786804199,
-16.9510936737061,48.1896972656250,
-40.4639053344727,18.3057422637939,
-33.2517242431641,-38.3367843627930,
-11.2994003295898,-72.5606460571289,
7.15167856216431,-51.7928733825684,
14.3057546615601,-11.0955476760864,
9.80239582061768,3.57282781600952,
-5.23140096664429,-6.88323545455933,
-18.4049930572510,-2.53695821762085,
-2.56518840789795,18.3603630065918,
35.8605155944824,23.0923633575439,
56.0335922241211,4.26714420318604,
29.0087852478027,-2.46972060203552,
-21.4559669494629,20.5976715087891,
-51.8498992919922,33.8353347778320,
-52.1152725219727,-0.810570240020752,
-40.7262382507324,-52.2777328491211,
-35.9006271362305,-56.4195404052734,
-36.9305152893066,-10.6171598434448,
-36.1817779541016,25.1636028289795,
-36.2265625000000,5.99644088745117,
-33.9795341491699,-39.4470024108887,
-18.8519153594971,-65.1496810913086,
7.48417711257935,-63.7376976013184,
23.6309871673584,-58.9323081970215,
18.0784645080566,-51.2300910949707,
1.44241058826447,-22.4642581939697,
-19.4191455841064,17.6930294036865,
-45.5572357177734,26.2119960784912,
-62.3404884338379,-13.3392810821533,
-35.5853805541992,-55.4147796630859,
31.0128822326660,-45.9538421630859,
79.2675781250000,4.62320423126221,
55.8786659240723,34.1914100646973,
-12.1378250122070,11.2575073242188,
-40.6799545288086,-32.6628417968750,
-4.35183382034302,-47.1170845031738,
29.0308322906494,-24.3400554656982,
3.00010824203491,-1.00057470798492,
-46.5107116699219,-5.33539628982544,
-43.9417381286621,-22.6494960784912,
14.5774707794189,-27.9222831726074,
57.0981254577637,-13.6681327819824,
45.2847442626953,-0.564868032932282,
15.0569162368774,-4.82756233215332,
13.4653196334839,-25.4282684326172,
30.9633502960205,-43.0845642089844,
26.8818950653076,-39.4383430480957,
2.12143707275391,-21.8590183258057,
-10.1298036575317,-11.3917675018311,
1.17571198940277,-16.4385452270508,
7.50333023071289,-27.7668170928955,
-12.1914529800415,-30.2099323272705,
-35.7882575988770,-26.3712539672852,
-33.7778816223145,-26.6884822845459,
-4.17641735076904,-29.9942550659180,
30.2465991973877,-23.2654914855957,
51.2579879760742,-8.61830902099609,
52.1892547607422,-7.23266315460205,
36.4940261840820,-19.9264907836914,
9.43214797973633,-20.0912170410156,
-16.8643836975098,9.47378349304199,
-29.7300739288330,42.6430435180664,
-33.8567657470703,38.4569435119629,
-39.7887229919434,-2.94017982482910,
-44.5572853088379,-34.2966995239258,
-27.9390144348145,-25.0168209075928,
9.87220954895020,9.61887645721436,
37.8430976867676,34.2591018676758,
21.6681308746338,40.4452819824219,
-25.9141616821289,39.7287826538086,
-61.0189704895020,31.0130443572998,
-53.5990867614746,3.83141183853149,
-22.7159519195557,-31.5245914459229,
-9.36859321594238,-45.0982322692871,
-25.3189525604248,-23.8271121978760,
-42.3138542175293,10.6881971359253,
-30.8088417053223,24.0554733276367,
-0.636928319931030,9.94328975677490,
23.2393016815186,-13.3863048553467,
27.5704765319824,-26.0020885467529,
25.5264854431152,-19.1103057861328,
33.1331443786621,3.15988945960999,
38.2472305297852,31.0171813964844,
15.1840343475342,44.2909126281738,
-41.1996459960938,24.5319957733154,
-89.3054122924805,-15.6574621200562,
-83.8349990844727,-38.5932083129883,
-33.2427787780762,-22.8453159332275,
5.39091539382935,12.8726463317871,
-7.63584518432617,24.4505500793457,
-44.0378646850586,-1.54310333728790,
-37.8247299194336,-36.2280769348145,
23.1665477752686,-43.4158363342285,
78.1962585449219,-20.5252914428711,
77.0092163085938,5.49344396591187,
37.1911239624023,17.4205551147461,
3.62185716629028,18.4340152740479,
-11.6778182983398,18.1659259796143,
-26.3371524810791,19.8872394561768,
-35.4469184875488,25.5581760406494,
-16.8134174346924,32.4775238037109,
21.7851085662842,34.5393333435059,
31.9171619415283,18.4581336975098,
-2.75431537628174,-10.5986862182617,
-27.8525905609131,-31.7279548645020,
-3.10062313079834,-27.9604606628418,
39.3936691284180,-3.79732632637024,
34.6541595458984,21.6534175872803,
-11.7183456420898,35.5174713134766,
-28.3652000427246,36.7869567871094,
13.8303871154785,23.7964706420898,
56.5894660949707,5.73681879043579,
42.4757499694824,3.21064257621765,
-5.82997941970825,29.6584033966064,
-22.6990470886230,63.9391403198242,
-0.951124429702759,67.1399917602539,
7.66995191574097,29.7003536224365,
-16.2471733093262,-21.7739944458008,
-29.4828796386719,-49.3305130004883,
7.44158172607422,-42.0151138305664,
59.1254577636719,-17.9988403320313,
65.2838973999023,2.24506354331970,
26.6255302429199,4.27449274063110,
-5.10177612304688,-16.5269317626953,
0.598963499069214,-42.1703643798828,
21.0046024322510,-41.3320159912109,
17.5110416412354,-13.3227539062500,
-9.49456501007080,5.60841274261475,
-28.0136966705322,-15.4739151000977,
-18.8887557983398,-44.2179832458496,
0.315580487251282,-25.0999946594238,
4.86654615402222,40.1184349060059,
-16.1218948364258,74.2822570800781,
-47.3208770751953,29.8175659179688,
-58.1527862548828,-44.9139595031738,
-34.4165344238281,-58.9867553710938,
0.847067832946777,1.66537845134735,
6.95672416687012,56.3077850341797,
-18.4853324890137,40.6406822204590,
-36.5845680236816,-16.8451614379883,
-12.6403636932373,-38.5915260314941,
37.9157867431641,-2.52029752731323,
64.4161987304688,43.2497253417969,
48.0230751037598,50.8277702331543,
21.3283214569092,31.1080741882324,
17.3854045867920,26.8817405700684,
28.3550968170166,51.5184745788574,
27.7301578521729,68.9201889038086,
12.2689170837402,44.1647262573242,
-0.724178314208984,-9.49781703948975,
-3.67469549179077,-45.1082572937012,
-4.79153394699097,-39.4769172668457,
-6.82104253768921,-10.7644376754761,
8.17210483551025,4.21495819091797,
41.7761917114258,-8.05541038513184,
68.3775711059570,-15.8395385742188,
60.4067764282227,4.68593883514404,
24.4227409362793,34.8541183471680,
-5.44692516326904,41.8500175476074,
-11.0399675369263,21.3592758178711,
-4.57498502731323,7.47426939010620,
-0.718230307102203,21.6823577880859,
4.94607162475586,42.9799957275391,
19.8542156219482,41.1124496459961,
31.3375492095947,19.6625366210938,
20.1040763854980,13.2069549560547,
-12.2101106643677,22.6603183746338,
-38.3305282592773,12.2212247848511,
-39.5497245788574,-35.1758804321289,
-21.2517242431641,-80.8213958740234,
-2.56421756744385,-72.6467590332031,
6.18266820907593,-16.8599720001221,
6.95671224594116,28.8317871093750,
-3.10253095626831,23.0210800170898,
-24.3964843750000,-16.7582225799561,
-37.8212814331055,-50.0165252685547,
-27.6593036651611,-56.2389564514160,
6.23097753524780,-37.3311424255371,
37.1863250732422,-1.14141082763672,
37.4840888977051,40.4815788269043,
8.23232841491699,60.3647384643555,
-16.1430625915527,37.1983032226563,
-4.33002758026123,-7.52104568481445,
34.7118225097656,-27.9728870391846,
59.6390342712402,-6.04049062728882,
34.6977767944336,23.8713092803955,
-21.8243446350098,18.7417697906494,
-48.0555000305176,-19.1150341033936,
-13.0191450119019,-46.4575614929199,
39.4841308593750,-33.4633712768555,
39.6144180297852,1.55412948131561,
-17.7243175506592,24.4130783081055,
-65.2475280761719,24.0965709686279,
-51.2727012634277,12.0861196517944,
-8.75729084014893,-1.18226838111877,
-0.128374218940735,-9.43252658843994,
-32.4193954467773,-10.7910451889038,
-49.2191085815430,0.301748573780060,
-13.6667699813843,10.1586036682129,
39.1824264526367,5.65817832946777,
57.2506713867188,-9.99324893951416,
37.4747276306152,-11.1390018463135,
13.8926410675049,21.1802253723145,
4.82217073440552,60.8323974609375,
-2.05029296875000,63.5091552734375,
-12.7806568145752,17.7920379638672,
-19.2917842864990,-40.2260322570801,
-14.6931095123291,-66.8443832397461,
-5.82478713989258,-49.6007041931152,
5.91636753082275,-12.9296302795410,
23.4635314941406,13.4896125793457,
37.3348999023438,25.0179824829102,
28.4116821289063,36.6392250061035,
-5.02455139160156,57.1361656188965,
-28.3467407226563,70.9660110473633,
-13.2224779129028,52.8207283020020,
12.2013130187988,3.02936744689941,
5.54605627059937,-44.3632583618164,
-24.9425048828125,-56.7881431579590,
-25.9288845062256,-37.6904296875000,
31.4715290069580,-20.4838867187500,
93.4933319091797,-17.3477611541748,
90.8036651611328,-5.14823150634766,
21.3230934143066,21.0861053466797,
-45.7055358886719,36.7620201110840,
-56.9300918579102,21.1693572998047,
-26.4266662597656,-7.72145700454712,
1.06473898887634,-13.2195167541504,
7.84912443161011,5.18935918807983,
4.38917160034180,15.1807994842529,
-6.95699977874756,6.35090160369873,
-30.7264442443848,-0.865526914596558,
-54.8461265563965,2.96133303642273,
-51.0626411437988,-5.09713983535767,
-9.22829246520996,-36.8587760925293,
45.3533363342285,-55.1532287597656,
75.7751693725586,-23.5985984802246,
71.2973709106445,33.4152793884277,
54.2877502441406,58.3327140808106,
43.5073928833008,32.0933723449707,
35.9550514221191,-3.98493719100952,
26.7187194824219,-17.8959255218506,
8.53926467895508,-25.5022525787354,
-10.2172117233276,-49.8315277099609,
-11.3046140670776,-75.5158004760742,
12.0950727462769,-67.7344970703125,
44.7675209045410,-30.5279521942139,
59.6201858520508,-5.87583875656128,
44.9774856567383,-9.43039417266846,
21.5802268981934,-10.7510166168213,
15.5474796295166,13.6960191726685,
17.9665412902832,46.1947746276856,
-0.0878022387623787,49.8167114257813,
-37.6159667968750,16.6090011596680,
-52.3206062316895,-25.4631309509277,
-16.4084663391113,-45.0532608032227,
43.7641143798828,-35.2421379089356,
71.8169555664063,-12.3368225097656,
55.3202133178711,0.314659655094147,
28.0526084899902,-10.6774358749390,
20.0197277069092,-36.8866806030273,
17.8053684234619,-45.3546905517578,
-2.59304976463318,-17.2169208526611,
-32.1393089294434,26.8023910522461,
-36.6536865234375,35.1138610839844,
-5.76242876052856,-2.82280611991882,
33.2730369567871,-46.0771598815918,
40.0139884948731,-44.1786308288574,
12.1019134521484,0.713084697723389,
-22.1552200317383,39.7915420532227,
-34.3067588806152,34.4568595886231,
-17.2237205505371,-1.64802157878876,
9.92430686950684,-34.5344352722168,
20.3383865356445,-48.3815078735352,
11.4288768768311,-46.4577903747559,
1.17621839046478,-34.6535186767578,
-2.14067959785461,-11.9638795852661,
-1.85554242134094,14.3753252029419,
-9.09121990203857,31.5180530548096,
-17.1117725372314,35.6948051452637,
-15.0772037506104,39.9337615966797,
-9.28640747070313,48.3230628967285,
-22.4465637207031,45.8564796447754,
-51.5091552734375,23.3216667175293,
-55.2515754699707,-7.21745061874390,
-10.8298349380493,-15.1723022460938,
43.4935569763184,7.03552150726318,
49.7091331481934,28.0139274597168,
2.35833859443665,24.6748371124268,
-34.4905967712402,3.52762269973755,
-14.5415534973145,-11.1831521987915,
34.0331306457520,-10.2086706161499,
54.5741691589356,-9.91999149322510,
34.8940773010254,-16.7060871124268,
14.4889898300171,-18.2909202575684,
18.8832836151123,-0.0956823825836182,
23.2461471557617,25.6200771331787,
2.51489686965942,28.1710910797119,
-25.8667278289795,-3.86313748359680,
-26.6852512359619,-51.1551513671875,
-1.14610016345978,-74.2970504760742,
19.5289268493652,-51.5282859802246,
10.6526393890381,3.55994915962219,
-18.8446159362793,46.7855873107910,
-42.9492454528809,46.3240394592285,
-39.1508102416992,11.4834556579590,
-6.85609292984009,-19.7605457305908,
32.4875488281250,-21.9916095733643,
42.5794982910156,-10.6821470260620,
6.94010925292969,-12.0435009002686,
-41.7206039428711,-20.8321571350098,
-51.2158393859863,-7.11249542236328,
-14.7567415237427,32.8707351684570,
20.0025844573975,59.7141952514648,
19.4737606048584,45.0470466613770,
9.60366058349609,9.36259937286377,
24.6890773773193,-6.15336275100708,
48.5187568664551,5.71567058563232,
37.1658782958984,10.4509115219116,
-13.5897922515869,-10.8868265151978,
-50.3379478454590,-31.9608039855957,
-32.5783462524414,-24.4381656646729,
13.6331081390381,1.80119442939758,
37.6210975646973,16.8663349151611,
26.6825962066650,14.9989690780640,
-2.49468088150024,17.1180191040039,
-36.2974395751953,23.7122879028320,
-63.1878738403320,11.2988262176514,
-60.7946968078613,-23.7600135803223,
-18.5510139465332,-48.5128059387207,
25.6872043609619,-30.2677669525147,
25.1806888580322,16.5278663635254,
-10.9030199050903,45.1120491027832,
-22.5452232360840,28.5422515869141,
15.1252765655518,-12.6123600006104,
49.3066825866699,-42.2697830200195,
27.1856327056885,-42.7372589111328,
-25.2039146423340,-22.1135730743408,
-31.4729328155518,0.617059469223023,
19.1332244873047,6.74316978454590,
53.8703804016113,-9.66009330749512,
24.8577785491943,-24.8997745513916,
-33.6073036193848,-11.2852106094360,
-55.8306083679199,28.7469749450684,
-27.7176589965820,57.3733367919922,
5.93653964996338,44.2265129089356,
7.94404935836792,1.72164702415466,
-15.0881576538086,-27.7161407470703,
-32.5739784240723,-18.8614959716797,
-29.4551315307617,10.2247819900513,
-11.4953289031982,25.7093524932861,
2.16378641128540,15.7333297729492,
-7.82320499420166,-9.75148391723633,
-38.8384132385254,-27.7725620269775,
-51.9986648559570,-19.4505138397217,
-15.7948160171509,10.4499940872192,
38.0188560485840,34.9922180175781,
44.6334381103516,29.8631515502930,
-7.36408901214600,2.63073301315308,
-50.6690101623535,-13.4416666030884,
-26.3108596801758,-2.02796506881714,
36.5074768066406,14.7849102020264,
55.4450988769531,10.9341802597046,
11.8326730728149,-1.45292687416077,
-34.7305259704590,9.06094837188721,
-38.8524169921875,37.3431587219238,
-28.1945152282715,41.1981887817383,
-40.4917068481445,2.79991555213928,
-59.6004486083984,-37.5813026428223,
-41.7796516418457,-34.0683784484863,
2.78153228759766,0.528551101684570,
23.6602725982666,13.0562734603882,
0.678470134735107,-15.4773960113525,
-27.2880096435547,-40.1452102661133,
-24.0229492187500,-21.7400398254395,
-5.40056467056274,20.5393142700195,
-3.99309372901917,33.4671134948731,
-18.8314933776855,-2.86160469055176,
-23.5450553894043,-48.3966903686523,
-13.4071683883667,-55.0652198791504,
-9.60302829742432,-19.1083793640137,
-18.0270977020264,23.5884513854980,
-28.1188411712647,33.8299217224121,
-32.0325508117676,3.84585165977478,
-29.7207984924316,-43.5942268371582,
-17.2887554168701,-69.8140716552734,
14.5482845306396,-58.4330291748047,
48.7041549682617,-20.1350116729736,
50.5904502868652,22.4689788818359,
6.18664264678955,49.9307708740234,
-45.3101959228516,52.0163650512695,
-50.4160156250000,30.0947761535645,
-10.3080720901489,-3.87466955184937,
27.3944435119629,-28.6123847961426,
32.6929702758789,-21.9012393951416,
21.8820934295654,4.56467485427856,
18.5658111572266,19.8472957611084,
23.1397418975830,17.7763042449951,
22.1777362823486,19.9963016510010,
11.2829608917236,41.4840927124023,
-3.11468100547791,59.3691139221191,
-17.3447341918945,45.0217895507813,
-31.0420131683350,10.1984214782715,
-33.0554275512695,-5.48938322067261,
-18.4424781799316,3.75257730484009,
-5.57493305206299,3.27500748634338,
-15.4769792556763,-26.6677532196045,
-37.2008666992188,-50.3235702514648,
-37.9149551391602,-22.4990959167480,
-16.0560913085938,34.5991020202637,
-7.83947610855103,58.4433364868164,
-22.7097549438477,25.6694030761719,
-28.3769798278809,-16.7100925445557,
3.06738042831421,-21.4140090942383,
41.7672233581543,-3.66485691070557,
39.7481117248535,-5.45623922348023,
2.36249828338623,-31.4972438812256,
-17.2333793640137,-39.6483497619629,
1.32460093498230,-12.3614416122437,
15.7690124511719,18.1609897613525,
-5.60425996780396,13.7686815261841,
-36.0994415283203,-17.2428493499756,
-33.1069946289063,-40.6886482238770,
-3.92829751968384,-43.4720916748047,
16.0515804290772,-38.1265945434570,
19.7465934753418,-33.9446830749512,
28.6594791412354,-23.5236606597900,
45.2473945617676,-7.78796148300171,
43.6877136230469,2.29411745071411,
18.0179805755615,7.21397113800049,
-3.08532547950745,19.6875591278076,
-3.10310053825378,42.9116096496582,
-4.24569749832153,54.5619773864746,
-26.2954139709473,31.9444923400879,
-47.1972389221191,-9.70279693603516,
-35.9508361816406,-29.9044437408447,
-8.26738452911377,-14.2188844680786,
-4.43582630157471,13.8984584808350,
-28.7151718139648,24.3982639312744,
-39.0069160461426,17.3163528442383,
-13.9967479705811,15.6374740600586,
13.1646575927734,27.4689273834229,
-2.99349164962769,34.4472084045410,
-47.4961318969727,15.5745286941528,
-63.2604866027832,-21.7195777893066,
-26.4472370147705,-39.9442062377930,
22.9775924682617,-19.5751495361328,
28.1754093170166,20.2058963775635,
-8.06362342834473,42.8687973022461,
-41.0385665893555,33.4137573242188,
-40.8132362365723,9.63838577270508,
-26.0566902160645,-6.89800548553467,
-25.5662422180176,-13.8632688522339,
-37.1620559692383,-18.4821605682373,
-38.9956283569336,-12.0994024276733,
-29.0560951232910,8.84037399291992,
-23.8641681671143,18.4857368469238,
-22.7582492828369,-12.4126033782959,
-3.80297827720642,-62.4091453552246,
34.6120300292969,-71.0212326049805,
54.3553848266602,-16.5637931823730,
26.1797351837158,46.2214050292969,
-28.0652999877930,49.8834457397461,
-60.5979614257813,0.851349830627441,
-53.0197525024414,-35.5223999023438,
-33.1884269714356,-33.5669898986816,
-20.2866134643555,-30.3128318786621,
-5.83794879913330,-52.5906219482422,
18.4152412414551,-66.4069824218750,
36.6884002685547,-36.4750137329102,
29.5936203002930,6.62232875823975,
12.7623701095581,8.53896331787109,
10.2147893905640,-24.3686103820801,
22.8576908111572,-30.8395843505859,
23.9454383850098,12.2721843719482,
-0.855430364608765,51.2745437622070,
-33.5049438476563,37.7151184082031,
-44.8121986389160,0.588465690612793,
-29.3954925537109,-3.43382549285889,
-5.32181167602539,28.2505302429199,
13.3827838897705,40.4822463989258,
25.5121841430664,6.91979503631592,
35.6918411254883,-29.6581897735596,
44.0388488769531,-30.3138771057129,
34.0125617980957,-9.86004447937012,
-3.67859649658203,-3.42338466644287,
-49.8111000061035,-11.9898796081543,
-62.5250892639160,-7.71102476119995,
-28.0248622894287,17.1008358001709,
20.5744094848633,35.2131652832031,
32.3687705993652,24.9108371734619,
2.54011726379395,-0.469221591949463,
-30.7582550048828,-16.0505447387695,
-36.0804443359375,-14.7475137710571,
-21.8893089294434,-6.64293003082275,
-13.0571393966675,5.45279502868652,
-7.47619724273682,9.24309444427490,
7.06236600875855,-5.64834403991699,
25.0684223175049,-33.9081535339356,
27.9752864837647,-44.1189613342285,
17.1323051452637,-15.8075828552246,
12.8846435546875,33.6081314086914,
21.5777606964111,56.6804618835449,
30.8100643157959,38.5253105163574,
33.9018516540527,7.79669189453125,
40.2116050720215,-0.623613178730011,
47.8217582702637,13.2779130935669,
32.0630683898926,29.8353939056397,
-17.6307792663574,40.0335197448731,
-68.7693557739258,41.1882209777832,
-75.5570602416992,23.6190509796143,
-37.2833213806152,-21.2346897125244,
0.330258965492249,-71.0152511596680,
6.32871246337891,-84.0707015991211,
-3.92595028877258,-50.8393211364746,
-1.65581631660461,-11.2482576370239,
8.38261985778809,-11.0200138092041,
-1.51747107505798,-47.4856719970703,
-27.1437873840332,-74.6070175170898,
-35.4289741516113,-62.2653503417969,
-3.45933771133423,-29.3199062347412,
46.2225990295410,-10.7309255599976,
64.2983779907227,-17.3820285797119,
35.1552047729492,-23.5747203826904,
-6.58615541458130,-4.37498188018799,
-17.3268489837647,30.1399269104004,
4.00029706954956,47.2488632202148,
23.9831848144531,29.6531085968018,
19.4503231048584,-7.02432155609131,
1.77624595165253,-28.4010696411133,
0.394834786653519,-17.7010059356689,
13.2681121826172,7.40170478820801,
4.44045639038086,18.7761783599854,
-39.7613983154297,-1.76846683025360,
-78.0943298339844,-34.9551353454590,
-62.4979171752930,-46.6079940795898,
-2.19208717346191,-23.1090145111084,
37.8353385925293,12.7275753021240,
16.0493240356445,26.7376251220703,
-32.0909919738770,7.04057073593140,
-37.6356658935547,-24.9289398193359,
1.18101429939270,-39.3296623229981,
29.1874523162842,-31.0727329254150,
18.5062713623047,-16.0179080963135,
5.83263063430786,-6.73748445510864,
27.7297344207764,-5.97135305404663,
55.0130996704102,-4.40539264678955,
35.9230079650879,6.45900058746338,
-16.9693679809570,23.4834194183350,
-32.9625511169434,32.8661079406738,
11.2170295715332,19.8743438720703,
55.7486381530762,-6.40053653717041,
41.5184402465820,-14.3378419876099,
-1.42744064331055,8.23735427856445,
-4.14077377319336,33.9920845031738,
40.1349525451660,26.5239162445068,
66.1348648071289,-8.81558418273926,
35.1551742553711,-26.0430431365967,
-11.7531585693359,-1.69335293769836,
-22.9558944702148,31.3074073791504,
-6.69520187377930,32.6191406250000,
-3.97650742530823,2.70526862144470,
-29.5685672760010,-24.2103691101074,
-53.3510322570801,-30.6512088775635,
-46.8685684204102,-23.0860824584961,
-14.9950199127197,-10.5876770019531,
18.8020744323730,1.56959128379822,
40.4706497192383,5.14032888412476,
41.2018928527832,-13.5389118194580,
17.2002048492432,-40.4114761352539,
-13.8796854019165,-42.6516036987305,
-28.6059265136719,-13.4842138290405,
-28.2612991333008,12.3617897033691,
-24.9918422698975,2.99394893646240,
-13.3099174499512,-19.8390617370605,
19.0241127014160,-20.9327850341797,
56.9529228210449,-5.46205902099609,
58.8578224182129,-7.07733106613159,
11.3935852050781,-27.8185195922852,
-38.3283576965332,-28.9469738006592,
-35.7468948364258,7.87103176116943,
3.04919528961182,41.4633407592773,
16.7252082824707,23.1991729736328,
-3.54317188262939,-27.8638725280762,
-8.88204002380371,-52.7052116394043,
23.1353778839111,-29.3886966705322,
49.9141502380371,4.19014167785645,
25.8216609954834,12.5606298446655,
-20.6698246002197,14.3116502761841,
-32.6410865783691,37.6806068420410,
-11.3720855712891,64.5014495849609,
-4.61876821517944,59.0728187561035,
-22.4503536224365,15.3725385665894,
-19.1294879913330,-26.3484649658203,
26.5720157623291,-28.8949489593506,
65.8942337036133,-2.32617282867432,
45.7607612609863,11.7620859146118,
-4.91670846939087,-7.88216829299927,
-21.6479301452637,-38.6822853088379,
-0.313454151153564,-42.0633735656738,
6.63476657867432,-6.02944946289063,
-27.0219135284424,38.4921264648438,
-63.6328887939453,37.4625892639160,
-56.7266159057617,-21.4043350219727,
-15.3293676376343,-73.5657424926758,
20.1217594146729,-52.9314727783203,
29.9167118072510,28.0470104217529,
24.7223796844482,83.2334747314453,
8.77962303161621,62.3957023620606,
-15.9152832031250,9.61745643615723,
-26.0440425872803,-4.00394201278687,
-0.832300901412964,21.2148399353027,
38.3124160766602,27.7947502136230,
40.3224754333496,2.05416679382324,
2.95565414428711,-7.85556411743164,
-27.1001281738281,22.3335361480713,
-10.9797992706299,45.6392021179199,
27.7475128173828,21.1496810913086,
37.1675987243652,-21.2822170257568,
9.77084350585938,-18.5989875793457,
-15.0482902526855,30.4124393463135,
-15.3695926666260,65.4414978027344,
-12.0531454086304,56.9191932678223,
-20.5563755035400,33.7246589660645,
-27.3712234497070,26.4581642150879,
-16.5312175750732,23.8774356842041,
6.53903388977051,4.97411298751831,
32.6505317687988,-14.4878158569336,
58.2646255493164,-10.2655410766602,
77.8703918457031,5.88192224502564,
71.7455596923828,-1.13994479179382,
32.4040946960449,-28.7527885437012,
-9.41330623626709,-49.2092018127441,
-16.7344875335693,-50.9242744445801,
2.88730287551880,-51.2583084106445,
7.58145236968994,-57.0038604736328,
-14.7108154296875,-55.7440071105957,
-28.8459892272949,-40.1461677551270,
-15.4655342102051,-30.1504688262939,
-0.256216317415237,-39.7817420959473,
-8.53956317901611,-51.1520729064941,
-15.0176191329956,-33.7838020324707,
17.6175270080566,-0.124116897583008,
71.5307464599609,20.2221927642822,
89.7524566650391,24.7180900573730,
43.7599868774414,39.6409339904785,
-21.6851081848145,65.7816009521484,
-50.3263702392578,73.0266799926758,
-33.6477546691895,46.7665061950684,
-6.20357704162598,14.2245855331421,
9.09994983673096,10.9147405624390,
13.8100700378418,34.4378280639648,
11.9135894775391,49.8994789123535,
5.44932651519775,44.4320716857910,
-0.693093657493591,28.4114170074463,
-9.74921798706055,8.89800071716309,
-26.8358230590820,-21.4421653747559,
-45.0808753967285,-51.6881942749023,
-36.6975479125977,-53.6309089660645,
11.2233953475952,-25.3490619659424,
64.6989669799805,-2.67944097518921,
70.4014358520508,-10.1748809814453,
22.0067443847656,-25.2376594543457,
-21.0449047088623,-11.2350282669067,
-20.6396446228027,23.9169139862061,
-8.02218914031982,39.5896568298340,
-17.4658660888672,15.6499719619751,
-30.6448287963867,-14.6737270355225,
-6.95357561111450,-15.8519754409790,
38.0108146667481,6.42600297927856,
38.4258842468262,23.2157211303711,
-23.0514068603516,27.1843719482422,
-80.2653808593750,18.6518859863281,
-75.0821685791016,-3.56200957298279,
-34.2261962890625,-36.1551513671875,
-21.4121360778809,-55.1199417114258,
-30.8366222381592,-43.8097457885742,
-9.03116703033447,-19.5467548370361,
47.4974975585938,-7.17691802978516,
67.3772125244141,-7.23103857040405,
9.71710491180420,3.04651117324829,
-63.3335533142090,21.7313117980957,
-67.9162979125977,17.4868450164795,
-6.92122650146484,-12.6038217544556,
40.4061660766602,-21.5229206085205,
28.3359355926514,14.0513057708740,
-12.3211135864258,53.4621009826660,
-34.6233406066895,50.1084213256836,
-38.2606201171875,19.2115097045898,
-43.3454895019531,3.89115643501282,
-40.3939933776856,5.13010358810425,
-10.3069400787354,-12.2264289855957,
26.1515254974365,-43.4562072753906,
35.7130126953125,-36.7393074035645,
16.9478034973145,17.3343238830566,
3.27573752403259,55.6974716186523,
13.7336091995239,24.5751209259033,
30.8220844268799,-31.0348739624023,
30.5694923400879,-31.9374866485596,
12.1491422653198,16.7801322937012,
-6.42603683471680,44.9985771179199,
-19.2082233428955,22.6963806152344,
-24.3360481262207,-2.26930546760559,
-14.8564815521240,7.22478103637695,
1.12505578994751,26.9919185638428,
-2.01401162147522,18.8728103637695,
-30.2118225097656,-6.05358028411865,
-56.1622848510742,-8.28410339355469,
-48.5414657592773,9.57880401611328,
-21.5908279418945,14.5529041290283,
-8.68595027923584,5.93496513366699,
-16.6624870300293,13.4472789764404,
-18.0986328125000,33.4972648620606,
-0.0371239781379700,23.0846157073975,
12.9402360916138,-30.2383365631104,
1.76948428153992,-73.8888244628906,
-9.48955249786377,-68.0441436767578,
2.37730550765991,-39.5771331787109,
18.0218887329102,-36.6462326049805,
7.06239366531372,-58.2741203308106,
-21.5439929962158,-55.7510261535645,
-33.6889839172363,-13.6398353576660,
-26.6822738647461,21.0626640319824,
-25.6776084899902,12.3117895126343,
-30.4237136840820,-16.3478183746338,
-12.7854728698730,-25.9193000793457,
31.5287303924561,-19.0171241760254,
59.4966506958008,-22.9430141448975,
38.6786651611328,-37.6146774291992,
4.13957595825195,-43.1042022705078,
5.98659706115723,-33.4419937133789,
34.3751564025879,-20.2918071746826,
36.5904273986816,-4.63805150985718,
1.56263625621796,20.8274688720703,
-21.8939456939697,44.5315437316895,
-8.97496414184570,34.5815010070801,
10.7900638580322,-11.9335079193115,
4.15128707885742,-54.9388961791992,
-3.39201164245605,-56.6422500610352,
26.2481613159180,-30.2530555725098,
78.2922363281250,-4.48362731933594,
88.9596252441406,16.1406269073486,
39.5426521301270,38.3363647460938,
-17.7231864929199,46.1391258239746,
-26.8780746459961,23.8978309631348,
3.87738013267517,-10.4460725784302,
23.5502986907959,-18.3622112274170,
14.1006708145142,4.44574594497681,
-9.98641872406006,20.1881275177002,
-31.2808399200439,2.96965885162354,
-47.3535881042481,-19.4501266479492,
-60.2302932739258,-15.5551834106445,
-66.5097122192383,1.32806515693665,
-63.8830184936523,-1.57292830944061,
-59.5366973876953,-15.3449287414551,
-55.8621177673340,-15.1511716842651,
-46.1835212707520,-9.04748344421387,
-27.5509185791016,-22.3705215454102,
-10.3484039306641,-48.4584999084473,
5.24572849273682,-42.4026374816895,
32.8488349914551,4.97203111648560,
58.2587051391602,44.4876632690430,
50.0077438354492,36.6451797485352,
2.93808794021606,6.22987365722656,
-37.6129722595215,4.05478096008301,
-22.0970458984375,23.1613655090332,
29.7164955139160,17.6107006072998,
50.8130493164063,-13.5842552185059,
17.5515556335449,-16.5011863708496,
-18.2775459289551,27.8971309661865,
-15.4625110626221,69.4623947143555,
-2.49217438697815,58.3660202026367,
-28.5692062377930,8.34524726867676,
-75.8704605102539,-30.3651695251465,
-74.7966842651367,-43.0184478759766,
-10.0445880889893,-47.4579391479492,
58.1327438354492,-44.4509925842285,
70.5090942382813,-16.9533882141113,
44.6370811462402,28.3317127227783,
36.7636604309082,47.6255722045898,
57.4748802185059,22.5371570587158,
69.9865951538086,-10.0415229797363,
47.9630584716797,-18.3346138000488,
15.5414199829102,-14.3347215652466,
8.69315052032471,-22.8804168701172,
27.6956844329834,-35.2699966430664,
51.4656372070313,-24.9462966918945,
63.1036224365234,7.69302415847778,
53.1178016662598,36.4166526794434,
22.3306045532227,42.7434806823731,
-13.6035108566284,36.8399429321289,
-31.7200889587402,26.0279312133789,
-27.9692401885986,-1.50211429595947,
-15.8317461013794,-34.3270492553711,
-12.9319801330566,-40.2237167358398,
-21.3048171997070,-12.3416938781738,
-27.7731781005859,9.07066631317139,
-34.1788253784180,-7.04557418823242,
-41.1112899780273,-33.4478034973145,
-36.3969726562500,-25.6568222045898,
-2.79694867134094,10.6469507217407,
36.7893066406250,24.3008365631104,
46.2267074584961,0.725301504135132,
25.4483337402344,-15.9363403320313,
9.53204536437988,3.99938249588013,
15.5273132324219,23.0627956390381,
17.7673225402832,-9.44641113281250,
-3.46361660957336,-63.6365203857422,
-23.3048381805420,-67.7525253295898,
-4.71342992782593,-7.55021667480469,
34.5732536315918,45.2573318481445,
44.0809402465820,32.8110389709473,
22.3866310119629,-15.4626789093018,
16.7978801727295,-33.1781349182129,
42.6898765563965,-4.34230470657349,
52.3203506469727,24.2937450408936,
12.6591377258301,15.0446071624756,
-33.5229034423828,-18.2861137390137,
-20.5878524780273,-39.0940475463867,
35.3746337890625,-34.9191207885742,
59.9688072204590,-14.4791774749756,
26.2643394470215,12.7868862152100,
-7.53245353698731,35.1344490051270,
16.3658924102783,39.3956871032715,
67.3746871948242,30.9240608215332,
73.6817550659180,23.2289543151855,
22.7823867797852,18.7291946411133,
-24.6967258453369,9.66091918945313,
-20.3092327117920,-5.04632949829102,
17.2253570556641,-15.3736305236816,
42.4754219055176,-6.73361873626709,
39.2606964111328,10.6851692199707,
27.3053054809570,18.9937648773193,
25.7367115020752,20.6545028686523,
35.0799293518066,24.7775783538818,
43.2358016967773,21.4274635314941,
44.3774566650391,-1.50650000572205,
32.8325195312500,-21.9507141113281,
7.78198480606079,-7.74055290222168,
-20.0414752960205,36.3981132507324,
-31.1574974060059,59.7502059936523,
-20.4425029754639,34.5251350402832,
-5.08939170837402,1.83918845653534,
1.34702670574188,16.2145748138428,
-0.560872077941895,66.5222091674805,
-5.45971775054932,88.2457656860352,
-12.0475521087646,51.6596755981445,
-21.1696434020996,-0.675368010997772,
-22.9244022369385,-15.5462808609009,
-3.90871548652649,2.56861257553101,
26.1354789733887,15.8011646270752,
38.2662124633789,13.1318788528442,
12.7571277618408,17.6535263061523,
-29.2990875244141,38.6073036193848,
-49.0530853271484,49.0040626525879,
-25.6113414764404,29.6411705017090,
21.7393627166748,-3.62519836425781,
49.0307044982910,-19.3156719207764,
29.4920234680176,-9.78602027893066,
-21.4981517791748,0.998028635978699,
-58.0093765258789,-4.44162654876709,
-50.2073898315430,-16.0505752563477,
-11.9267101287842,-16.2761878967285,
13.2155809402466,-8.35906028747559,
5.08508396148682,-4.92691802978516,
-10.1106433868408,-19.0013256072998,
-4.71182680130005,-40.2992439270020,
14.9092006683350,-47.9440269470215,
15.5266456604004,-37.9147262573242,
-9.53879928588867,-25.8424358367920,
-22.7592773437500,-29.0226669311523,
3.65803194046021,-42.2811622619629,
48.1535797119141,-41.4632034301758,
63.7279815673828,-10.9225759506226,
35.7987403869629,30.7310867309570,
0.557502150535584,44.4768142700195,
-0.718612551689148,18.5355453491211,
29.6279850006104,-14.8285284042358,
51.3158569335938,-14.0048122406006,
29.8018932342529,23.6197853088379,
-23.5241489410400,52.4659576416016,
-66.4198455810547,37.6907691955566,
-63.2090148925781,-8.87759876251221,
-18.4738006591797,-43.6082229614258,
24.1407623291016,-43.7539100646973,
22.9238491058350,-27.0504837036133,
-14.8391819000244,-13.8564004898071,
-45.2540206909180,-0.825403928756714,
-42.0329055786133,24.4376106262207,
-23.3121051788330,50.3664855957031,
-17.9863834381104,50.7002487182617,
-19.9954948425293,16.4431114196777,
-6.83922719955444,-22.1378803253174,
23.3351840972900,-26.7085952758789,
34.9005699157715,7.13735151290894,
11.2669324874878,53.9152679443359,
-16.2362022399902,80.9200820922852,
-14.9327802658081,73.2975158691406,
4.14626979827881,39.7852516174316,
3.11527347564697,4.42216491699219,
-26.0380058288574,-6.23359012603760,
-46.7774467468262,13.3498497009277,
-35.1808700561523,40.2480926513672,
-7.21178054809570,46.1931457519531,
5.92783117294312,29.6268997192383,
-2.78379821777344,17.3831863403320,
-19.7209205627441,23.2839374542236,
-34.4456977844238,27.5148220062256,
-47.1500625610352,4.97365713119507,
-51.2343444824219,-32.9795875549316,
-38.8009147644043,-44.6011505126953,
-15.3594188690186,-14.9046707153320,
1.86004602909088,19.9484348297119,
7.29870939254761,18.0235939025879,
12.2554311752319,-15.7422733306885,
17.8152103424072,-34.6690368652344,
12.2896480560303,-12.3922986984253,
-12.6572027206421,30.0680694580078,
-38.5897865295410,50.1514663696289,
-41.4144134521484,31.6893157958984,
-15.3735294342041,-3.52412390708923,
14.5584716796875,-28.1555213928223,
23.1822090148926,-32.9965553283691,
12.6291942596436,-21.7425918579102,
-0.520758688449860,-4.94106769561768,
-2.41947817802429,11.0342044830322,
4.07197189331055,20.6917057037354,
5.11316204071045,18.7607383728027,
-7.06037807464600,3.39435887336731,
-28.4570007324219,-20.2652206420898,
-41.8281097412109,-37.2285232543945,
-41.2386970520020,-33.8872566223145,
-35.4076728820801,-11.5918951034546,
-40.2280883789063,6.74314498901367,
-50.9383544921875,-4.17605447769165,
-44.2233352661133,-37.4546318054199,
-7.38275384902954,-54.8067817687988,
43.8951911926270,-31.0425987243652,
75.1460266113281,18.1036472320557,
67.6292419433594,50.2352371215820,
33.5824470520020,44.9411048889160,
-0.883311271667481,26.6087131500244,
-17.9827308654785,23.4682769775391,
-18.8997650146484,30.3279418945313,
-11.5896797180176,22.1968421936035,
0.348040938377380,-2.06458926200867,
18.5178890228272,-16.0086479187012,
40.4151115417481,-5.72094345092773,
52.2689590454102,8.99064159393311,
36.2746887207031,4.93670225143433,
0.0850623846054077,-8.74186992645264,
-24.5132369995117,-5.98681497573853,
-13.1406116485596,9.35428333282471,
16.9286308288574,10.9461622238159,
32.8560295104981,-8.22699737548828,
20.2887630462647,-23.4091320037842,
1.11815261840820,-10.9070291519165,
-3.19982361793518,12.2999067306519,
-2.86523771286011,13.9280452728271,
-9.21314144134522,-2.78156328201294,
-15.1377372741699,-10.1278867721558,
-4.34926748275757,5.85308837890625,
11.8978643417358,23.3141059875488,
9.28419208526611,22.1425514221191,
-13.2272396087646,9.64553165435791,
-24.6692104339600,9.14690113067627,
-7.77476882934570,28.7254505157471,
13.7279052734375,49.4933242797852,
3.85751175880432,50.2555656433106,
-36.3877296447754,29.2408008575439,
-70.2069702148438,-0.0802018418908119,
-67.7107086181641,-18.9024658203125,
-35.0710105895996,-17.1573638916016,
0.548156619071960,0.391855508089066,
23.8469734191895,17.2352504730225,
29.1129341125488,22.8835716247559,
14.7834224700928,14.9228372573853,
-17.2797622680664,-0.882970154285431,
-52.7946166992188,-18.7083568572998,
-66.9162216186523,-25.5405750274658,
-49.9142990112305,-13.0230474472046,
-20.6580467224121,12.4817590713501,
-5.05419301986694,29.2796554565430,
-5.93179702758789,18.6076202392578,
-7.06660985946655,-9.42801666259766,
1.03614044189453,-29.2445526123047,
6.01875448226929,-28.1494064331055,
1.43041849136353,-14.6922330856323,
3.98413085937500,-8.41939353942871,
25.8241729736328,-13.8453035354614,
49.2761650085449,-28.1931991577148,
37.0000991821289,-43.9425048828125,
-6.01362991333008,-46.5401687622070,
-34.4255561828613,-21.6488456726074,
-23.3767890930176,21.9613647460938,
1.81611061096191,54.5255393981934,
3.54707288742065,52.8890953063965,
-11.1874179840088,25.5830078125000,
-7.08335638046265,-2.06488132476807,
19.0154991149902,-22.4511756896973,
33.1860694885254,-40.3004035949707,
20.6147499084473,-46.9574623107910,
7.59571266174316,-25.9096565246582,
17.0793247222900,23.8426246643066,
26.1996994018555,64.1399536132813,
0.326937198638916,64.3298950195313,
-43.2151718139648,33.9938774108887,
-56.8795242309570,7.92901134490967,
-24.1818504333496,5.33795928955078,
18.7069225311279,12.5162563323975,
35.1996421813965,11.5541191101074,
25.9705371856689,2.86790657043457,
11.4663639068604,-4.94734239578247,
-3.29308700561523,-3.28812861442566,
-26.0979003906250,9.57238578796387,
-48.5484008789063,19.4077720642090,
-54.3143157958984,10.4105377197266,
-45.3202476501465,-21.3703422546387,
-36.5426254272461,-58.3310890197754,
-25.0072937011719,-73.1961746215820,
7.14498090744019,-58.3027572631836,
50.1221733093262,-26.9572544097900,
65.8386840820313,7.71294546127319,
34.8554306030273,46.8955535888672,
-10.2169198989868,71.6745910644531,
-24.4157886505127,57.3381042480469,
-0.0712192505598068,12.0797653198242,
27.5363140106201,-18.9173564910889,
35.4978675842285,-4.11250495910645,
34.6747474670410,27.1212482452393,
36.5654029846191,23.2989768981934,
33.3700942993164,-11.6310214996338,
16.9190273284912,-23.8184032440186,
1.61279785633087,10.5518503189087,
1.61652028560638,41.6130371093750,
4.70993614196777,21.6818523406982,
-3.08328270912170,-19.3640708923340,
-19.3153572082520,-15.4536209106445,
-28.1397762298584,38.9334983825684,
-26.7304363250732,74.1004867553711,
-21.9073543548584,40.4984474182129,
-21.3848934173584,-28.5298500061035,
-18.6331233978272,-64.5842895507813,
-13.6694173812866,-50.3064041137695,
-15.2381439208984,-15.8298053741455,
-13.2913808822632,9.80433845520020,
6.25517463684082,25.8490371704102,
29.8430099487305,30.8103866577148,
26.7711715698242,13.3581628799438,
-2.54627656936646,-21.8795890808105,
-15.2763767242432,-38.6712989807129,
10.5239076614380,-14.6070938110352,
36.3279953002930,20.9577045440674,
17.3512516021729,25.6950187683105,
-24.9528408050537,-3.02474951744080,
-24.2618503570557,-31.9981479644775,
29.3690834045410,-33.6484298706055,
64.8147201538086,-14.9532165527344,
28.3749351501465,1.92640542984009,
-42.0075531005859,10.3675708770752,
-70.7475585937500,18.2270355224609,
-46.0449333190918,22.4648914337158,
-17.8831939697266,25.8189239501953,
-15.0378961563110,32.7876625061035,
-15.3952980041504,37.3828048706055,
3.42640972137451,30.7593517303467,
23.6347713470459,14.5407247543335,
22.8016242980957,10.5539703369141,
11.6244258880615,30.0366458892822,
13.9966545104980,45.0173606872559,
29.2956180572510,21.7638950347900,
34.1499633789063,-29.8231925964355,
18.6608695983887,-59.1129837036133,
2.37206530570984,-41.4995727539063,
-2.43901252746582,-17.2458667755127,
-2.48076963424683,-33.3041229248047,
0.731350541114807,-73.0982742309570,
11.3727245330811,-71.2684249877930,
26.0604972839355,-4.12117671966553,
35.4085578918457,68.9906387329102,
28.0856113433838,77.6123352050781,
9.95355319976807,22.4512462615967,
-3.01797437667847,-25.6311950683594,
-0.444852709770203,-20.1897277832031,
16.1391563415527,16.3513107299805,
36.4628295898438,32.2490196228027,
40.9861106872559,15.2770862579346,
14.7023830413818,-1.61648356914520,
-29.2512054443359,2.70944595336914,
-52.3909072875977,14.9220323562622,
-27.6763286590576,13.4296035766602,
17.5050773620605,-2.45227169990540,
32.6698760986328,-13.0467538833618,
2.74522972106934,-9.24077606201172,
-33.6356239318848,2.75624799728394,
-33.3253326416016,13.1962060928345,
1.87072670459747,24.2072238922119,
30.5908756256104,35.3049697875977,
20.9047870635986,35.7743873596191,
-9.99579048156738,18.3331775665283,
-29.4467964172363,-11.1070384979248,
-20.5448551177979,-28.0283031463623,
5.67417144775391,-10.5886716842651,
24.8987045288086,37.5866737365723,
18.7190151214600,79.0190200805664,
-9.89628219604492,73.9564056396484,
-38.5357246398926,18.2756938934326,
-40.3247261047363,-48.5895843505859,
-14.6567344665527,-76.7417602539063,
5.81767272949219,-52.4423065185547,
-5.66258192062378,-4.60552597045898,
-33.9893875122070,23.4866104125977,
-31.6240539550781,12.1176490783691,
18.7253417968750,-18.7224178314209,
72.5892333984375,-31.2009162902832,
77.2094802856445,-11.6525592803955,
32.3578186035156,19.1369686126709,
-13.8203716278076,21.2409191131592,
-28.1666221618652,-12.4195890426636,
-18.2208862304688,-44.0036354064941,
-9.03746986389160,-36.3204460144043,
-3.81635332107544,-0.776662349700928,
4.36109590530396,18.7271556854248,
5.19895315170288,12.6851606369019,
-12.0064849853516,14.5057411193848,
-28.3296318054199,35.8656692504883,
-17.1860580444336,44.1448287963867,
13.8542327880859,13.8677396774292,
26.2943553924561,-22.6262741088867,
3.88915467262268,-12.3438291549683,
-24.4689483642578,34.7533378601074,
-34.6479415893555,56.6593360900879,
-37.9413833618164,29.4248332977295,
-50.4158439636231,-1.27651381492615,
-59.5291404724121,1.55487227439880,
-33.7068557739258,9.42121791839600,
14.1609191894531,-13.4210653305054,
39.0741653442383,-39.7272071838379,
25.8178710937500,-20.9090461730957,
10.5487327575684,31.5114097595215,
17.2574081420898,54.5352172851563,
26.8213272094727,23.9306201934814,
11.4156951904297,-14.7470684051514,
-15.5976066589355,-18.7973308563232,
-24.2344493865967,-7.83013010025024,
-17.3273601531982,-13.0255088806152,
-18.4655075073242,-19.1716365814209,
-28.6222305297852,5.33174943923950,
-21.2620334625244,36.8068466186523,
15.5269737243652,26.5911483764648,
53.5371932983398,-15.8103828430176,
65.4968185424805,-28.8165149688721,
52.2514190673828,16.6316204071045,
29.7535705566406,68.8358383178711,
-4.88990545272827,66.5496215820313,
-48.9240188598633,22.2770919799805,
-76.7768249511719,-8.98640727996826,
-72.3958969116211,-6.04945611953735,
-46.4716606140137,0.0891063958406448,
-22.2621097564697,-9.89445400238037,
-6.11979818344116,-15.7634410858154,
5.61707210540772,-5.13510799407959,
7.47015523910523,-2.48879981040955,
-11.8170576095581,-25.4737186431885,
-32.9675102233887,-46.8930511474609,
-24.7141323089600,-30.6213169097900,
5.11066293716431,15.4462604522705,
9.87638187408447,45.1947326660156,
-25.1109046936035,24.4219188690186,
-46.5900802612305,-25.8701725006104,
-10.5090236663818,-55.4804992675781,
53.3671989440918,-44.0866165161133,
73.7638092041016,-7.65085029602051,
37.5378112792969,25.2378501892090,
3.73581814765930,34.6643104553223,
12.3796167373657,24.3932476043701,
32.5169448852539,18.2716770172119,
9.90788269042969,25.7403907775879,
-44.2529067993164,29.1187648773193,
-70.7640380859375,4.42041635513306,
-44.5587005615234,-30.8511772155762,
-3.21618652343750,-30.6728725433350,
12.5305137634277,13.8736572265625,
9.73353004455566,54.3880577087402,
12.5230398178101,35.5591049194336,
19.1052589416504,-31.7596855163574,
11.7976436614990,-80.5308761596680,
-6.30032920837402,-72.5720443725586,
-9.58017158508301,-37.8171501159668,
15.2078094482422,-14.2633514404297,
45.5314750671387,-1.31231594085693,
47.9644317626953,17.7353744506836,
23.5051403045654,38.5674743652344,
-4.49685382843018,48.1994781494141,
-17.9043922424316,48.3485488891602,
-11.3958187103271,47.1729316711426,
7.10220432281494,32.4463920593262,
15.4268274307251,-7.63305616378784,
3.81789112091064,-43.2899208068848,
-12.8759346008301,-31.6979007720947,
-9.09273910522461,12.3685302734375,
15.4624691009521,20.9850711822510,
27.4885807037354,-30.6019058227539,
8.02146053314209,-70.5861740112305,
-16.7113456726074,-29.2884445190430,
-6.96144866943359,48.4182662963867,
22.3906383514404,63.8026008605957,
21.1157417297363,-3.55952310562134,
-14.8636875152588,-65.2340927124023,
-28.4153938293457,-47.5472030639648,
6.69268894195557,16.2766761779785,
41.5525360107422,47.3804397583008,
13.5434522628784,28.6907176971436,
-55.8215599060059,7.78896427154541,
-91.8085327148438,3.76543474197388,
-67.0915222167969,-1.50568580627441,
-26.2605895996094,-16.8376159667969,
-10.7622280120850,-17.4404544830322,
-1.84010803699493,0.467583298683167,
28.0889472961426,7.55999660491943,
55.9720916748047,-9.77008056640625,
44.4971084594727,-23.0525321960449,
7.70065402984619,-10.0942945480347,
-7.54863882064819,14.7886762619019,
11.6076602935791,20.9033412933350,
31.5912113189697,15.3642673492432,
23.7388992309570,25.9356040954590,
-4.30066537857056,43.4520034790039,
-33.2305870056152,27.5972347259522,
-53.4515762329102,-21.3875255584717,
-54.2022705078125,-56.3181076049805,
-21.0475540161133,-50.7343559265137,
33.8315620422363,-32.6917381286621,
66.4378280639648,-34.2763328552246,
38.6751861572266,-41.4684715270996,
-18.1812419891357,-22.5646247863770,
-39.6068572998047,7.21086883544922,
-8.63964843750000,0.858620762825012,
26.6693134307861,-49.3237342834473,
22.2563896179199,-91.8366699218750,
-11.8385114669800,-75.6277313232422,
-30.8940792083740,-19.8911552429199,
-16.6903533935547,15.1036357879639,
4.89609241485596,4.93399572372437,
2.33567333221436,-22.7399044036865,
-18.6385955810547,-29.5131759643555,
-26.7526187896729,-12.5246448516846,
-3.35565090179443,7.72018337249756,
41.7063789367676,16.9962081909180,
71.8249053955078,21.0836429595947,
62.1647033691406,34.3209304809570,
20.7678012847900,49.8468704223633,
-17.2757759094238,47.6373443603516,
-22.3445701599121,15.9385166168213,
-5.27982425689697,-28.0894145965576,
4.62515354156494,-52.7928886413574,
-3.59587407112122,-38.7546653747559,
-10.1941070556641,-1.19098067283630,
2.05865955352783,24.3967666625977,
18.3387622833252,26.0986022949219,
7.35371541976929,17.2472305297852,
-28.9970455169678,11.2438163757324,
-50.6642227172852,5.02495479583740,
-29.0033950805664,-1.97947072982788,
14.3137893676758,-0.404771327972412,
35.1296501159668,15.6352796554565,
15.7298555374146,28.8855876922607,
-14.5151672363281,18.5998115539551,
-19.6072311401367,-5.86423015594482,
-2.47778654098511,-9.72481441497803,
12.2574253082275,17.3617534637451,
7.61322402954102,41.7811317443848,
-10.5645694732666,37.1429405212402,
-28.1958999633789,19.9097938537598,
-32.8374633789063,20.2076511383057,
-18.0252189636230,24.9422016143799,
6.59803009033203,4.68071174621582,
17.4714431762695,-34.4987945556641,
-1.18067741394043,-52.8940200805664,
-25.2348899841309,-36.2874526977539,
-15.7637901306152,-23.2353115081787,
25.2197399139404,-38.9121017456055,
53.7326927185059,-48.6203269958496,
34.5337677001953,-11.8526229858398,
-9.04504585266113,42.6152572631836,
-22.6860294342041,47.2412376403809,
1.99167668819428,-3.50578069686890,
24.6148738861084,-41.1044349670410,
15.7824821472168,-22.9333057403564,
-7.48846054077148,5.20505046844482,
-13.0395059585571,-11.0334014892578,
10.0915966033936,-53.0307807922363,
39.5418205261231,-55.4553604125977,
54.0132713317871,-6.78535938262939,
39.6797752380371,35.6204681396484,
3.89660024642944,32.2528381347656,
-26.9639549255371,13.0624771118164,
-26.0545825958252,21.6874294281006,
3.79155874252319,47.1983413696289,
23.1826801300049,51.9049263000488,
2.28680300712585,31.1459674835205,
-36.3179168701172,14.5570735931396,
-45.1166305541992,15.9561243057251,
-17.0784130096436,23.8396606445313,
3.33678674697876,28.7733993530273,
-12.5270557403564,30.8454418182373,
-45.7590751647949,29.4240226745605,
-64.0881118774414,15.2336015701294,
-63.5313186645508,-8.84439182281494,
-63.0571403503418,-21.5052833557129,
-59.0662117004395,-7.22422409057617,
-30.1153507232666,13.1466903686523,
15.6232357025146,22.1981601715088,
38.3820838928223,23.0294914245605,
14.1299304962158,24.9077568054199,
-29.2241878509522,21.6265659332275,
-42.7017059326172,5.70223093032837,
-13.8622932434082,-9.34391021728516,
29.6869850158691,-7.05003595352173,
58.5560379028320,5.47775030136108,
65.3986511230469,2.03086805343628,
49.5523452758789,-18.4756011962891,
16.3990192413330,-26.4603595733643,
-23.0237770080566,-5.88285827636719,
-47.7961006164551,8.32698249816895,
-44.3567504882813,-17.8177032470703,
-24.2498283386230,-68.6020355224609,
-7.40771245956421,-91.6430282592773,
-4.32835006713867,-70.1717224121094,
-5.56527519226074,-37.5514755249023,
-3.46167087554932,-26.3144149780273,
0.845201373100281,-29.0960655212402,
6.85475015640259,-16.9704494476318,
10.8133239746094,10.4316902160645,
13.2116365432739,29.7843475341797,
21.1693992614746,30.2742710113525,
38.2220687866211,23.9166889190674,
52.6693038940430,16.1455707550049,
46.9770507812500,-2.75564670562744,
19.6025009155273,-34.6157455444336,
-4.41757869720459,-58.2588806152344,
-4.17987632751465,-54.0990829467773,
8.08038425445557,-34.8169021606445,
2.98622083663940,-23.5520935058594,
-15.5768775939941,-17.5323467254639,
-11.7458219528198,-1.75239646434784,
23.0673217773438,24.5724754333496,
51.1856155395508,32.0918960571289,
42.1419143676758,10.6526031494141,
15.9497079849243,-8.22581386566162,
12.0171880722046,8.52688980102539,
24.8813953399658,42.9464302062988,
15.9724903106689,46.6715927124023,
-17.0620365142822,6.06613302230835,
-28.7236652374268,-35.9408340454102,
8.83082008361816,-33.0005722045898,
52.2985305786133,6.20916271209717,
50.9210128784180,34.0261650085449,
14.1825141906738,19.9981040954590,
-1.79605865478516,-17.1453857421875,
25.9443187713623,-40.1506423950195,
52.2046356201172,-36.0115890502930,
35.0575370788574,-13.0307302474976,
-9.00082683563232,11.7473745346069,
-35.1272125244141,26.7171726226807,
-29.4290866851807,22.7725582122803,
-13.5864238739014,2.61075019836426,
-6.82117223739624,-19.1251525878906,
2.70757555961609,-22.0962600708008,
23.2203941345215,0.500306606292725,
36.7422409057617,33.5293426513672,
15.1940212249756,47.8600692749023,
-28.1797866821289,28.4265270233154,
-49.0913848876953,-10.9724731445313,
-17.8471527099609,-40.4234352111816,
42.1759719848633,-40.0171737670898,
78.7393569946289,-12.2582244873047,
61.9976844787598,19.9444713592529,
16.0004997253418,40.0341300964356,
-15.5734262466431,42.5362129211426,
-15.2376432418823,32.3872032165527,
1.60222482681274,15.3876476287842,
14.9495601654053,2.88352966308594,
22.3392200469971,5.97847700119019,
34.3290824890137,14.6569328308105,
45.5008392333984,14.8333644866943,
36.9278335571289,6.40678930282593,
-3.23243975639343,7.04115962982178,
-54.5284347534180,25.1787776947022,
-79.1491241455078,37.2377548217773,
-58.4464797973633,10.5541400909424,
-16.4808826446533,-40.8404045104981,
8.29164505004883,-66.8692779541016,
-3.41726207733154,-41.5924491882324,
-32.2136878967285,-0.439703226089478,
-43.8849678039551,2.46066141128540,
-28.6962451934814,-30.5056552886963,
-3.77461838722229,-42.4508323669434,
4.78134775161743,3.88853788375855,
-8.68048286437988,66.6307678222656,
-28.2049102783203,79.9317703247070,
-38.1802482604981,36.1568031311035,
-36.3112792968750,-5.25523328781128,
-38.8016128540039,-3.04638981819153,
-53.4861373901367,15.0240087509155,
-61.4591369628906,-0.311780571937561,
-35.7982101440430,-44.1058006286621,
14.5048103332520,-64.2623138427734,
43.9319267272949,-35.8748245239258,
26.9269008636475,-0.895984113216400,
-9.89365196228027,-1.02765238285065,
-20.2188167572022,-17.8918952941895,
0.765910923480988,-9.33245372772217,
13.6024818420410,26.7709465026855,
1.69353294372559,48.5864601135254,
-0.846728086471558,36.1440124511719,
28.4921627044678,18.5191860198975,
50.2215538024902,23.1686458587647,
22.4042167663574,27.8419361114502,
-32.3352928161621,7.19117927551270,
-44.3581504821777,-23.4846534729004,
4.28957843780518,-26.3651752471924,
57.9784774780273,0.402932882308960,
58.2951545715332,16.4824428558350,
23.4441738128662,-2.77819538116455,
-1.51291525363922,-32.0920410156250,
-10.9819316864014,-31.1314239501953,
-26.9664802551270,-4.35567617416382,
-43.5842437744141,13.7923603057861,
-27.9971904754639,8.01007652282715,
13.0304574966431,-2.03858613967896,
23.3660964965820,7.16072416305542,
-23.9262237548828,33.1775245666504,
-76.9312438964844,46.1310272216797,
-68.4361877441406,26.0297698974609,
-14.9561882019043,-12.1422119140625,
11.5493288040161,-30.8745803833008,
-24.2269325256348,-17.8164730072022,
-70.0944976806641,4.78097009658814,
-57.9175987243652,1.37346994876862,
3.45851302146912,-30.9583034515381,
46.5991058349609,-60.5051879882813,
39.4630393981934,-62.1975555419922,
11.4721517562866,-47.2401542663574,
3.37706398963928,-38.2230186462402,
13.3959655761719,-30.8038635253906,
8.64571857452393,-12.9143695831299,
-17.0015048980713,7.97914600372314,
-29.8584194183350,7.11037826538086,
-3.44398665428162,-15.1363668441772,
48.4217300415039,-23.9386711120605,
80.5146179199219,4.71375894546509,
66.8303756713867,48.4383010864258,
22.2065811157227,68.7040939331055,
-10.2949228286743,57.9897308349609,
-6.92658376693726,38.1307182312012,
12.9177198410034,27.1451644897461,
7.45690631866455,17.2305622100830,
-34.0637588500977,-1.18902313709259,
-73.0134124755859,-19.2063274383545,
-60.0952301025391,-14.9823675155640,
0.205504179000855,9.63905620574951,
43.5728874206543,37.6879997253418,
15.9914150238037,46.3751869201660,
-53.6013641357422,29.6620140075684,
-85.7361831665039,-0.720198094844818,
-45.4294700622559,-17.8459796905518,
16.3918590545654,-13.4600524902344,
30.3310890197754,-3.46848535537720,
-8.16024208068848,-7.48342561721802,
-35.2521667480469,-21.0528011322022,
-13.3018264770508,-25.2622013092041,
30.4947490692139,-13.9047098159790,
42.0922737121582,-12.8889398574829,
15.9794616699219,-33.2475585937500,
-8.18124389648438,-48.7624397277832,
0.518362045288086,-25.4058494567871,
33.0467720031738,19.0527019500732,
57.6677093505859,34.2082290649414,
61.7724189758301,8.92246246337891,
47.4789772033691,-9.64089870452881,
24.2141799926758,19.0284976959229,
4.97914314270020,67.5292739868164,
-3.38997793197632,78.1114501953125,
-0.143920540809631,41.0778808593750,
9.86505126953125,3.88677072525024,
20.9129295349121,3.15528464317322,
38.3166732788086,21.5939865112305,
58.3849449157715,27.0654239654541,
62.3426017761231,20.0217170715332,
38.9210166931152,23.8770847320557,
1.08036708831787,35.6053237915039,
-28.4795284271240,37.5453567504883,
-40.4002990722656,25.5312042236328,
-42.6787147521973,18.1571960449219,
-38.6463356018066,22.2414760589600,
-26.1777286529541,28.0484981536865,
-12.5110473632813,28.3852901458740,
-16.6193637847900,34.3533668518066,
-36.9884872436523,46.6227912902832,
-49.6260681152344,44.2124176025391,
-29.8364124298096,15.3506221771240,
9.30487632751465,-16.9074440002441,
32.8908309936523,-18.7016925811768,
25.0518436431885,-3.64954280853272,
-2.59581398963928,-14.4853153228760,
-23.8164520263672,-52.5545654296875,
-24.8857460021973,-71.5196685791016,
-2.14982056617737,-43.0718269348145,
24.0163612365723,-2.84850597381592,
26.0382537841797,-1.79768931865692,
0.921893835067749,-37.4531631469727,
-22.1272830963135,-51.0113067626953,
-14.2380361557007,-12.9297561645508,
9.13563156127930,40.7155838012695,
9.70984840393066,59.8422279357910,
-23.7725811004639,36.9130668640137,
-48.8074302673340,-1.44359731674194,
-32.6699943542481,-24.9922256469727,
3.91580939292908,-19.0629520416260,
21.2188205718994,14.5456571578980,
21.4595508575439,43.6550102233887,
31.0199127197266,32.9940795898438,
45.6904983520508,-13.7852277755737,
34.5549964904785,-41.1048011779785,
-2.17040824890137,-9.56002807617188,
-19.4018421173096,49.9148521423340,
4.20508480072022,60.6227645874023,
27.5345478057861,3.45867037773132,
8.49131393432617,-57.1837806701660,
-28.3468017578125,-67.1962051391602,
-23.2057285308838,-44.5732955932617,
28.0888519287109,-27.0679149627686,
60.5674018859863,-18.6881408691406,
33.5704956054688,-3.02136898040772,
-14.5321817398071,9.67842388153076,
-28.1114883422852,-11.4510507583618,
-6.68017959594727,-50.9273490905762,
9.56978988647461,-59.3483467102051,
2.93828272819519,-29.0904502868652,
-7.52283668518066,-10.0859594345093,
-6.19608402252197,-28.1094474792480,
0.821525216102600,-40.5290489196777,
1.67564797401428,2.71593213081360,
1.30658650398254,66.8488388061523,
3.31315183639526,69.5417098999023,
0.307512402534485,6.68546485900879,
-7.20750093460083,-42.1616058349609,
-4.19720649719238,-18.2680778503418,
10.9320325851440,40.7903709411621,
13.9042139053345,50.1689224243164,
-10.4440908432007,-3.59489727020264,
-39.4148597717285,-54.7100601196289,
-44.2117156982422,-52.8538932800293,
-26.7257270812988,-20.0089969635010,
-11.4818849563599,-8.93077087402344,
-9.38707828521729,-36.7363929748535,
-3.87864518165588,-68.9173202514648,
16.0522632598877,-68.1110763549805,
33.6338081359863,-25.7483501434326,
27.6947650909424,35.5586547851563,
4.73593044281006,74.2661666870117,
-12.5160655975342,63.2831344604492,
-12.1709547042847,12.9746379852295,
-0.371900737285614,-34.6648254394531,
9.29956722259522,-40.3994750976563,
6.16557264328003,-13.7012767791748,
-10.7220163345337,-4.52181911468506,
-23.7331848144531,-32.3465957641602,
-10.3465833663940,-60.0557479858398,
22.4652748107910,-41.7277679443359,
40.3008766174316,14.9204740524292,
23.4524078369141,54.3276290893555,
-7.92504978179932,41.0633392333984,
-11.6799898147583,-0.923603415489197,
14.2041168212891,-29.2724552154541,
33.0018882751465,-34.0534629821777,
21.8462829589844,-32.1858444213867,
1.99721062183380,-29.9191989898682,
-4.90264749526978,-17.6358585357666,
-5.75878381729126,0.672261714935303,
-15.7003736495972,-3.93191170692444,
-22.4728679656982,-36.6753921508789,
-8.18005371093750,-64.3446502685547,
12.7618427276611,-50.7600517272949,
6.16309499740601,-4.83395338058472,
-27.1208782196045,23.6489353179932,
-40.5617256164551,6.04952383041382,
-5.36113214492798,-35.7495994567871,
45.5144462585449,-50.0713005065918,
60.1202049255371,-19.3321857452393,
31.2768096923828,29.2514820098877,
2.78842568397522,53.8429718017578,
5.63114070892334,33.5030326843262,
23.6381149291992,-6.74550628662109,
30.2503681182861,-25.8062877655029,
27.1026134490967,-3.66629147529602,
29.7347640991211,38.2461090087891,
32.6998977661133,59.0303115844727,
18.1430625915527,39.6105690002441,
-7.25739574432373,-0.464471578598022,
-9.65863609313965,-30.9681148529053,
27.6315593719482,-33.4697151184082,
70.0378265380859,-14.9926614761353,
65.5010986328125,10.5639686584473,
13.1024990081787,31.1103210449219,
-33.3729362487793,37.4325256347656,
-30.4661140441895,25.2818565368652,
5.61624765396118,0.525205552577972,
24.8237514495850,-24.1407852172852,
3.34613060951233,-32.0769805908203,
-23.9525070190430,-13.7629356384277,
-20.5666027069092,19.1495780944824,
6.97979545593262,36.4924774169922,
26.0406436920166,14.1030235290527,
16.4759445190430,-29.6470260620117,
-1.85589933395386,-47.3997650146484,
-1.95625603199005,-24.4717960357666,
18.8477783203125,1.63529896736145,
36.5768890380859,-11.0505504608154,
30.4450016021729,-51.4844169616699,
4.96493434906006,-62.8471603393555,
-13.4513254165649,-25.3668441772461,
-10.2123069763184,17.1322822570801,
2.06205415725708,17.7561264038086,
-6.80474805831909,-11.1170063018799,
-44.2056236267090,-22.3840255737305,
-69.9845733642578,-8.72105312347412,
-44.9318313598633,-3.51796221733093,
18.5211811065674,-19.8691139221191,
63.3481178283691,-28.2132530212402,
51.5300025939941,-6.55940532684326,
8.57037258148193,13.9661664962769,
-13.2363090515137,-4.49438524246216,
1.61549103260040,-47.0659255981445,
23.5270023345947,-60.1685409545898,
29.1707553863525,-20.9042396545410,
23.8794326782227,31.7205333709717,
20.0288219451904,51.2192039489746,
17.2762660980225,35.1014328002930,
10.0665063858032,14.0836105346680,
8.65885162353516,2.93646955490112,
23.9957447052002,-2.78509902954102,
43.0862007141113,-4.63030004501343,
43.5131340026856,1.38888669013977,
21.4447402954102,12.3859338760376,
-1.41604363918304,19.3349151611328,
-10.1711626052856,18.4448223114014,
-8.62921714782715,18.1837253570557,
-17.1459045410156,24.8358421325684,
-36.8617324829102,25.8983898162842,
-50.0833129882813,10.6883420944214,
-40.3699417114258,-9.63767242431641,
-12.5164623260498,-13.0703420639038,
12.0444650650024,5.35411500930786,
11.9842948913574,32.5473976135254,
-8.65359020233154,50.8920707702637,
-22.7364501953125,44.1407012939453,
-9.34928798675537,16.3424873352051,
17.6757907867432,-15.4130277633667,
27.5144195556641,-23.5984954833984,
14.9221200942993,0.616729259490967,
4.64446878433228,32.0275573730469,
13.5016736984253,31.8750820159912,
27.3347778320313,-5.52029037475586,
21.6421298980713,-36.7539176940918,
4.34691095352173,-29.3932476043701,
2.07433915138245,1.03042840957642,
21.2660732269287,15.7839584350586,
30.3971939086914,13.4873571395874,
11.5117053985596,24.4276618957520,
-19.2722740173340,54.4303779602051,
-35.4212188720703,68.9499130249023,
-37.7840805053711,40.4518089294434,
-35.4738388061523,-6.95787334442139,
-21.3480377197266,-27.0404129028320,
9.19998359680176,-21.2271518707275,
36.2935714721680,-20.2315406799316,
34.1643981933594,-26.8094043731689,
11.1854524612427,-9.87329578399658,
-3.55918765068054,34.5749435424805,
-3.51292634010315,64.0727233886719,
-17.0524406433105,48.1713600158691,
-49.3526000976563,16.2104015350342,
-60.9205169677734,7.07240819931030,
-31.7995605468750,9.80657958984375,
-3.41454052925110,-9.43789863586426,
-18.4165477752686,-38.6755409240723,
-47.2714233398438,-29.1429080963135,
-33.3920288085938,20.7724685668945,
17.5840320587158,47.3336486816406,
41.7918128967285,5.42008399963379,
11.3175468444824,-54.2795982360840,
-22.6228351593018,-63.3437576293945,
-14.6385946273804,-27.0478019714355,
4.35392236709595,-2.37187218666077,
-15.3433904647827,-14.5069408416748,
-52.2727432250977,-31.1521759033203,
-44.1485404968262,-19.4841403961182,
5.46573066711426,9.95727920532227,
30.8853416442871,27.6635932922363,
5.48052501678467,26.8707637786865,
-18.8560142517090,10.9698095321655,
0.721725702285767,-13.7811536788940,
35.1723289489746,-28.4424228668213,
30.8487110137939,-4.61707305908203,
-0.870165288448334,48.8263931274414,
-11.2002210617065,78.6540298461914,
10.0814285278320,58.3053321838379,
18.9609909057617,27.9670352935791,
-2.30878615379334,32.4962387084961,
-15.3688364028931,50.1662559509277,
5.33662319183350,28.0366077423096,
26.5453910827637,-32.5686187744141,
10.9042186737061,-58.5611457824707,
-21.6650886535645,-13.7061071395874,
-23.9840660095215,51.1262779235840,
6.54291963577271,64.4459609985352,
23.8204441070557,34.6014747619629,
1.61497640609741,19.3717365264893,
-36.2025566101074,33.2399139404297,
-52.2748947143555,36.3317489624023,
-45.5423278808594,7.51132297515869,
-41.3414459228516,-22.4461765289307,
-43.8606185913086,-20.8840332031250,
-34.8995971679688,-1.60080826282501,
-6.99763727188110,5.97547388076782,
22.4104576110840,-1.94832193851471,
36.7574386596680,1.35226500034332,
31.4354343414307,22.7557201385498,
15.2982816696167,44.0727386474609,
-1.15551531314850,53.2127227783203,
-15.7415752410889,56.0248718261719,
-34.1487808227539,53.8470840454102,
-53.7575798034668,32.9713668823242,
-56.0289268493652,-2.04480695724487,
-29.8816375732422,-19.6044692993164,
11.5677108764648,-1.55250620841980,
29.2037696838379,27.4727287292480,
6.47781467437744,29.5872650146484,
-18.5818862915039,5.84992074966431,
-0.309561252593994,-4.51995229721069,
51.5651473999023,14.4271879196167,
69.6685104370117,28.3619480133057,
27.0476150512695,9.12674236297607,
-26.2020244598389,-19.6030158996582,
-35.7280082702637,-14.1057376861572,
-10.5767936706543,22.5625114440918,
0.977624297142029,42.8459854125977,
-10.7005290985107,25.0462684631348,
-5.10018730163574,-4.87904167175293,
32.3265266418457,-11.4479789733887,
60.2651710510254,0.473575562238693,
49.1379013061523,2.96010112762451,
27.0797233581543,-8.71521854400635,
23.5805282592773,-12.6729831695557,
15.1330480575562,-3.51559019088745,
-28.6162548065186,3.44909429550171,
-70.8081130981445,-3.07394957542419,
-42.9317703247070,-18.2004051208496,
43.3594055175781,-28.1270351409912,
85.8114624023438,-22.8487091064453,
28.9612102508545,2.26196908950806,
-53.7236633300781,32.0742568969727,
-57.0482864379883,36.1287002563477,
14.4978971481323,3.98892068862915,
54.4368019104004,-28.2118377685547,
12.5157375335693,-14.7406702041626,
-40.8441619873047,41.7030448913574,
-26.1998748779297,73.2108001708984,
28.4729766845703,34.6458663940430,
41.9954414367676,-36.0579147338867,
-1.75720286369324,-66.2462005615234,
-39.7297439575195,-38.9674301147461,
-22.1249504089355,3.28325319290161,
20.7717323303223,25.7428054809570,
26.6827411651611,29.0512924194336,
-17.2913208007813,23.1967811584473,
-63.6948585510254,8.41522979736328,
-69.0666198730469,-9.44173049926758,
-35.3800926208496,-11.3520889282227,
7.54163885116577,2.82763099670410,
22.4278755187988,-0.172748774290085,
2.14121580123901,-37.9675865173340,
-16.9739742279053,-74.4308776855469,
5.92711687088013,-65.3177185058594,
53.4549751281738,-23.7277011871338,
68.2574920654297,-0.838022768497467,
22.9915332794189,-10.1932964324951,
-32.7953453063965,-7.73954439163208,
-30.6958503723145,23.3681449890137,
19.3980827331543,45.7939414978027,
40.8054771423340,24.5306720733643,
3.64324760437012,-14.4711284637451,
-33.2082481384277,-15.4373331069946,
-9.48552608489990,21.0587711334229,
45.9381484985352,43.7957916259766,
62.3152618408203,26.0256156921387,
22.3261013031006,1.69279801845551,
-20.4173736572266,8.89999008178711,
-29.0644207000732,33.3686561584473,
-26.7415084838867,34.3095588684082,
-44.9585456848145,5.47460842132568,
-65.6741638183594,-25.0305023193359,
-55.0797348022461,-37.7325019836426,
-16.5625629425049,-30.5337104797363,
10.9239091873169,-10.2140007019043,
9.41920566558838,17.1313533782959,
-3.37089180946350,40.1465492248535,
-14.6290855407715,46.1129875183106,
-28.9502601623535,32.4934539794922,
-39.6898231506348,15.1501922607422,
-29.9664764404297,4.71922683715820,
-2.94764542579651,-2.81886458396912,
16.9071884155273,-3.31778597831726,
13.2145767211914,18.5358619689941,
1.98354351520538,50.3369140625000,
10.0189132690430,54.7524452209473,
31.4129047393799,21.9218578338623,
40.4152488708496,-12.0698547363281,
41.2942199707031,-11.6578712463379,
49.8233108520508,7.19024658203125,
62.0798301696777,2.55005764961243,
47.8165473937988,-24.9672470092773,
12.2768783569336,-25.4869651794434,
-3.50110054016113,11.5217380523682,
13.1164331436157,33.5717430114746,
23.7243022918701,4.43450212478638,
-4.70704221725464,-30.4675083160400,
-46.7280387878418,-13.7858152389526,
-51.7212524414063,31.1748886108398,
-14.3562564849854,30.3255290985107,
16.7642803192139,-27.0331859588623,
16.9479618072510,-66.5387268066406,
11.5516901016235,-37.4740219116211,
27.4607295989990,14.4961786270142,
53.8237304687500,22.2704830169678,
69.9326477050781,-2.87882566452026,
74.4411773681641,1.82173645496368,
60.4804725646973,43.2092361450195,
16.2954196929932,58.1272544860840,
-43.2305297851563,20.1289100646973,
-60.8095054626465,-22.9319324493408,
-11.0974073410034,-21.4807472229004,
51.6271514892578,3.18284988403320,
50.7938194274902,4.42059516906738,
-14.4755325317383,-15.8805532455444,
-67.6656417846680,-16.6531677246094,
-61.8600120544434,3.07878947257996,
-36.0567855834961,2.66396117210388,
-27.6997871398926,-30.7787933349609,
-15.2603940963745,-54.4002380371094,
29.1912822723389,-31.9721546173096,
73.7561264038086,5.01224517822266,
65.9806900024414,13.4214248657227,
16.0146961212158,8.21860694885254,
-19.9171733856201,29.5743865966797,
-16.8896045684814,69.0433883666992,
-8.14305973052979,72.4747009277344,
-14.8785343170166,21.8968372344971,
-11.3812112808228,-30.1492309570313,
19.0852451324463,-19.9165496826172,
40.4742813110352,38.9962615966797,
13.4294843673706,76.5307769775391,
-37.3354721069336,53.5627403259277,
-53.4691085815430,-2.22423768043518,
-30.1373329162598,-42.7477111816406,
-7.55521726608276,-42.1631050109863,
-10.3306913375855,-13.1810922622681,
-20.8964900970459,11.5374975204468,
-21.5390319824219,5.23064994812012,
-18.2456970214844,-21.3822898864746,
-14.8766832351685,-33.3602066040039,
-0.668193101882935,-8.75141334533691,
30.8687877655029,25.3042240142822,
52.0791320800781,19.3861770629883,
33.8340492248535,-26.1377124786377,
-3.32855463027954,-54.8027381896973,
-26.0601654052734,-25.9280700683594,
-32.5084114074707,21.7884140014648,
-42.9753341674805,18.6177444458008,
-50.5221481323242,-33.6077804565430,
-28.0957794189453,-68.8752059936523,
16.1309967041016,-44.0006065368652,
36.6870689392090,-0.267433404922485,
11.7366046905518,0.542136967182159,
-18.6332283020020,-35.2508392333984,
-9.61492824554443,-51.2200393676758,
22.6253623962402,-17.4218120574951,
27.1200675964355,29.0031223297119,
2.35915732383728,35.9217758178711,
2.40009522438049,6.24806594848633,
49.2289962768555,-16.9260692596436,
94.0609893798828,-5.56931591033936,
78.5673522949219,25.0355587005615,
16.9828109741211,41.1637039184570,
-31.5580368041992,29.0925064086914,
-31.5255279541016,7.12791728973389,
-5.96177053451538,8.18616104125977,
11.2357721328735,29.8144531250000,
11.7599401473999,35.6129302978516,
7.19166469573975,-0.796052455902100,
2.20861887931824,-52.8401756286621,
-1.39925551414490,-58.7972259521484,
1.58896589279175,2.13177824020386,
7.29760456085205,70.8592453002930,
-1.81565320491791,72.8383941650391,
-30.2905158996582,12.3742790222168,
-51.3342933654785,-37.7902641296387,
-44.5751304626465,-30.1529064178467,
-24.3874874114990,3.75173091888428,
-24.6178359985352,12.4873285293579,
-44.7985534667969,-2.62036871910095,
-52.5800056457520,-2.12914609909058,
-25.4264106750488,30.2737312316895,
8.06613922119141,61.3180694580078,
8.16181087493897,58.3271217346191,
-18.5722751617432,30.0058078765869,
-37.4889678955078,8.59507083892822,
-30.7476711273193,10.8168210983276,
-12.3334207534790,24.1821575164795,
6.86463451385498,27.5086994171143,
28.6975727081299,11.8107833862305,
51.3087539672852,-13.0880203247070,
58.8266296386719,-20.3631706237793,
40.1948242187500,10.6677122116089,
12.8618335723877,52.5801506042481,
-4.53716897964478,53.2882575988770,
-12.9290981292725,0.345860958099365,
-20.4711227416992,-56.8849830627441,
-12.8985052108765,-64.1513595581055,
24.6002044677734,-27.4278182983398,
67.9431915283203,0.647681176662445,
71.9127197265625,-4.42593383789063,
35.2720298767090,-12.0029621124268,
9.48154926300049,5.37897491455078,
27.7845954895020,28.8677768707275,
55.1092529296875,27.3530368804932,
29.5955123901367,9.06381034851074,
-39.8758430480957,3.55070137977600,
-81.3037719726563,14.9028091430664,
-56.0651588439941,24.1731929779053,
-3.45502686500549,23.4754142761230,
13.7649965286255,19.1293010711670,
-2.99694538116455,11.7285652160645,
-14.4785099029541,-4.48763132095337,
-10.3674459457397,-19.9796772003174,
-13.1715526580811,-16.4658088684082,
-32.7593994140625,-0.402075260877609,
-40.8327217102051,-3.58809971809387,
-22.5302200317383,-31.4329414367676,
-1.03183031082153,-41.7665481567383,
-9.16312503814697,-10.6742296218872,
-38.5010299682617,21.1933593750000,
-51.1408615112305,1.55671119689941,
-28.5440101623535,-44.6429710388184,
11.1342887878418,-48.4239273071289,
43.4382133483887,7.14274454116821,
55.5392990112305,53.7788276672363,
39.2410774230957,34.1028671264648,
9.30590057373047,-16.0073146820068,
-5.03844308853149,-23.3286972045898,
12.9596166610718,16.7692794799805,
46.0499267578125,36.9526100158691,
61.6101531982422,4.73613214492798,
48.1894378662109,-37.1922073364258,
23.2726917266846,-39.1642189025879,
3.00371360778809,-9.55721092224121,
-12.5162410736084,14.1531019210815,
-22.3790607452393,25.3441772460938,
-14.5633935928345,43.0813865661621,
3.90698862075806,63.4385185241699,
-3.24040961265564,57.1497230529785,
-39.1946792602539,16.1760673522949,
-59.5496292114258,-26.1050033569336,
-26.1472320556641,-42.1332740783691,
33.5522193908691,-42.6617393493652,
62.2906837463379,-39.2308807373047,
52.1343383789063,-17.2350997924805,
39.2782516479492,29.8856449127197,
40.7006607055664,63.3442802429199,
27.7569656372070,41.8390769958496,
-8.76469612121582,-13.2007522583008,
-29.0887107849121,-37.3026237487793,
-4.01046371459961,-5.99537944793701,
24.2074317932129,29.9585323333740,
1.14531028270721,22.1089820861816,
-53.9150085449219,-3.58292460441589,
-71.7675018310547,4.94806337356567,
-39.4172477722168,44.3735542297363,
-12.2169237136841,51.2961196899414,
-27.1612834930420,1.12318873405457,
-46.4228820800781,-59.0007743835449,
-22.1118221282959,-73.4182739257813,
25.4911537170410,-43.1457710266113,
37.9001464843750,-12.0819053649902,
2.72693204879761,-3.09626007080078,
-29.3142299652100,-5.03374767303467,
-24.6291007995605,-6.23067617416382,
0.700935006141663,-11.8140745162964,
12.8441524505615,-28.5663051605225,
15.2810144424438,-39.7061882019043,
18.8790645599365,-29.8412513732910,
12.0695838928223,-1.38804531097412,
-17.7062988281250,27.4347515106201,
-48.9536895751953,40.7912330627441,
-45.7771530151367,31.4848594665527,
0.700983762741089,10.5618543624878,
50.3069686889648,-3.03282046318054,
57.4791717529297,0.301131695508957,
26.6897125244141,13.6822471618652,
-4.77312898635864,23.8197555541992,
-11.7584466934204,26.8358955383301,
-4.39900064468384,34.8040809631348,
-8.55674648284912,46.2927894592285,
-36.4535331726074,43.2898483276367,
-71.1537094116211,11.8715972900391,
-80.9573974609375,-32.6111450195313,
-53.3899879455566,-57.7823677062988,
-9.56065940856934,-48.6937026977539,
14.7753944396973,-26.8088264465332,
3.59974741935730,-18.1438961029053,
-16.3438377380371,-29.7545108795166,
-4.98877620697022,-43.0119400024414,
44.8773651123047,-37.5938453674316,
92.4421539306641,-7.13094615936279,
92.9263153076172,21.9882431030273,
47.6346893310547,23.6618995666504,
0.719576358795166,-4.42196702957153,
-9.82168388366699,-34.1164627075195,
9.57186317443848,-37.0110626220703,
25.1919708251953,-19.8601760864258,
22.7398586273193,-11.4956178665161,
14.9171514511108,-16.9961757659912,
11.4680624008179,-12.6945762634277,
2.79766058921814,19.3694057464600,
-15.8839378356934,49.6689949035645,
-28.5449962615967,38.4561080932617,
-13.8095340728760,-3.49632382392883,
18.2104454040527,-20.4685611724854,
33.0953598022461,22.4663391113281,
13.8254642486572,89.3100585937500,
-17.9275798797607,112.700706481934,
-34.6202239990234,69.8488540649414,
-31.4464263916016,-2.92196130752563,
-26.7248668670654,-53.0581092834473,
-23.7289924621582,-57.7157249450684,
-11.9478769302368,-29.0616092681885,
10.8806962966919,9.81085681915283,
28.2913646697998,36.5179901123047,
24.8527584075928,34.1073570251465,
3.25348520278931,6.22706890106201,
-20.5552101135254,-25.1628780364990,
-33.8578605651856,-36.3500022888184,
-31.5890350341797,-25.3808956146240,
-15.1526985168457,-6.38239145278931,
8.21946239471436,9.15284347534180,
23.1772193908691,11.8924016952515,
16.6638069152832,-0.310096025466919,
-2.33294820785522,-19.8401355743408,
-14.3094396591187,-31.6761779785156,
-10.6216316223145,-15.0933780670166,
4.59490156173706,22.1799488067627,
14.8339624404907,48.5950088500977,
11.2145700454712,39.6708297729492,
-7.79173183441162,1.96038889884949,
-30.0639209747314,-35.3827018737793,
-38.5332260131836,-48.3971366882324,
-23.4418029785156,-33.6173667907715,
2.37422060966492,-1.54450213909149,
9.64330673217773,23.8980693817139,
-11.6303672790527,20.9983196258545,
-32.2382469177246,-8.40464687347412,
-20.5261459350586,-36.8333740234375,
14.3425045013428,-33.0239219665527,
28.4143981933594,-4.66371297836304,
0.761223316192627,14.3588361740112,
-39.2861671447754,8.77581596374512,
-52.6238899230957,0.285157799720764,
-36.8523674011231,15.3103256225586,
-22.2961826324463,42.0603027343750,
-27.5958118438721,49.1305122375488,
-35.9860038757324,31.6699409484863,
-28.2968692779541,11.3586578369141,
-6.63208580017090,2.60189509391785,
17.8316078186035,-1.89744532108307,
36.2534828186035,-12.2801151275635,
42.5798530578613,-18.9874801635742,
28.0596332550049,-6.87472963333130,
-0.286096602678299,18.7074508666992,
-16.1868515014648,37.4192619323731,
-4.85875844955444,39.9785079956055,
12.4281415939331,27.2237529754639,
9.04356193542481,6.99747276306152,
-7.78561115264893,-13.8120880126953,
-5.84823274612427,-19.5767860412598,
24.2642440795898,-7.66352653503418,
44.5469017028809,0.880168616771698,
29.0656414031982,-13.5385828018188,
-5.28746509552002,-34.3628654479981,
-20.9368114471436,-27.1312294006348,
-14.6074342727661,14.4485778808594,
-7.80333375930786,43.5101776123047,
-10.0077123641968,22.1667079925537,
-9.48211193084717,-22.4362144470215,
-1.44274747371674,-27.9580993652344,
3.43340921401978,17.5176734924316,
1.78193640708923,62.0692749023438,
2.78987288475037,64.8907623291016,
12.2562036514282,43.0580863952637,
13.4502620697021,31.6072044372559,
-4.73529052734375,29.9630832672119,
-31.8234272003174,11.6391181945801,
-48.2971267700195,-17.5484066009522,
-49.9259262084961,-20.3019866943359,
-42.4601936340332,12.1743822097778,
-24.3641414642334,38.8667602539063,
-2.11093759536743,34.1848487854004,
3.74652957916260,19.5626201629639,
-16.6563796997070,27.1885566711426,
-35.9183082580566,42.9010734558106,
-20.3754577636719,29.5638217926025,
20.7297668457031,-2.13292074203491,
39.0657272338867,-8.85434818267822,
7.19827461242676,20.0942916870117,
-46.4503288269043,36.9571571350098,
-72.9555130004883,11.4822635650635,
-59.6139144897461,-23.4884281158447,
-31.0919265747070,-14.0894737243652,
-7.72358036041260,23.4336547851563,
5.17226219177246,26.0712356567383,
6.21287202835083,-24.8967590332031,
-0.989154338836670,-75.7020568847656,
-1.32855403423309,-70.0114898681641,
21.6112785339355,-22.5290412902832,
49.8891181945801,18.2594146728516,
50.2872047424316,33.9554443359375,
11.5200614929199,45.5430374145508,
-37.6320457458496,55.6104698181152,
-64.4415283203125,40.7671928405762,
-62.1585121154785,-9.27324199676514,
-44.6496429443359,-56.3400688171387,
-23.5186500549316,-63.4782600402832,
0.718189477920532,-40.8646316528320,
24.6595325469971,-25.1148891448975,
38.9715232849121,-24.5495605468750,
43.8331794738770,-13.6020193099976,
40.4505386352539,22.2504920959473,
23.0100212097168,61.8734703063965,
-12.3052167892456,70.8560333251953,
-46.8741836547852,45.6522979736328,
-57.0691413879395,19.1443881988525,
-41.7431335449219,13.0130586624146,
-22.7699985504150,27.7998657226563,
-17.2532024383545,44.8838233947754,
-33.3778686523438,41.7260246276856,
-59.9724845886231,11.9998178482056,
-77.8616333007813,-26.3757476806641,
-66.6003341674805,-39.0177764892578,
-18.7782039642334,-14.4839382171631,
31.8927688598633,18.4096641540527,
34.6711502075195,25.3995780944824,
-12.7085113525391,6.10976314544678,
-46.6345329284668,-4.09353590011597,
-18.2396392822266,9.75980186462402,
36.5433082580566,19.1664581298828,
42.7875862121582,-6.90049743652344,
-2.70915794372559,-43.7475433349609,
-26.0593452453613,-50.3888778686523,
18.1002178192139,-24.3298721313477,
79.2885742187500,-3.35185456275940,
79.6181640625000,-7.07736682891846,
24.2722492218018,-19.5881977081299,
-13.5456037521362,-17.6920280456543,
-3.44648528099060,-9.26826286315918,
5.39658355712891,-6.61505031585693,
-20.9978275299072,-2.85474324226379,
-50.1591224670410,7.77683353424072,
-33.2482757568359,9.55548572540283,
14.1525001525879,-8.48293113708496,
40.8672180175781,-21.0730972290039,
36.3791236877441,4.03142023086548,
36.0592765808106,46.5881500244141,
50.7494812011719,49.4452400207520,
53.7972373962402,8.79588699340820,
30.7451915740967,-20.8953285217285,
11.2449855804443,1.17151272296906,
21.3508129119873,46.2551727294922,
34.6527748107910,58.3768119812012,
16.0223159790039,26.4593353271484,
-14.0097656250000,-14.8026437759399,
-15.3898639678955,-37.5568389892578,
8.15935897827148,-47.5201721191406,
18.2372970581055,-48.5640449523926,
3.49356794357300,-36.5666084289551,
-1.31156671047211,-21.5307064056397,
23.5313072204590,-19.0069160461426,
49.3706741333008,-16.4247283935547,
39.1632461547852,16.3874797821045,
7.76668691635132,71.5372238159180,
-7.01339578628540,97.0816726684570,
-6.97751855850220,69.7505722045898,
-17.8373165130615,29.7782363891602,
-37.3210029602051,23.3944606781006,
-33.6874961853027,35.3862075805664,
-5.81172704696655,16.6423168182373,
6.14079618453980,-36.8391265869141,
-18.5014343261719,-63.6366271972656,
-46.2681198120117,-32.5238914489746,
-36.5556488037109,17.4425468444824,
3.06137752532959,37.8073234558106,
29.5606079101563,27.6889247894287,
26.0690708160400,16.8841476440430,
21.8751335144043,9.50831127166748,
32.0575790405273,-2.51074337959290,
36.9496345520020,-9.03329849243164,
18.2999649047852,8.41402912139893,
-12.5687131881714,35.9190711975098,
-36.2720603942871,38.5872726440430,
-44.9684257507324,15.7722129821777,
-41.6117134094238,9.12109184265137,
-24.8449420928955,40.0549468994141,
-7.76127433776856,70.5588836669922,
-9.88647842407227,56.2483749389648,
-33.7182922363281,10.7803344726563,
-38.6245193481445,-17.2808952331543,
7.07381772994995,-14.5416946411133,
71.7785949707031,-3.75839996337891,
83.9356307983398,-1.95034217834473,
27.6970272064209,0.387300223112106,
-31.0900249481201,10.8894824981689,
-27.3470802307129,13.1059961318970,
20.1193618774414,-2.02062344551086,
41.1698722839356,-12.0484142303467,
10.1086788177490,2.45914649963379,
-35.4646186828613,20.8151760101318,
-49.9900131225586,11.5238780975342,
-38.7494468688965,-20.2164058685303,
-39.0186576843262,-32.7964668273926,
-59.8626937866211,-13.3548641204834,
-72.0549163818359,6.85889863967896,
-50.6545829772949,-1.04041361808777,
-8.68998432159424,-23.5122528076172,
16.3946475982666,-25.8483791351318,
4.80736446380615,-5.11068820953369,
-23.7786483764648,13.3473377227783,
-29.2503013610840,16.7951869964600,
5.37721014022827,20.9969253540039,
42.2680358886719,36.0468444824219,
35.0476264953613,42.4130401611328,
-12.3445816040039,18.0231876373291,
-47.8318786621094,-21.6021881103516,
-32.5897521972656,-42.0221672058106,
12.8908615112305,-33.4176139831543,
36.5162467956543,-22.5200691223145,
20.8879375457764,-33.1360702514648,
0.828069329261780,-55.7442131042481,
7.39007520675659,-53.1217308044434,
22.0418682098389,-11.5399284362793,
17.7539558410645,37.3976402282715,
-3.06371784210205,54.2913932800293,
-10.9666442871094,33.8499603271484,
3.79618406295776,4.38874340057373,
22.7788658142090,-0.168696522712708,
26.9300689697266,18.4328575134277,
22.0983505249023,25.7470798492432,
17.6610145568848,-0.623412847518921,
10.4552097320557,-34.5290985107422,
-0.389364600181580,-36.4733276367188,
-0.389422059059143,-8.41091060638428,
19.7299499511719,4.29502916336060,
36.3206481933594,-20.9123516082764,
17.7348175048828,-46.2320785522461,
-20.7351913452148,-21.8719902038574,
-36.6869087219238,35.7524299621582,
-18.9723434448242,52.6473350524902,
-4.20717620849609,6.63262033462524,
-20.9569454193115,-44.9871597290039,
-48.9434852600098,-44.7340164184570,
-48.0463066101074,-18.0068874359131,
-17.9836997985840,-25.4503860473633,
8.95000839233398,-63.6091270446777,
25.2863903045654,-70.1925277709961,
47.5144577026367,-21.8407955169678,
62.4908981323242,33.7033576965332,
36.3617935180664,45.8629112243652,
-19.8650627136230,28.1215000152588,
-42.9211120605469,17.5584259033203,
-1.63500988483429,16.1355915069580,
47.7050819396973,-1.75119829177856,
35.9254150390625,-29.5810413360596,
-15.0058393478394,-42.0383987426758,
-24.9974002838135,-43.3462638854981,
20.4676742553711,-54.9408378601074,
48.2215881347656,-65.9181594848633,
10.5539379119873,-49.6414031982422,
-41.1423606872559,-16.7276306152344,
-36.8021011352539,-11.1355361938477,
-1.64526724815369,-42.9263229370117,
-2.82864189147949,-60.0189094543457,
-41.2579231262207,-29.1957969665527,
-50.8522567749023,17.9181938171387,
-0.884625911712647,24.5103969573975,
47.2686767578125,4.92385578155518,
36.8102302551270,15.4952268600464,
-9.20580673217773,52.1077308654785,
-23.1793022155762,55.3059806823731,
10.7426319122314,4.42354249954224,
48.8973350524902,-42.0214805603027,
57.0102577209473,-31.2364063262939,
42.6553153991699,17.2595233917236,
13.0332288742065,44.8507843017578,
-29.4742317199707,33.4914245605469,
-62.1875991821289,1.14007580280304,
-53.9308815002441,-33.1822814941406,
-8.83262443542481,-66.2444534301758,
26.1803379058838,-75.7539520263672,
17.9717292785645,-37.5379791259766,
-15.6526317596436,22.5196876525879,
-35.3268394470215,39.4509735107422,
-33.6898078918457,0.706225156784058,
-34.8189239501953,-34.5470962524414,
-39.5421066284180,-23.9116115570068,
-30.1843509674072,4.17717361450195,
-17.5067558288574,5.56285762786865,
-27.9963912963867,-10.6213569641113,
-53.2295913696289,-7.34329986572266,
-56.1572380065918,7.34806680679321,
-24.4668483734131,-8.33834171295166,
9.38949775695801,-52.9505691528320,
21.3748416900635,-60.4683189392090,
31.4182052612305,-8.33587646484375,
54.3000717163086,40.5517158508301,
68.3085174560547,27.3820705413818,
43.2163658142090,-24.5669593811035,
3.12869811058044,-45.6376495361328,
2.63679742813110,-30.6564884185791,
36.9042816162109,-25.0607547760010,
45.7640419006348,-38.4540176391602,
8.94447040557861,-27.4163532257080,
-25.4469032287598,24.0369625091553,
-11.1832342147827,65.4049682617188,
24.0727787017822,50.9043350219727,
28.3289661407471,18.2575263977051,
2.29613232612610,30.2506694793701,
-16.4557743072510,77.4657135009766,
-17.9255065917969,87.4246063232422,
-29.3100070953369,30.0975074768066,
-51.6305427551270,-38.6505928039551,
-44.5123977661133,-62.7221679687500,
6.97945404052734,-45.4694595336914,
55.0374679565430,-25.6552715301514,
45.8836631774902,-19.6624622344971,
-0.562799215316773,-11.4520978927612,
-22.6841449737549,4.70209693908691,
1.48606407642365,13.7168245315552,
35.2631301879883,10.9078931808472,
38.6256294250488,10.3933992385864,
11.6135139465332,23.7218227386475,
-14.9775190353394,37.4111442565918,
-20.3676776885986,38.5547103881836,
-9.99380111694336,29.0536079406738,
2.06566882133484,10.0099773406982,
1.49273788928986,-17.5098114013672,
-15.0579347610474,-41.0689582824707,
-30.7864398956299,-45.1754722595215,
-25.8067798614502,-21.2286968231201,
-2.24053931236267,15.9298877716064,
8.78883552551270,39.0510902404785,
-7.05752134323120,44.7319221496582,
-22.4732627868652,42.0918159484863,
-5.64369535446167,37.1938133239746,
33.5669250488281,28.8365192413330,
49.6086807250977,23.2325706481934,
22.6969833374023,31.8436527252197,
-14.3214006423950,48.8264656066895,
-14.2518959045410,46.2891540527344,
22.9144439697266,14.1479187011719,
55.0207901000977,-22.0538196563721,
48.6079139709473,-25.5173110961914,
16.5897140502930,7.93328189849854,
-8.86637783050537,37.8914833068848,
-12.1432037353516,26.8755130767822,
-5.52287435531616,-17.5531558990479,
-7.58475112915039,-48.9234733581543,
-21.0215091705322,-40.3412055969238,
-25.0789146423340,-6.36039495468140,
-4.72788047790527,17.0147972106934,
24.2867202758789,5.75860214233398,
29.2519760131836,-23.1515903472900,
1.69054388999939,-33.4951858520508,
-25.9393081665039,-2.15049433708191,
-20.4982795715332,51.0785293579102,
8.06002712249756,80.9691162109375,
10.7480077743530,58.6652717590332,
-32.1821975708008,9.31013107299805,
-72.1590576171875,-16.0559501647949,
-57.0408706665039,-0.176687955856323,
-5.07188034057617,17.9280815124512,
22.3509197235107,-4.53319072723389,
-1.46831357479095,-46.4761238098145,
-33.2249565124512,-50.5988540649414,
-26.8226871490479,-6.03899192810059,
6.45144462585449,38.7861938476563,
23.0564746856689,36.0747833251953,
14.3347845077515,7.92249107360840,
7.13282728195190,6.46039867401123,
8.60648250579834,42.1007766723633,
0.631256818771362,70.1253967285156,
-16.5718574523926,59.9651107788086,
-9.15164375305176,27.9738426208496,
31.2916164398193,5.54693078994751,
58.0419082641602,1.75749063491821,
30.8808040618897,6.79557180404663,
-24.4161148071289,15.7535943984985,
-45.3108634948731,18.9736347198486,
-21.2855930328369,1.32272875308990,
1.44431757926941,-31.3702259063721,
-6.35321903228760,-52.8208351135254,
-14.9619369506836,-49.4876518249512,
4.55787515640259,-40.3241882324219,
30.1987857818604,-50.8375091552734,
28.8803272247314,-68.6890258789063,
15.0902433395386,-57.4165687561035,
18.6357192993164,-16.9694442749023,
29.5601882934570,12.9966106414795,
13.0903587341309,12.0987644195557,
-22.9671058654785,7.86500072479248,
-27.6449470520020,17.2378711700439,
17.0819911956787,25.3288688659668,
54.6928367614746,13.8698749542236,
34.7395324707031,2.77040052413940,
-14.1924610137939,14.3528108596802,
-25.8575439453125,33.2654266357422,
8.79946517944336,27.6462955474854,
37.6842269897461,-0.218456983566284,
32.3523521423340,-12.6272830963135,
21.7971458435059,0.300528407096863,
27.2229881286621,2.59613204002380,
31.6078624725342,-17.5246505737305,
12.5904655456543,-24.4370975494385,
-13.1935396194458,12.3778190612793,
-18.5943145751953,54.9877014160156,
-16.7431545257568,58.2841033935547,
-37.8057250976563,28.0065574645996,
-74.6382293701172,3.67202615737915,
-79.9952087402344,-6.37832069396973,
-32.9694519042969,-26.6251525878906,
26.9715213775635,-51.8110046386719,
56.2489547729492,-36.0513687133789,
52.0141792297363,28.9770393371582,
25.7513389587402,79.7071151733398,
-14.9306907653809,59.1669807434082,
-58.1664352416992,-0.789803028106690,
-81.0293884277344,-27.6987342834473,
-68.9219055175781,-16.7213039398193,
-37.6636886596680,-22.9048080444336,
-12.3107509613037,-66.7657470703125,
6.40057945251465,-92.1058959960938,
33.5719833374023,-54.1214332580566,
60.5730552673340,15.2924947738647,
63.4079475402832,50.3645896911621,
48.3148422241211,36.5597839355469,
44.6361732482910,20.6753864288330,
53.2301864624023,30.2173023223877,
34.5366821289063,43.8148002624512,
-17.1528854370117,37.2006225585938,
-57.3400077819824,17.9838371276855,
-44.1170272827148,5.85487318038940,
-2.16298627853394,-6.35830211639404,
8.02789306640625,-22.5888462066650,
-19.6295127868652,-38.4594078063965,
-36.0298843383789,-46.4772033691406,
-11.9039869308472,-48.9434776306152,
13.9875631332397,-49.5532112121582,
9.74713802337647,-40.0559883117676,
-5.16381454467773,-15.8372364044189,
2.22897100448608,12.7313480377197,
17.2413196563721,20.0704154968262,
1.49217176437378,8.69526672363281,
-29.1932334899902,-1.76155567169189,
-23.9343414306641,-4.52766799926758,
29.2582073211670,-7.14909410476685,
68.7577743530273,-2.11597800254822,
47.4241905212402,27.5615119934082,
-5.19476652145386,64.6224136352539,
-23.1207141876221,68.6316375732422,
-0.260331481695175,31.4418678283691,
7.13270521163940,-4.09049320220947,
-24.6713905334473,-0.686589241027832,
-57.6891136169434,23.0866088867188,
-55.1633949279785,15.5981788635254,
-25.4929389953613,-26.8951110839844,
0.876776278018951,-62.5944557189941,
13.9672079086304,-68.0360565185547,
25.5463714599609,-62.9353981018066,
31.7383937835693,-58.0422897338867,
20.9146709442139,-31.5690078735352,
0.0608549416065216,12.7403640747070,
-12.5237522125244,32.6356315612793,
-19.4843025207520,2.23178148269653,
-34.4914588928223,-32.3141670227051,
-45.0357589721680,-12.3704462051392,
-20.6824893951416,41.5247306823731,
25.5835342407227,50.9718284606934,
38.5944747924805,-4.11014938354492,
-1.08362674713135,-54.0061607360840,
-42.4216766357422,-36.0073394775391,
-24.7942657470703,15.9668369293213,
37.2748222351074,29.4884433746338,
73.1015548706055,4.83303928375244,
50.1865997314453,3.93575906753540,
5.30128955841064,47.7889556884766,
-14.9152307510376,83.8905105590820,
-11.5599088668823,57.6567115783691,
-13.4874181747437,-6.63132619857788,
-23.7276210784912,-48.0404701232910,
-25.7094306945801,-40.2908248901367,
-12.8853254318237,-12.0106582641602,
4.87560939788818,5.04032611846924,
16.6675662994385,6.75900411605835,
23.0533771514893,2.26166486740112,
27.8431968688965,-6.51039743423462,
36.2218360900879,-17.8304691314697,
46.9226913452148,-13.4455881118774,
48.8123130798340,9.99948215484619,
30.6441268920898,34.3022651672363,
-3.49228429794312,37.5160026550293,
-28.2178249359131,16.4434318542480,
-17.6012058258057,-9.35420608520508,
15.4452028274536,-25.6429805755615,
38.6033782958984,-37.4312744140625,
37.0789222717285,-53.6225700378418,
25.5605545043945,-58.7376136779785,
20.4012966156006,-35.1236534118652,
16.5525398254395,8.33245658874512,
5.80274534225464,37.7119789123535,
-4.88457059860230,24.3935241699219,
-2.27677011489868,-21.4162788391113,
9.90719318389893,-57.3590011596680,
16.5220947265625,-52.1993446350098,
10.6052703857422,-12.1342649459839,
4.55041265487671,24.8551902770996,
6.17647171020508,31.8287277221680,
14.1866731643677,10.8763751983643,
21.5873680114746,-11.1580514907837,
26.8166790008545,-12.8230171203613,
23.3428573608398,-0.132246613502502,
-0.348793745040894,3.69073891639709,
-42.1018562316895,-7.14348793029785,
-73.0830230712891,-16.6198844909668,
-70.5997772216797,-10.7893342971802,
-40.9144477844238,-3.04163074493408,
-12.5168418884277,-9.09799194335938,
0.510133981704712,-24.7415275573730,
10.8282756805420,-29.1230049133301,
30.5231914520264,-18.0765266418457,
46.8106765747070,-16.1508369445801,
40.6545104980469,-36.7262878417969,
21.9597244262695,-55.3046646118164,
13.7819433212280,-49.8619537353516,
19.1330642700195,-30.8846836090088,
25.0766696929932,-26.0574398040772,
27.6246051788330,-32.0242195129395,
33.9709205627441,-21.9642410278320,
40.2135963439941,5.95802164077759,
30.1266956329346,18.5006275177002,
4.30185985565186,-1.61071681976318,
-4.02033615112305,-27.7635345458984,
19.9917831420898,-29.6674194335938,
43.4079208374023,-12.6159114837646,
24.4249973297119,-6.97219467163086,
-12.4492568969727,-15.0567770004272,
-10.0987796783447,-12.3829860687256,
36.1460151672363,9.21539306640625,
61.8293228149414,25.0369243621826,
22.4420948028564,19.0514411926270,
-33.0329399108887,3.57640910148621,
-38.0016021728516,-4.50117826461792,
-1.22501957416534,2.12536454200745,
3.65506434440613,16.7922534942627,
-44.3813056945801,28.0153026580811,
-78.5299758911133,20.2593460083008,
-45.1353874206543,-11.0275411605835,
19.9317321777344,-40.6813240051270,
44.0265083312988,-32.9127960205078,
24.0281238555908,13.7507152557373,
15.3199739456177,49.8677253723145,
41.4250831604004,34.5757980346680,
61.1770782470703,-3.36006069183350,
38.7215881347656,-7.47924995422363,
-9.52417755126953,21.4168376922607,
-44.1143798828125,29.0955162048340,
-57.6768722534180,-6.94050407409668,
-67.7417068481445,-41.4585113525391,
-71.8571319580078,-31.2820415496826,
-54.2610359191895,5.20492839813232,
-22.0079021453857,22.8988113403320,
-1.58229327201843,16.3132266998291,
1.84428620338440,18.9102878570557,
9.26719856262207,33.9497718811035,
23.2303867340088,32.8718986511231,
27.5031261444092,5.59599399566650,
10.4846143722534,-14.3418445587158,
-12.8167448043823,-4.59782743453980,
-23.4605197906494,10.7447032928467,
-26.1221370697022,0.346028864383698,
-33.2350120544434,-21.3656406402588,
-32.7458801269531,-25.1684703826904,
-3.76593375205994,-13.3256540298462,
37.6294059753418,-12.2363328933716,
57.0986824035645,-22.0164489746094,
46.2085380554199,-15.8642807006836,
27.4125499725342,16.9863548278809,
13.8667840957642,48.7907066345215,
-2.51262855529785,51.2062988281250,
-28.9469413757324,39.4931869506836,
-44.5810699462891,41.6184654235840,
-34.9111747741699,56.4163475036621,
-18.8875408172607,59.9431076049805,
-19.4639492034912,45.8914718627930,
-25.0507545471191,26.1674365997314,
-3.04429316520691,12.6455173492432,
41.1407127380371,2.59201121330261,
56.6110229492188,-5.92638683319092,
18.7892742156982,-10.8203420639038,
-34.5624923706055,-13.1547870635986,
-48.7970733642578,-19.5911369323730,
-20.9991607666016,-23.2354640960693,
1.91185402870178,-8.37633705139160,
-13.0848884582520,25.6438064575195,
-46.7975349426270,47.4662208557129,
-60.6137924194336,29.3752403259277,
-41.3196067810059,-8.51119327545166,
-7.35450172424316,-24.2499389648438,
15.8712072372437,2.59044647216797,
19.0200710296631,43.2331771850586,
0.979137957096100,61.0345687866211,
-28.9270324707031,47.9786758422852,
-53.0449523925781,23.2464866638184,
-58.8155136108398,3.47023701667786,
-52.6910934448242,-9.01958370208740,
-48.5661239624023,-22.5495433807373,
-48.8203735351563,-38.4102668762207,
-40.6648254394531,-52.5303535461426,
-16.2084732055664,-60.2901115417481,
14.0223951339722,-51.2084617614746,
29.1780090332031,-23.8556632995605,
20.6838264465332,11.9037876129150,
0.348346590995789,40.8974380493164,
-19.9481544494629,51.5171546936035,
-26.2000579833984,36.8785476684570,
-14.3121376037598,-2.79850244522095,
10.9288940429688,-47.9244155883789,
28.2323360443115,-63.8928070068359,
21.0968608856201,-31.5126228332520,
-2.79257082939148,25.5354690551758,
-14.0932579040527,51.2610244750977,
2.05576086044312,21.5692138671875,
34.4519309997559,-20.5511703491211,
52.3353080749512,-15.6935348510742,
44.3031349182129,34.5908851623535,
14.8899288177490,68.4781723022461,
-18.9731082916260,44.2010650634766,
-47.0645599365234,-12.2082958221436,
-55.2801055908203,-43.1122131347656,
-43.9382514953613,-34.7804069519043,
-33.0715904235840,-17.7227401733398,
-36.6770248413086,-14.2967052459717,
-48.9233703613281,-10.4074916839600,
-48.4887390136719,2.60952520370483,
-36.3669967651367,1.85289049148560,
-27.3999958038330,-24.1409339904785,
-21.4176311492920,-51.4941177368164,
-0.585846185684204,-44.8186721801758,
39.2381706237793,-14.5495910644531,
65.0164566040039,-3.31001591682434,
51.7278099060059,-18.0410003662109,
25.5787963867188,-27.6001815795898,
35.6271286010742,-13.7115545272827,
72.3342056274414,0.836102128028870,
77.3656463623047,-8.55026245117188,
26.7056045532227,-26.3169059753418,
-35.9748077392578,-20.0588264465332,
-59.2929573059082,-0.104378342628479,
-52.4154548645020,-1.82804656028748,
-51.8502197265625,-29.1403045654297,
-55.1419906616211,-50.9629287719727,
-31.1117172241211,-46.5234375000000,
18.3843784332275,-26.9801025390625,
45.7408256530762,-5.01716184616089,
37.3169059753418,21.0435543060303,
32.2867813110352,40.7084350585938,
53.1736831665039,34.5735664367676,
65.4595336914063,5.31731891632080,
34.9034271240234,-12.0468063354492,
-4.54027652740479,9.60884380340576,
0.788794577121735,39.6415290832520,
41.2034530639648,29.1012935638428,
50.7428512573242,-14.9940338134766,
12.6405591964722,-43.1986274719238,
-17.6879673004150,-29.2143669128418,
3.97666501998901,3.20126175880432,
32.0112724304199,25.9853935241699,
10.4681358337402,30.5157985687256,
-41.4413490295410,17.1980972290039,
-49.2062110900879,-9.22116947174072,
0.879863262176514,-28.6577529907227,
40.5360908508301,-10.8099784851074,
23.8985843658447,35.3092155456543,
-16.5797863006592,48.7063293457031,
-23.3438816070557,-7.54086637496948,
1.49070250988007,-81.5291366577148,
14.5802755355835,-86.6487274169922,
-1.13271141052246,-16.3085498809814,
-15.2975959777832,47.2064704895020,
-6.42094087600708,43.5536117553711,
1.62779438495636,10.3650598526001,
-18.4899253845215,7.89401197433472,
-53.2427864074707,34.6731109619141,
-68.3500366210938,39.7621421813965,
-47.4576416015625,9.60047435760498,
-2.31239080429077,-11.2025165557861,
38.1778640747070,4.10758638381958,
46.8282318115234,24.5496330261230,
24.6430168151855,12.5695896148682,
-2.68565750122070,-19.5645217895508,
-13.3356027603149,-36.4997749328613,
-6.24892711639404,-34.5649032592773,
0.0532192364335060,-42.6340560913086,
-1.11188650131226,-62.5691795349121,
8.21732234954834,-66.3894271850586,
33.9671897888184,-47.4345817565918,
48.8003730773926,-32.9167175292969,
30.2625694274902,-43.9851417541504,
0.129999458789825,-60.6687164306641,
-5.62648153305054,-46.9563903808594,
7.16081237792969,-10.8211469650269,
0.289384722709656,10.4607696533203,
-30.3211917877197,1.97420799732208,
-38.9303283691406,-8.88472747802734,
1.76149368286133,3.26417970657349,
52.6193084716797,31.2439422607422,
54.7946662902832,49.8641357421875,
9.38755226135254,45.3524360656738,
-24.9762096405029,20.1606025695801,
-13.7857637405396,-16.9394321441650,
15.4370660781860,-53.0017814636231,
23.2705669403076,-68.6767272949219,
7.94768762588501,-54.9258270263672,
-4.57351779937744,-24.4650688171387,
-5.57211112976074,-9.25860595703125,
-3.03958916664124,-18.4875831604004,
2.95480060577393,-36.6510887145996,
17.5206851959229,-44.0130195617676,
28.2551269531250,-39.7980690002441,
13.2613363265991,-29.8811511993408,
-25.2723693847656,-19.2867374420166,
-52.4071578979492,-13.2836542129517,
-36.5386314392090,-11.0929698944092,
4.55016756057739,-3.87232542037964,
23.8944149017334,16.2293872833252,
5.61026573181152,42.0652236938477,
-30.2937412261963,43.2267417907715,
-53.1755065917969,8.33272933959961,
-49.2570037841797,-35.1222000122070,
-23.3591823577881,-46.3085517883301,
8.16886138916016,-20.3923835754395,
29.6471405029297,4.64866304397583,
32.9742965698242,7.71449232101440,
25.8784465789795,0.903267085552216,
25.3911495208740,0.0806511640548706,
29.5994167327881,-4.22351837158203,
16.6110477447510,-22.8067493438721,
-15.5656118392944,-39.9173202514648,
-35.6797790527344,-29.1694717407227,
-12.5364913940430,4.62649917602539,
29.5560092926025,28.1086082458496,
46.2491035461426,28.9368724822998,
27.9321651458740,27.0781040191650,
11.6780757904053,37.9344406127930,
24.6098918914795,42.9531364440918,
43.7141914367676,24.9172325134277,
36.7528839111328,3.10928845405579,
14.2937641143799,4.53357505798340,
9.36308956146240,21.7363033294678,
26.2505607604980,24.4951343536377,
32.7202453613281,3.78086376190186,
10.3076343536377,-12.7473983764648,
-21.5643272399902,-6.30274868011475,
-38.5970535278320,6.94161558151245,
-42.3605499267578,5.58166551589966,
-50.1826820373535,-5.62981081008911,
-59.3786735534668,-10.7195177078247,
-54.0818023681641,-16.0834407806397,
-28.1774482727051,-39.1070861816406,
9.76571846008301,-65.7469940185547,
40.2878150939941,-57.3768997192383,
51.0944175720215,-6.06533765792847,
38.4622230529785,41.9459762573242,
9.89087295532227,39.3311691284180,
-20.5920333862305,-5.79913711547852,
-29.7553558349609,-36.1627922058106,
-12.4386978149414,-18.2416667938232,
16.7902851104736,20.1407146453857,
34.7650947570801,30.4144363403320,
25.3874359130859,9.50394821166992,
-9.57015037536621,-10.7938070297241,
-43.0014266967773,-3.67543697357178,
-39.0091667175293,22.5602741241455,
5.31334209442139,34.4600219726563,
48.5766677856445,15.1632385253906,
44.2157630920410,-20.9150524139404,
-2.28137207031250,-42.3943367004395,
-27.4356613159180,-32.1860847473145,
9.97080039978027,-5.06701660156250,
70.3516387939453,11.7407608032227,
76.9999542236328,8.03084659576416,
12.6744003295898,3.74225640296936,
-53.7336235046387,16.3487758636475,
-57.4215812683106,24.3073005676270,
-12.6066331863403,-6.85084009170532,
18.4538021087647,-64.5847015380859,
12.0333080291748,-87.9203796386719,
2.28915500640869,-43.1248168945313,
20.2045459747314,30.5936298370361,
45.5564651489258,65.4214019775391,
41.9232788085938,44.4302330017090,
12.5309638977051,15.5209159851074,
-14.6320428848267,18.8100051879883,
-25.8347129821777,36.6571998596191,
-32.3029212951660,33.5072937011719,
-34.1658859252930,2.87668895721436,
-19.2754116058350,-23.3508987426758,
9.91881179809570,-20.9666347503662,
21.8730792999268,5.01617813110352,
5.39028835296631,31.5448169708252,
-18.4125862121582,34.1944274902344,
-22.7773666381836,4.96331071853638,
-9.91911506652832,-34.7320213317871,
-6.29602718353272,-44.3439369201660,
-8.83185291290283,-9.81022167205811,
7.48494338989258,34.2937355041504,
39.7300796508789,42.1620254516602,
53.9822998046875,5.13350915908814,
31.7883033752441,-40.9826202392578,
2.01764678955078,-59.2303390502930,
3.91671395301819,-49.9975547790527,
36.4711608886719,-33.2750930786133,
61.6017532348633,-15.2412776947021,
61.3174667358398,0.548370480537415,
45.0355453491211,6.82483959197998,
23.5489711761475,-2.48591279983521,
-7.25337886810303,-18.7438507080078,
-36.2911224365234,-29.2699241638184,
-32.6279449462891,-35.4683227539063,
8.40159606933594,-44.0301437377930,
41.3519859313965,-48.5094261169434,
21.5736846923828,-40.4320297241211,
-30.0806941986084,-27.0846004486084,
-47.1177024841309,-19.9084930419922,
-6.08628749847412,-18.5081844329834,
38.3891410827637,-8.08831977844238,
30.4111766815186,16.5662708282471,
-16.7707366943359,35.5884475708008,
-45.8928680419922,38.3172187805176,
-35.3773345947266,36.1463737487793,
-21.2741260528564,36.3780937194824,
-26.7459297180176,25.1462993621826,
-33.9105148315430,-5.24766635894775,
-17.7048206329346,-33.2415733337402,
7.19654226303101,-35.5731239318848,
8.50350189208984,-20.1190567016602,
-12.5830669403076,-15.7364425659180,
-25.3509941101074,-24.3745956420898,
-14.3292274475098,-14.9754390716553,
0.514220714569092,18.7420196533203,
-6.94421768188477,39.6422615051270,
-28.4791164398193,18.6676921844482,
-33.3996620178223,-16.5106105804443,
-11.1423168182373,-13.6927347183228,
21.9849338531494,29.7060031890869,
41.6366310119629,55.6240463256836,
36.4874191284180,31.2078876495361,
13.6481208801270,-11.0503225326538,
-11.9237375259399,-11.3857707977295,
-26.6042346954346,33.7458000183106,
-25.1770458221436,67.4156494140625,
-9.95549774169922,50.7280731201172,
6.01559782028198,9.78334236145020,
5.63596057891846,-6.37566518783569,
-15.9882469177246,5.73080348968506,
-37.1436347961426,9.79423046112061,
-31.4394454956055,-17.8175563812256,
-0.477912873029709,-50.7866935729981,
23.8434963226318,-53.5594367980957,
18.0425796508789,-25.4033641815186,
0.151073932647705,13.3245334625244,
8.50581359863281,46.7709770202637,
36.7189559936523,64.4672927856445,
44.4551811218262,50.2010269165039,
16.0611972808838,-0.519849300384522,
-6.15652465820313,-49.5639762878418,
7.52723550796509,-46.4392089843750,
25.5948009490967,1.89837074279785,
5.69241476058960,31.4772472381592,
-35.4770393371582,9.44884204864502,
-37.7015113830566,-27.2906303405762,
5.34035015106201,-21.6321964263916,
29.7348308563232,18.7332725524902,
-7.79625606536865,36.1412467956543,
-53.3804092407227,8.89028263092041,
-35.3624000549316,-21.6009826660156,
30.2955894470215,-20.6414394378662,
64.4086685180664,-4.74337720870972,
39.6169738769531,-1.35520637035370,
14.9673604965210,-12.5718364715576,
32.2043876647949,-23.9501438140869,
52.8399620056152,-28.1661891937256,
27.3423213958740,-22.2295532226563,
-22.8188877105713,1.43298995494843,
-37.0916519165039,33.6299934387207,
-17.6452770233154,47.4856681823731,
-22.9733409881592,24.5546894073486,
-68.6812744140625,-11.3271570205688,
-90.6748962402344,-25.2522869110107,
-42.7756767272949,-22.7277336120605,
26.0753631591797,-35.3232841491699,
38.1446189880371,-60.8486671447754,
-5.42176723480225,-58.4236984252930,
-38.7850875854492,-18.3322544097900,
-30.2401409149170,16.7018966674805,
-14.8854198455811,11.6358528137207,
-21.5009117126465,-12.9087810516357,
-27.1272583007813,-20.1500320434570,
1.70301163196564,-7.77182722091675,
40.8479881286621,-5.58679676055908,
43.0957527160645,-22.7145919799805,
15.7374000549316,-40.4654388427734,
8.21331977844238,-39.3204231262207,
32.3885498046875,-20.8843517303467,
48.1356391906738,3.11672139167786,
23.7652130126953,28.9113292694092,
-17.5027046203613,41.1475143432617,
-41.1924934387207,26.7853832244873,
-40.7354698181152,3.94552969932556,
-38.4519042968750,2.18458271026611,
-40.0817718505859,15.8507308959961,
-33.1750946044922,4.22953891754150,
-23.9796581268311,-38.5207557678223,
-30.2589702606201,-66.6239395141602,
-40.2944107055664,-46.0223007202148,
-29.0185146331787,-10.1866989135742,
-0.364120483398438,-14.9586114883423,
11.4103116989136,-48.3068504333496,
-3.16346788406372,-44.0872840881348,
-15.6901378631592,16.6717624664307,
-2.92537927627563,69.2133255004883,
8.62941741943359,58.9997711181641,
-12.2660551071167,15.0463743209839,
-52.1148033142090,-3.53849005699158,
-66.1078262329102,5.98088884353638,
-48.2729110717773,-1.16239202022553,
-37.3072891235352,-31.9582672119141,
-46.7530822753906,-43.7487487792969,
-43.7056922912598,-15.7906188964844,
-5.23197555541992,16.1687240600586,
38.3142852783203,12.6477851867676,
42.3049201965332,-12.3399772644043,
13.0360298156738,-19.9749641418457,
-4.26755189895630,-3.32894539833069,
10.2542734146118,5.88873481750488,
33.7328948974609,-0.821642458438873,
42.6125602722168,-0.218752086162567,
38.1405525207520,19.4480075836182,
29.9022712707520,35.3822402954102,
13.6164999008179,25.7839298248291,
-6.10197210311890,-1.96948027610779,
-3.58373069763184,-16.7101917266846,
37.8246498107910,-3.36101412773132,
81.0752334594727,24.2856426239014,
73.8308944702148,41.5008392333984,
7.71494245529175,36.7440948486328,
-61.9825820922852,19.3376865386963,
-78.5676574707031,4.30507040023804,
-43.5674362182617,4.69626569747925,
-6.50472164154053,22.1277198791504,
-6.20251417160034,39.2556953430176,
-28.9255237579346,42.6298637390137,
-42.4339599609375,34.9616584777832,
-34.3760833740234,22.5708103179932,
-18.7274761199951,7.67981195449829,
-16.0518608093262,-4.71949672698975,
-26.7865295410156,-6.32434225082398,
-38.3420028686523,4.42464733123779,
-37.2752037048340,14.3171138763428,
-27.9496650695801,0.952993631362915,
-24.2497730255127,-28.5502738952637,
-31.1146430969238,-37.0746879577637,
-35.2475814819336,-7.42214632034302,
-31.1440925598145,25.1304931640625,
-23.7118053436279,10.8184814453125,
-24.4191036224365,-42.9871101379395,
-34.4085922241211,-70.4214172363281,
-35.4646110534668,-32.7574424743652,
-21.7120056152344,26.7318477630615,
-7.05841493606567,34.7546463012695,
-0.0380263924598694,-16.4672145843506,
7.06289720535278,-57.7254753112793,
24.4707164764404,-34.2152290344238,
34.6899566650391,28.1021862030029,
24.7193889617920,64.3175506591797,
7.67036628723145,47.9385528564453,
9.47350311279297,0.590498328208923,
23.7683448791504,-45.1473350524902,
18.1843757629395,-71.8024673461914,
-15.2556724548340,-65.4919586181641,
-33.4662704467773,-26.2738628387451,
-6.76422405242920,17.1451377868652,
32.0065956115723,23.5329494476318,
28.4333820343018,-5.36968708038330,
-11.7185850143433,-21.0157852172852,
-35.9546470642090,3.22366762161255,
-25.5183582305908,34.3174743652344,
-24.4379787445068,25.2939720153809,
-59.0633888244629,-10.5197706222534,
-89.5716552734375,-21.3070850372314,
-62.6943855285645,7.03842926025391,
3.77678728103638,34.9679718017578,
37.3244552612305,35.5294456481934,
7.37454843521118,29.4032039642334,
-40.9202880859375,40.8967628479004,
-56.8889007568359,47.8716964721680,
-41.4932594299316,13.3160114288330,
-28.5352859497070,-42.9142494201660,
-26.2909297943115,-64.4408264160156,
-17.2314071655273,-26.7248744964600,
-0.886649191379547,21.9737777709961,
7.20750617980957,27.1014556884766,
7.97682666778564,-4.66806840896606,
15.1306934356689,-22.2770996093750,
30.1852283477783,-0.107887744903564,
30.9195671081543,38.4994621276856,
0.428954601287842,53.6897392272949,
-40.8399238586426,28.2760601043701,
-51.4422988891602,-13.6131744384766,
-17.5458431243897,-38.8057746887207,
31.2117481231689,-38.6323661804199,
54.3388862609863,-26.2103557586670,
32.6312522888184,-23.0038719177246,
-19.7410678863525,-30.9801616668701,
-60.6371345520020,-32.3057708740234,
-64.0964584350586,-12.1103916168213,
-40.8509902954102,12.8642616271973,
-24.0312442779541,18.6475048065186,
-29.4138469696045,11.3675327301025,
-36.7051239013672,15.9932403564453,
-23.7382755279541,30.6902332305908,
3.21932601928711,25.1314964294434,
22.1865673065186,-16.2936115264893,
28.3922653198242,-54.5156860351563,
39.5032997131348,-36.5904273986816,
55.0071144104004,22.0397205352783,
41.4275779724121,51.1448402404785,
-9.20513820648193,19.7816772460938,
-55.7489242553711,-24.0661582946777,
-55.8482551574707,-16.9184818267822,
-16.2655143737793,29.1292037963867,
10.2394742965698,47.2753715515137,
-4.85752296447754,11.5238828659058,
-35.7954788208008,-29.5440216064453,
-51.7141609191895,-33.6884918212891,
-50.8877601623535,-18.4657154083252,
-42.9245033264160,-25.2967281341553,
-16.9980545043945,-51.7493515014648,
28.6522121429443,-52.8670845031738,
59.1889610290527,-12.9679355621338,
31.4722366333008,26.0516014099121,
-36.5184974670410,19.4795932769775,
-68.2102203369141,-22.4137420654297,
-20.2687873840332,-47.6068038940430,
51.9286613464356,-26.6270446777344,
64.8355484008789,17.8311252593994,
12.9865493774414,36.5893211364746,
-31.2160949707031,7.85192489624023,
-14.5719251632690,-38.3236732482910,
26.8439044952393,-58.0386276245117,
25.9377765655518,-40.2358055114746,
-18.2453479766846,-12.6933813095093,
-40.7468070983887,-5.60911989212036,
-9.59056377410889,-18.3914394378662,
33.8877410888672,-22.1664505004883,
32.8593406677246,-2.06724357604980,
-5.62690353393555,24.6530036926270,
-24.7066783905029,33.4732933044434,
1.59168338775635,26.0807247161865,
33.7239456176758,14.7450895309448,
18.6258239746094,4.67698383331299,
-25.1995639801025,-7.66752052307129,
-35.3498115539551,-23.8978939056397,
4.41165542602539,-33.7462387084961,
46.2147407531738,-30.6756896972656,
32.7820091247559,-22.8664321899414,
-20.7371921539307,-15.5865907669067,
-46.1836242675781,-0.605953454971314,
-15.6048431396484,25.6806697845459,
19.2676715850830,44.7211227416992,
4.01071548461914,30.8343944549561,
-39.6644477844238,-10.8735580444336,
-48.6609954833984,-38.3293418884277,
-8.01377487182617,-18.7265682220459,
24.5381603240967,24.1466197967529,
2.15969824790955,39.1871414184570,
-40.5397300720215,9.82987880706787,
-34.2009239196777,-22.8043708801270,
27.6274909973145,-18.7633342742920,
80.4863815307617,8.24895954132080,
73.0988388061523,16.1918048858643,
28.8754787445068,-0.623363375663757,
4.29856967926025,-4.58716821670532,
11.6962375640869,23.8277053833008,
13.9454965591431,58.8920440673828,
-15.9381999969482,61.4222488403320,
-60.2131423950195,31.9152927398682,
-81.1368179321289,3.18076729774475,
-61.2695999145508,-5.88344430923462,
-14.4423294067383,3.03383708000183,
26.3287868499756,19.5052375793457,
31.8412513732910,38.1075744628906,
4.37316942214966,46.2592964172363,
-24.9443817138672,32.2810478210449,
-19.8241882324219,7.27142858505249,
16.8323650360107,-0.588143944740295,
39.7483024597168,13.2919569015503,
16.2030010223389,20.2418212890625,
-27.6077213287354,-0.439264297485352,
-41.9049377441406,-30.7548065185547,
-10.3470792770386,-37.7393112182617,
31.5366878509522,-13.2493801116943,
44.4935760498047,16.2794857025147,
27.1855068206787,22.4197235107422,
4.49524974822998,7.56046056747437,
-7.15579700469971,-14.9894752502441,
-12.2143478393555,-33.6124763488770,
-6.71160125732422,-41.8980789184570,
14.5727424621582,-38.8340377807617,
39.6677474975586,-26.7382202148438,
43.9116592407227,-10.2375087738037,
18.3593959808350,11.4696350097656,
-13.1265687942505,34.2696723937988,
-22.9679107666016,38.2184257507324,
-11.8744211196899,9.17450046539307,
-1.38049697875977,-35.8973159790039,
0.415646344423294,-55.4875259399414,
1.21873486042023,-28.2784538269043,
3.01403379440308,17.9890880584717,
-4.53263759613037,36.2238388061523,
-19.1876335144043,15.7833595275879,
-17.2088966369629,-14.9943809509277,
10.5501852035522,-27.3441181182861,
34.9952583312988,-20.4027843475342,
22.9579086303711,-2.37846398353577,
-14.2752628326416,21.6842918395996,
-29.9605598449707,47.2933273315430,
-6.18220043182373,53.3570213317871,
19.4786357879639,32.0707855224609,
5.78962326049805,-2.02244400978088,
-35.3539848327637,-22.4255123138428,
-53.6797485351563,-18.6337547302246,
-27.9513359069824,-1.35931527614594,
13.0202903747559,11.5780124664307,
27.7057132720947,12.5051002502441,
7.84544563293457,-0.229715585708618,
-23.1893386840820,-25.7269935607910,
-37.8245353698731,-51.6184883117676,
-23.9742088317871,-59.0128593444824,
12.5264616012573,-46.8351936340332,
48.3996238708496,-26.7486820220947,
56.0024185180664,-4.13286876678467,
30.6283721923828,25.6186180114746,
-2.12182283401489,57.7931289672852,
-7.38402557373047,66.0594863891602,
14.3793907165527,32.7538719177246,
29.5177154541016,-12.0112161636353,
17.7869529724121,-22.6725463867188,
-6.74631977081299,13.1799802780151,
-19.0356521606445,53.4671478271484,
-15.6739740371704,51.6735458374023,
-11.3907995223999,14.6085290908813,
-13.4100027084351,-9.61779594421387,
-11.6328582763672,4.53905200958252,
0.103699445724487,33.4470787048340,
9.98170948028565,34.7713317871094,
7.78604030609131,0.614641666412354,
-4.57348442077637,-38.5232925415039,
-18.7944717407227,-42.4193267822266,
-29.8908519744873,-11.9273843765259,
-36.9158325195313,11.2577428817749,
-29.0683727264404,-6.39928865432739,
-5.54797220230103,-48.9342689514160,
22.7470207214355,-59.8829536437988,
40.0125160217285,-17.0495815277100,
42.5674705505371,39.0576744079590,
38.6297416687012,47.4531784057617,
29.8616771697998,0.0770401954650879,
8.18126296997070,-45.7633361816406,
-20.4260768890381,-44.2058639526367,
-32.5310134887695,-14.6860179901123,
-15.8879108428955,-2.19715523719788,
8.57468032836914,-13.0581245422363,
16.6739273071289,-13.4337759017944,
10.8964147567749,16.9048652648926,
6.28698253631592,55.7039489746094,
0.617741525173187,66.2753143310547,
-22.3622188568115,43.4866485595703,
-55.9014472961426,7.07795381546021,
-60.5046157836914,-22.0359477996826,
-21.5047950744629,-30.8115959167480,
26.4326438903809,-15.5217437744141,
35.2782325744629,8.72669029235840,
10.8633308410645,14.8677730560303,
-4.60055828094482,-11.4345560073853,
4.41567993164063,-41.9337081909180,
6.31452560424805,-40.0849037170410,
-14.5177936553955,-11.9799089431763,
-30.0708160400391,2.12073302268982,
-11.3981132507324,-18.7620124816895,
23.4517459869385,-48.8690948486328,
28.9201240539551,-50.1266708374023,
-4.46071910858154,-26.5776920318604,
-36.4275779724121,-11.5995645523071,
-32.9811820983887,-18.6599712371826,
0.173789262771606,-23.7556419372559,
34.3596420288086,-15.1311292648315,
50.7976646423340,-2.18111324310303,
52.8530769348145,1.11270868778229,
44.7509078979492,2.10937142372131,
37.0353088378906,13.2946395874023,
40.8334655761719,22.0527820587158,
51.6513519287109,11.9130191802979,
52.4310073852539,-4.35257673263550,
30.7261543273926,4.26229000091553,
-3.69423985481262,39.6074752807617,
-22.4036045074463,61.7807693481445,
-8.09877490997315,41.8314018249512,
26.2604694366455,7.18184852600098,
45.8613357543945,6.15263795852661,
27.8176746368408,38.9666557312012,
-17.6524791717529,55.9615402221680,
-51.5752220153809,24.7122421264648,
-38.5098571777344,-24.5059223175049,
9.75921821594238,-39.8940124511719,
44.3231620788574,-14.3316001892090,
32.1956748962402,15.0327224731445,
-10.0725975036621,21.4868736267090,
-32.3915519714356,18.9823513031006,
-17.9079380035400,25.3990230560303,
10.8130817413330,32.5104713439941,
29.0144367218018,23.5366363525391,
30.6610412597656,7.70392370223999,
29.0799274444580,11.4642314910889,
25.2433300018311,33.8171958923340,
10.3346481323242,50.6393775939941,
-9.03445720672607,40.7303276062012,
-17.8094520568848,15.0416898727417,
-10.1662445068359,-1.54013311862946,
4.90840911865234,-4.51429128646851,
16.8824920654297,-9.64130401611328,
20.6787967681885,-21.4246234893799,
11.8311929702759,-31.9054508209229,
-16.1077251434326,-33.3462333679199,
-49.6183090209961,-27.1161460876465,
-54.2004814147949,-19.6990642547607,
-11.2516908645630,-16.7398452758789,
51.5639305114746,-9.98204135894775,
82.9376373291016,11.0364780426025,
56.3583641052246,40.3657531738281,
0.193489551544189,55.6213264465332,
-43.6886024475098,35.0150032043457,
-58.3349037170410,-11.3830595016480,
-52.6147079467773,-44.9394035339356,
-34.3216781616211,-34.2612113952637,
-10.2270622253418,4.20948934555054,
7.15145587921143,34.5490608215332,
6.14899492263794,42.0756874084473,
-5.98817777633667,41.6807327270508,
-6.65503120422363,36.0230140686035,
9.74416732788086,7.98899555206299,
21.5261821746826,-40.3974876403809,
15.2095394134521,-69.6984176635742,
7.91581439971924,-43.0066223144531,
22.2823333740234,17.8806533813477,
44.2133903503418,54.1018447875977,
38.3640174865723,40.4442863464356,
5.25236129760742,8.93706989288330,
-14.6079711914063,1.15128898620605,
5.77735233306885,15.4654750823975,
40.4760665893555,26.5233078002930,
44.1693496704102,30.0334014892578,
10.8280315399170,39.7565460205078,
-24.4548397064209,50.7286071777344,
-30.4827251434326,46.4311523437500,
-11.7371902465820,27.0003166198730,
5.97016620635986,8.56509590148926,
7.66942453384399,3.90658998489380,
-7.87134742736816,5.34617137908936,
-32.9323196411133,2.97711586952209,
-52.1380844116211,1.38453948497772,
-51.8415756225586,-3.83898806571960,
-38.2408523559570,-27.0685825347900,
-25.8101158142090,-67.4479522705078,
-10.0357179641724,-82.6366195678711,
17.8264579772949,-46.7767219543457,
47.9497299194336,4.67299985885620,
53.7837028503418,14.1164045333862,
28.9932212829590,-15.1823549270630,
4.11340284347534,-25.2526016235352,
12.4093275070190,10.4433727264404,
39.2691574096680,38.5355453491211,
46.3756790161133,8.66067504882813,
32.1216278076172,-48.0433959960938,
24.4325294494629,-54.4274711608887,
27.1010150909424,-2.33800053596497,
12.8711690902710,40.5815353393555,
-18.2695083618164,32.1091690063477,
-25.8665180206299,7.66422653198242,
13.1631145477295,10.8822956085205,
53.2816848754883,27.0914154052734,
41.2648124694824,19.7688159942627,
-6.75039482116699,-1.90514862537384,
-22.2996063232422,-1.09926569461823,
10.2099819183350,22.0485324859619,
33.9965095520020,30.7201766967773,
9.41732978820801,11.5327548980713,
-24.1060791015625,-3.24601674079895,
-19.6706218719482,8.84199047088623,
3.31086254119873,20.9427509307861,
-10.4000701904297,0.367183446884155,
-52.1772308349609,-35.2851104736328,
-55.4603958129883,-44.0363273620606,
3.08009147644043,-21.2238082885742,
57.4747467041016,2.44191145896912,
43.5303192138672,3.67547607421875,
-8.79842948913574,-7.94591331481934,
-20.9028892517090,-10.4567794799805,
18.8019599914551,6.41225242614746,
42.4223442077637,28.1210002899170,
7.40024948120117,37.2257385253906,
-36.3390235900879,25.7325286865234,
-24.4261989593506,5.99952650070190,
33.3474388122559,-3.84887814521790,
65.9015045166016,2.44834184646606,
37.1550331115723,10.7052822113037,
-11.4413642883301,5.90763139724731,
-27.4543609619141,-3.19251680374146,
-8.90593528747559,-1.06839275360107,
11.5890083312988,6.05287313461304,
19.1023597717285,0.638836562633514,
19.6700000762939,-7.28247880935669,
13.7369260787964,9.88312721252441,
-4.13908100128174,51.6198616027832,
-20.2644004821777,80.8476257324219,
-22.9504795074463,72.9516983032227,
-22.6714363098145,47.9245452880859,
-38.4180564880371,38.3812141418457,
-60.4092521667481,37.5793838500977,
-55.5092811584473,15.5625181198120,
-8.66223526000977,-23.8157844543457,
43.2099151611328,-42.0056991577148,
56.8831176757813,-26.7455806732178,
42.8444747924805,-12.6224231719971,
33.6942481994629,-20.1258163452148,
38.4480667114258,-18.3622589111328,
36.6588668823242,15.8702278137207,
12.6816186904907,49.5544548034668,
-22.1865272521973,34.2010650634766,
-48.6247482299805,-17.6028633117676,
-51.2811431884766,-36.5283584594727,
-27.4017715454102,3.26144218444824,
4.62853813171387,42.2987861633301,
12.9041881561279,24.5826816558838,
-19.3770751953125,-21.7690715789795,
-58.1471862792969,-30.7466011047363,
-50.4528160095215,-2.83511495590210,
8.91438293457031,4.93156671524048,
56.5470314025879,-20.2839450836182,
48.2386093139648,-22.2871627807617,
14.2982940673828,27.1948280334473,
-4.21607828140259,70.9644622802734,
-13.8307008743286,44.7748603820801,
-39.9104537963867,-21.3519287109375,
-59.0393676757813,-44.1711044311523,
-28.4557533264160,-4.54818010330200,
34.7612686157227,28.9532833099365,
54.8768539428711,11.6258430480957,
1.77689647674561,-13.7591199874878,
-55.7517127990723,2.13799834251404,
-52.9658164978027,35.8341331481934,
-19.9349803924561,32.9965972900391,
-23.0956249237061,-1.42375493049622,
-51.1199684143066,-21.6306095123291,
-38.1099090576172,-7.93434333801270,
20.9237155914307,11.3588113784790,
51.0698165893555,16.0176162719727,
14.5135049819946,15.2419624328613,
-33.1605339050293,10.9238252639771,
-26.8866748809814,-15.0914964675903,
11.6815919876099,-59.3428611755371,
13.4821434020996,-72.0282211303711,
-25.0793399810791,-27.5115566253662,
-44.9706802368164,27.3476467132568,
-18.8200073242188,34.4153785705566,
8.24252986907959,-4.23667621612549,
-4.79234552383423,-37.6096534729004,
-27.7620830535889,-40.3307113647461,
-13.6192188262939,-36.0213546752930,
27.4042224884033,-47.4262657165527,
49.4073410034180,-57.8882179260254,
32.1999359130859,-43.7034530639648,
1.91161704063416,-15.4524822235107,
-12.3408708572388,3.87704968452454,
-11.7328481674194,12.6533164978027,
-16.4875774383545,20.4299793243408,
-27.5865306854248,20.2244930267334,
-25.0479164123535,0.113557934761047,
-1.65324139595032,-25.8818569183350,
30.9744224548340,-26.9866828918457,
49.0723114013672,-0.868689775466919,
37.8743591308594,23.8122615814209,
4.76881217956543,23.1720352172852,
-18.5329627990723,7.35638952255249,
-9.94042205810547,6.37268066406250,
15.5099992752075,20.9933147430420,
26.8503189086914,28.3779830932617,
20.3055992126465,17.9760589599609,
17.7323226928711,2.75964403152466,
28.9000473022461,-6.31367778778076,
32.2255897521973,-13.7235937118530,
4.73792028427124,-17.8128604888916,
-35.8327598571777,-11.4252920150757,
-51.8334312438965,5.70119714736939,
-38.9132957458496,17.0104370117188,
-30.2504138946533,12.9244537353516,
-31.3743247985840,8.53421974182129,
-13.2866210937500,18.4049377441406,
32.4756355285645,30.2458801269531,
65.6776275634766,15.5395336151123,
45.3619003295898,-22.2633037567139,
-1.36404800415039,-45.4514350891113,
-14.1068410873413,-42.5854682922363,
13.1417284011841,-36.9380874633789,
28.8220138549805,-41.5681266784668,
5.51105213165283,-34.3081016540527,
-18.6572341918945,1.81980741024017,
-0.827805161476135,40.9749183654785,
29.7555255889893,40.3531341552734,
14.5170879364014,5.63282871246338,
-40.4712829589844,-18.9589366912842,
-69.8356323242188,-19.3189983367920,
-40.0822067260742,-21.3349685668945,
14.9441461563110,-37.1167640686035,
44.1121520996094,-36.3619003295898,
43.8298912048340,-6.71093082427979,
36.9890060424805,9.90077686309815,
33.8847579956055,-20.9357490539551,
30.0370903015137,-60.6513442993164,
23.7515945434570,-46.7275543212891,
21.7842884063721,12.7271909713745,
9.48929119110107,45.4559211730957,
-23.8217792510986,12.0369024276733,
-51.4655952453613,-39.3125724792481,
-34.6407890319824,-43.1594924926758,
12.5389537811279,-0.972715377807617,
37.1478462219238,36.2870521545410,
19.0086498260498,45.8079071044922,
-10.2860355377197,38.8785858154297,
-19.0820007324219,23.1781425476074,
-17.9489498138428,-2.77729654312134,
-31.4699077606201,-25.0189647674561,
-36.9761695861816,-20.8864707946777,
2.63078689575195,1.15561306476593,
58.1631164550781,13.4682178497314,
62.3408317565918,8.25892353057861,
7.70784568786621,5.66706895828247,
-36.3437500000000,12.3643579483032,
-24.5004558563232,7.04261064529419,
3.43898820877075,-24.9421367645264,
-10.9094495773315,-52.5965309143066,
-40.8152465820313,-37.6610374450684,
-19.7857151031494,2.80100774765015,
42.9726524353027,26.7082328796387,
64.7146759033203,24.0434284210205,
8.83983325958252,16.9555568695068,
-50.5822944641113,14.7979803085327,
-33.8852462768555,2.27806401252747,
28.7601604461670,-19.9870471954346,
40.8420982360840,-26.9281139373779,
-19.7745323181152,-12.3288202285767,
-71.8793792724609,-1.27019524574280,
-50.5304908752441,-13.7358980178833,
5.82496356964111,-24.8836574554443,
21.5096836090088,-2.95179557800293,
-23.4030952453613,30.2254257202148,
-68.7000122070313,24.7617835998535,
-60.9528045654297,-24.5092697143555,
-18.8332519531250,-66.0970993041992,
5.61756610870361,-63.7397003173828,
-5.84000110626221,-36.5917053222656,
-22.2432327270508,-19.3960437774658,
-10.0115222930908,-17.3176040649414,
30.1767082214355,-12.3552789688110,
56.4673118591309,-9.23470211029053,
37.5229644775391,-24.4186172485352,
0.653633356094360,-48.3888778686523,
-4.13890314102173,-47.9243736267090,
25.3546848297119,-15.2972545623779,
37.3237800598145,11.9990663528442,
-5.24266386032105,5.71156978607178,
-68.8028030395508,-15.4578313827515,
-78.8197097778320,-15.7634992599487,
-21.5623359680176,-3.01737761497498,
33.7636528015137,-9.43494796752930,
28.9389133453369,-38.9314956665039,
-6.63722085952759,-53.0841407775879,
-8.44890022277832,-25.1963825225830,
29.8698253631592,21.8257942199707,
47.9022560119629,43.1851577758789,
12.2481298446655,28.7986068725586,
-33.8665351867676,8.04813003540039,
-30.4820251464844,2.61620330810547,
10.9613456726074,2.85187697410584,
33.6187934875488,-8.11061286926270,
8.01595401763916,-26.1820755004883,
-30.5023841857910,-34.9000892639160,
-39.9439315795898,-21.4625663757324,
-24.6540393829346,10.3986330032349,
-15.7051668167114,42.6023178100586,
-23.7752914428711,57.8656997680664,
-30.3002452850342,52.6653900146484,
-22.0182304382324,34.2201385498047,
-4.88971185684204,12.1836032867432,
11.0687379837036,-11.4104232788086,
19.0595836639404,-31.7304725646973,
20.1282424926758,-37.8445701599121,
20.0741233825684,-16.1466655731201,
28.2783527374268,15.4282560348511,
50.7970619201660,26.8857612609863,
69.4773635864258,12.6670331954956,
53.6841163635254,0.300021111965179,
1.66182279586792,9.53542995452881,
-45.3046417236328,17.2898197174072,
-48.5351638793945,-3.85904312133789,
-22.4473590850830,-41.8468894958496,
-10.3838176727295,-51.6403007507324,
-28.7042369842529,-20.2056903839111,
-48.0585975646973,15.8866615295410,
-42.0734786987305,20.4346542358398,
-23.6929588317871,4.18015384674072,
-22.1085147857666,5.83107519149780,
-34.5758972167969,29.5041790008545,
-30.2161369323730,46.7624855041504,
0.365286350250244,40.0669746398926,
32.4862365722656,19.2778301239014,
42.3464202880859,-2.77670383453369,
23.3196010589600,-25.9656829833984,
-10.1499013900757,-44.0406379699707,
-39.1892433166504,-44.3386421203613,
-41.1890182495117,-25.2629528045654,
-15.8312816619873,-12.5952434539795,
6.84615373611450,-25.7971935272217,
-1.11833095550537,-43.6203536987305,
-28.9379005432129,-29.7054080963135,
-35.2128677368164,7.15815067291260,
-7.22789859771729,19.8591308593750,
10.0373430252075,-4.53277015686035,
-17.6886215209961,-23.9226226806641,
-52.2246170043945,-8.90345478057861,
-33.7716865539551,13.7123098373413,
29.5817565917969,3.98084926605225,
65.4702529907227,-18.9299716949463,
43.7395629882813,-3.51446938514709,
7.27801799774170,44.4342155456543,
5.79692935943604,59.2127952575684,
23.1426715850830,17.6017837524414,
21.2949409484863,-18.8932685852051,
3.54877424240112,5.49946880340576,
-0.799350023269653,51.9761238098145,
8.18376541137695,44.6236152648926,
-6.22853755950928,-13.9134359359741,
-47.8104438781738,-45.7307319641113,
-76.6094055175781,-20.1141376495361,
-63.3191413879395,9.51214694976807,
-30.7180747985840,-9.22371101379395,
-4.31348609924316,-45.0531349182129,
15.9317283630371,-39.3547744750977,
34.3943939208984,2.85233235359192,
38.4413452148438,21.2524929046631,
26.1279315948486,0.591148972511292,
23.8022594451904,-13.2944192886353,
44.9266662597656,6.24682521820068,
55.3824996948242,33.7892227172852,
16.9838542938232,39.2930755615234,
-49.2016296386719,24.9085464477539,
-78.5969696044922,7.19458675384522,
-56.8732986450195,-12.8076333999634,
-38.9389038085938,-35.5472831726074,
-56.4303283691406,-40.8597793579102,
-67.9577713012695,-15.6752920150757,
-29.2370071411133,17.8110523223877,
30.8792762756348,25.8305492401123,
48.4436874389648,19.7921619415283,
11.0562591552734,35.6275138854981,
-29.0902557373047,60.3834037780762,
-34.6883354187012,43.5692901611328,
-20.7981491088867,-20.0403900146484,
-10.2048673629761,-68.5097885131836,
3.53126597404480,-49.6782302856445,
28.6478137969971,8.10090446472168,
39.0375976562500,32.7468032836914,
6.58071041107178,-0.578115582466126,
-39.3986854553223,-46.8567733764648,
-42.2440719604492,-65.4698486328125,
3.12308979034424,-53.6309509277344,
49.1259918212891,-28.4418201446533,
49.0123939514160,2.44215703010559,
10.4880695343018,25.4471645355225,
-26.3657131195068,13.0279312133789,
-32.2984886169434,-35.4429359436035,
-13.2544250488281,-72.2584381103516,
12.7689914703369,-56.2752265930176,
23.9462471008301,-3.51560759544373,
5.24738216400147,29.7924709320068,
-31.5527820587158,19.6820793151855,
-42.1108551025391,-8.33907032012940,
-6.63792705535889,-11.7348299026489,
34.2578239440918,16.2999553680420,
26.8718605041504,50.3474349975586,
-20.5867938995361,66.1709060668945,
-42.0595436096191,58.8479576110840,
-2.33343744277954,36.4381904602051,
49.2696990966797,17.2038173675537,
45.7161750793457,11.5431451797485,
0.693902730941773,9.91904926300049,
-13.4225835800171,-4.73256921768189,
25.8426971435547,-26.0206604003906,
62.4398536682129,-28.8702812194824,
53.8582572937012,-10.3504295349121,
29.5674934387207,3.45480227470398,
36.3406639099121,-2.89917850494385,
54.4744682312012,-10.6628532409668,
28.0137977600098,1.03861916065216,
-36.8017997741699,15.7751350402832,
-65.6174163818359,-0.704109668731690,
-19.8348426818848,-36.7840347290039,
45.4647026062012,-37.1842308044434,
50.8896598815918,12.8264636993408,
-5.30700349807739,59.6592369079590,
-55.0539131164551,47.1512908935547,
-55.2105751037598,-6.70308828353882,
-30.4418144226074,-43.2759819030762,
-12.0395107269287,-39.5591583251953,
-2.71661043167114,-27.3821048736572,
9.52474689483643,-32.8166923522949,
21.5024948120117,-42.2973899841309,
20.0016326904297,-36.8707351684570,
4.53704547882080,-28.4539947509766,
-2.18940401077271,-32.2977981567383,
11.1124191284180,-32.0363540649414,
30.7986812591553,-4.42543077468872,
33.0712738037109,32.3631896972656,
12.0932083129883,34.4157333374023,
-14.1735048294067,-2.89992213249207,
-14.1332893371582,-32.4807701110840,
25.4594326019287,-18.1027278900147,
70.9817428588867,17.6257286071777,
72.4985961914063,29.1272792816162,
23.2575302124023,11.5800647735596,
-33.5104026794434,-2.14245247840881,
-53.2353668212891,2.97650575637817,
-41.7036705017090,-0.751783967018127,
-32.2697029113770,-25.4326877593994,
-36.3056716918945,-44.8847999572754,
-29.3320789337158,-31.0309581756592,
-2.49297356605530,-4.36064529418945,
17.1118507385254,0.720172882080078,
12.2796936035156,-12.6180467605591,
1.29394936561584,-7.27705955505371,
8.96021556854248,24.2700176239014,
21.9814319610596,44.2643127441406,
8.59750366210938,18.4129199981689,
-20.8991565704346,-31.8436679840088,
-26.3577728271484,-58.5666770935059,
3.07636690139771,-51.5588226318359,
28.6030464172363,-41.0771980285645,
20.5952415466309,-48.5433540344238,
0.522539854049683,-62.9043540954590,
12.4942836761475,-62.1770210266113,
54.9062881469727,-39.5576553344727,
78.6625213623047,-7.49373722076416,
53.2584648132324,16.4606037139893,
-2.67627358436584,19.9723224639893,
-45.9124794006348,6.33415699005127,
-55.2609443664551,-9.22240734100342,
-32.3825912475586,-8.53036975860596,
13.7647848129272,5.24537897109985,
59.5382347106934,12.7199449539185,
66.4430541992188,3.82007646560669,
23.6220054626465,-4.56958723068237,
-31.9169750213623,-0.204447060823441,
-44.4951477050781,3.06301760673523,
-4.24526453018189,-7.56839179992676,
35.6040191650391,-25.7395019531250,
18.5862216949463,-25.7068176269531,
-40.0936012268066,-5.36976718902588,
-75.9772033691406,10.4781932830811,
-50.0002212524414,2.96714425086975,
6.95596599578857,-11.1595706939697,
35.1198577880859,-7.64735126495361,
8.39624404907227,12.2181358337402,
-30.5542068481445,25.3205051422119,
-28.5669555664063,22.6469364166260,
19.2722339630127,18.8381385803223,
65.4821624755859,23.9873371124268,
61.6634521484375,24.0347938537598,
20.1824398040772,-0.0417905449867249,
-9.36265945434570,-37.7132606506348,
6.11598920822144,-55.2529716491699,
45.4424705505371,-34.2781219482422,
60.6204338073731,8.73540019989014,
35.5206832885742,38.4618339538574,
-2.45316600799561,38.3347396850586,
-21.2857627868652,21.1216239929199,
-19.4898109436035,6.80942344665527,
-14.1249933242798,1.85114061832428,
-23.3750114440918,4.57210636138916,
-40.5642433166504,12.8028488159180,
-48.7978096008301,20.8086109161377,
-37.5340080261231,20.1062927246094,
-12.1748008728027,1.73144912719727,
15.3181238174438,-27.9234161376953,
28.7064933776855,-42.8593940734863,
25.9714984893799,-24.5099983215332,
13.7138299942017,15.7982931137085,
4.50386047363281,43.1223678588867,
1.74563956260681,39.9483146667481,
-5.62158060073853,18.1531696319580,
-25.9580898284912,10.3244562149048,
-47.5653877258301,26.5494537353516,
-52.2574615478516,42.1668052673340,
-34.0506553649902,33.4315185546875,
-8.90535831451416,10.7275876998901,
7.05942678451538,7.56114339828491,
16.3741245269775,30.6334571838379,
31.6717967987061,47.5604858398438,
48.4533233642578,31.3479461669922,
48.2292900085449,-3.89909029006958,
31.4151096343994,-22.9707126617432,
15.3666162490845,-18.9867515563965,
8.59644126892090,-20.3377246856689,
1.95719015598297,-39.2257423400879,
-14.6795053482056,-51.2221527099609,
-29.3362865447998,-33.1788177490234,
-23.8534049987793,-6.91626548767090,
-2.69388198852539,-4.77412319183350,
14.2513542175293,-19.7523403167725,
24.3900451660156,-16.0839996337891,
33.4281196594238,18.6373348236084,
34.7148056030273,53.8119468688965,
8.89911365509033,65.6648025512695,
-30.3938751220703,62.1492652893066,
-40.5054931640625,58.1540908813477,
-6.39543533325195,46.5418281555176,
25.9816055297852,17.5083885192871,
7.23579692840576,-12.3829421997070,
-45.7695465087891,-20.5975761413574,
-69.5440826416016,-17.2750244140625,
-36.2115058898926,-35.3846015930176,
9.99213790893555,-72.9887847900391,
15.3013772964478,-86.2243804931641,
-14.4832468032837,-51.6363945007324,
-34.4562492370606,2.33608555793762,
-28.2885189056397,30.3251857757568,
-16.2920570373535,23.8693046569824,
-16.7182712554932,10.4117507934570,
-25.8405685424805,16.4363307952881,
-29.1512794494629,34.3758163452148,
-20.1538143157959,42.5672836303711,
2.60532760620117,38.7064056396484,
32.6635665893555,28.9934425354004,
49.7027778625488,25.8666973114014,
37.2516860961914,34.4246215820313,
8.31943798065186,46.1751060485840,
-3.10811471939087,38.1275825500488,
18.7825374603272,5.69221544265747,
36.8419837951660,-21.5193691253662,
17.8550090789795,-7.76110172271729,
-16.8933105468750,25.7226219177246,
-24.1613292694092,25.6859283447266,
0.536808967590332,-27.2870998382568,
18.2709922790527,-75.7667160034180,
6.04774951934814,-52.1447334289551,
-16.0247688293457,20.9113655090332,
-20.5178775787354,56.4883880615234,
-12.3582429885864,19.2831153869629,
-10.3687391281128,-29.6828804016113,
-10.6736135482788,-27.9286270141602,
-3.09253478050232,10.3066492080688,
-6.61948108673096,23.6327877044678,
-38.6923866271973,-1.80931162834167,
-75.0930023193359,-29.2736968994141,
-65.1112442016602,-38.3907966613770,
-7.95355892181397,-48.0334968566895,
38.9919815063477,-61.2740859985352,
40.5339508056641,-47.8621788024902,
23.8360843658447,4.40858173370361,
31.0277347564697,48.9040298461914,
54.1240615844727,37.9267959594727,
53.2407646179199,-7.29302644729614,
21.7203121185303,-23.8282546997070,
-4.28929376602173,-1.16092967987061,
-7.62288522720337,14.0749645233154,
-14.5271482467651,-4.95488500595093,
-38.6338005065918,-33.8415145874023,
-54.9135856628418,-35.4807167053223,
-42.4813842773438,-9.16561317443848,
-18.6756572723389,13.1242685317993,
-7.65332984924316,18.8808917999268,
-3.29420471191406,17.5388183593750,
14.3528633117676,9.24765014648438,
31.0657386779785,-9.38922119140625,
25.4566783905029,-23.2550067901611,
5.05928039550781,-18.4238395690918,
4.98396825790405,-8.90710544586182,
25.6085815429688,-10.7259788513184,
27.6533946990967,-9.48123931884766,
-8.64135265350342,16.6733989715576,
-40.1271247863770,49.4790077209473,
-24.8020992279053,39.2890014648438,
18.7318592071533,-19.1939792633057,
37.3784866333008,-58.1468849182129,
17.5245075225830,-23.3273944854736,
-3.39994025230408,39.2540435791016,
0.442335724830627,40.3443908691406,
21.9211330413818,-17.1757526397705,
36.4425010681152,-43.1615676879883,
36.5592575073242,6.01282024383545,
28.4531269073486,61.6363105773926,
18.5019607543945,41.9118995666504,
9.81419277191162,-25.9865016937256,
10.2445678710938,-52.9010314941406,
16.4136848449707,-14.1099300384521,
17.4798870086670,21.4050312042236,
12.8718414306641,9.45446777343750,
16.6641235351563,-11.2860069274902,
21.7597351074219,2.03569412231445,
0.779854774475098,23.7492160797119,
-39.3457717895508,5.75985622406006,
-54.0312767028809,-33.8107070922852,
-17.7872409820557,-32.5292358398438,
29.9075546264648,12.3307685852051,
30.2458496093750,39.1161994934082,
-9.49984931945801,13.7287588119507,
-22.9326591491699,-24.2084903717041,
18.4706306457520,-28.7161388397217,
59.7473068237305,-10.5300216674805,
48.2621612548828,-18.4401435852051,
11.4270858764648,-51.4203948974609,
9.20439529418945,-58.0819358825684,
38.7201080322266,-20.1388511657715,
37.6125869750977,21.6574821472168,
-16.8026275634766,23.9856891632080,
-69.9393615722656,-10.9924259185791,
-61.9013519287109,-43.2785949707031,
-5.69057941436768,-44.5354804992676,
38.9161071777344,-18.8191719055176,
43.1209640502930,3.32946562767029,
25.2655200958252,2.90795779228210,
11.4519824981689,-6.77194166183472,
-0.818914830684662,5.05451345443726,
-13.9503202438355,48.5668487548828,
-13.9423875808716,91.7218093872070,
2.13689112663269,80.9313430786133,
14.1360902786255,15.8151988983154,
9.29916286468506,-35.5186729431152,
1.55948328971863,-20.2129783630371,
4.98669147491455,27.7605781555176,
11.2654981613159,46.3575744628906,
6.14545869827271,30.9387283325195,
-5.85458803176880,29.1611099243164,
-7.94299602508545,57.1394500732422,
-6.27524805068970,69.4110107421875,
-27.8495445251465,29.7398929595947,
-63.8012580871582,-22.3523559570313,
-68.3585281372070,-35.4663429260254,
-30.1505088806152,-24.1901760101318,
8.07592296600342,-36.7126083374023,
6.90470361709595,-67.0027236938477,
-12.9709186553955,-57.5342521667481,
-8.44133090972900,-5.31798458099365,
15.7701673507690,23.5182876586914,
19.0175113677979,-8.35774993896484,
-4.69037103652954,-45.8528442382813,
-10.6049442291260,-28.5520553588867,
14.1191339492798,18.4128379821777,
28.2474250793457,24.9736862182617,
5.26050043106079,-21.7974376678467,
-13.5627479553223,-55.7706680297852,
10.3055934906006,-37.2463722229004,
38.8168716430664,-0.376169681549072,
9.89047813415527,8.83919715881348,
-58.4105072021484,-5.61699390411377,
-81.2659072875977,-20.5910644531250,
-30.0753974914551,-38.5546798706055,
24.9303112030029,-61.3960876464844,
16.5528526306152,-60.3790473937988,
-21.8779850006104,-15.6437311172485,
-12.6538372039795,37.0248260498047,
46.2046852111816,48.1025466918945,
81.3366470336914,21.4035644531250,
59.9739227294922,10.8138446807861,
26.1472682952881,38.7520446777344,
21.0193214416504,62.6730041503906,
26.7695980072022,35.8683929443359,
12.3899250030518,-24.2097606658936,
-3.46121168136597,-61.3602256774902,
15.1478815078735,-55.7695541381836,
55.1299705505371,-23.9249248504639,
62.1693267822266,6.96957683563232,
19.2958583831787,17.9385738372803,
-29.7757034301758,2.35046386718750,
-40.0035209655762,-28.9824638366699,
-24.7128868103027,-47.2495613098145,
-11.8652563095093,-31.6619510650635,
1.00749778747559,-0.172723531723022,
25.8795013427734,18.1495971679688,
47.7435035705566,18.1939601898193,
36.4387321472168,19.6928749084473,
-4.50035667419434,29.3181514739990,
-37.8009681701660,17.9234676361084,
-37.7014923095703,-27.4763259887695,
-19.9920425415039,-66.9685058593750,
-16.7913990020752,-57.8209228515625,
-30.4353771209717,-11.2837476730347,
-38.5899658203125,28.8356113433838,
-27.4371452331543,35.0088729858398,
-1.31667470932007,21.8596229553223,
29.7662315368652,9.90424537658691,
47.9265594482422,-0.218279242515564,
36.6716766357422,-7.85913419723511,
5.56268882751465,-0.512928724288940,
-21.0078754425049,17.9066352844238,
-26.8841342926025,18.8055953979492,
-24.5894412994385,-16.7533035278320,
-30.9740200042725,-54.7009353637695,
-34.1086616516113,-45.4136276245117,
-11.6053495407105,-1.45190882682800,
23.7016429901123,18.3286437988281,
27.9366893768311,-13.1843976974487,
-6.64878273010254,-50.0381011962891,
-34.4186744689941,-39.3339233398438,
-22.5122528076172,8.78429222106934,
-3.90505218505859,36.8465347290039,
-22.8554897308350,18.9916419982910,
-63.3236045837402,-12.7539768218994,
-65.5134582519531,-24.5054206848145,
-16.9453582763672,-19.3208103179932,
24.6356029510498,-8.02361679077148,
14.2878074645996,9.31103897094727,
-19.6808395385742,26.7731418609619,
-20.9405345916748,16.3015003204346,
10.7455253601074,-30.0719814300537,
30.8462486267090,-72.0681762695313,
23.8196296691895,-63.9194412231445,
13.5168304443359,-15.1988315582275,
16.9755973815918,23.8048362731934,
15.8778762817383,24.7997627258301,
1.06125974655151,12.0446653366089,
-11.6724920272827,9.28415775299072,
-9.18048667907715,-1.33013391494751,
-0.423087596893311,-34.3288002014160,
5.18188810348511,-63.4542121887207,
21.7346744537354,-54.0861587524414,
56.7231140136719,-14.0817356109619,
79.3518676757813,19.9856777191162,
50.1072769165039,32.6560783386231,
-14.3946647644043,36.9159851074219,
-49.1238136291504,35.9319763183594,
-27.4483089447022,17.9224281311035,
13.4350843429565,-11.4851531982422,
32.4672126770020,-17.1451625823975,
34.4975395202637,15.2302942276001,
39.2821197509766,47.1458244323731,
43.0903434753418,36.1171073913574,
25.5053710937500,-5.96309089660645,
-3.60172033309937,-34.8526344299316,
-11.8316411972046,-35.5011978149414,
8.71366119384766,-25.3103942871094,
32.1944618225098,-15.9725475311279,
38.3305511474609,1.11593401432037,
34.8121910095215,22.7041473388672,
26.1864337921143,28.5126781463623,
4.94969511032105,13.5040321350098,
-28.9301471710205,8.97079086303711,
-44.0128479003906,35.3020896911621,
-24.4509391784668,61.3338050842285,
0.418612897396088,46.8467788696289,
-8.27908611297607,1.54608035087585,
-48.3534851074219,-21.3303966522217,
-74.8747787475586,-5.00452709197998,
-58.2805213928223,6.05402469635010,
-18.0962104797363,-20.0399475097656,
9.26035881042481,-54.5060119628906,
15.3121690750122,-46.6835098266602,
18.2611370086670,2.50227189064026,
28.8565406799316,36.7844848632813,
39.1838912963867,25.4585552215576,
40.9480590820313,-0.0191547870635986,
31.2923679351807,8.47343158721924,
16.0435848236084,46.3939971923828,
2.29602241516113,66.1346511840820,
-2.02343726158142,40.6414031982422,
3.13557386398315,-5.86915779113770,
8.52777385711670,-33.2211189270020,
10.2550945281982,-25.4665679931641,
8.06478977203369,1.37686133384705,
2.35195302963257,18.2164859771729,
-7.70670366287231,14.2900829315186,
-24.6398200988770,0.837054312229157,
-32.6919975280762,-6.33595848083496,
-15.4816856384277,-5.05081510543823,
15.4913892745972,-5.48044061660767,
28.4386520385742,-20.9900779724121,
14.3074169158936,-38.3310546875000,
-1.76584851741791,-32.1532783508301,
3.75574135780334,-0.0834062099456787,
19.3892765045166,31.7264366149902,
17.0418796539307,44.2590522766113,
1.20491456985474,47.7626113891602,
2.71168184280396,52.3410949707031,
26.1387157440186,50.8535728454590,
32.1085433959961,25.8864288330078,
-7.75529623031616,-7.81991386413574,
-56.1348991394043,-15.4780168533325,
-55.8930168151856,5.96698284149170,
-8.52474975585938,15.8840494155884,
23.9333629608154,-10.1825799942017,
1.90216898918152,-45.1109199523926,
-44.7716445922852,-49.3706474304199,
-60.1467514038086,-29.4932956695557,
-38.7253875732422,-21.4454898834229,
-14.4278497695923,-28.7890567779541,
-10.7483596801758,-20.3004608154297,
-16.7102317810059,9.58917808532715,
-21.2042503356934,26.9061660766602,
-28.3940773010254,7.32599353790283,
-32.7885742187500,-26.9853916168213,
-12.4981374740601,-34.6304664611816,
31.8154125213623,-20.2395744323730,
61.1734848022461,-15.3805522918701,
45.5252380371094,-29.5210723876953,
10.3803453445435,-39.1753349304199,
4.08114480972290,-28.5229549407959,
34.6727371215820,-12.3397998809814,
65.4966964721680,0.150468111038208,
66.6448669433594,15.8589620590210,
50.4754600524902,29.1005859375000,
39.4692306518555,21.0321311950684,
27.0480041503906,-8.87651824951172,
4.91899967193604,-26.9272880554199,
-16.0159149169922,-0.923769950866699,
-15.1980466842651,49.9856414794922,
-0.969789981842041,70.8819732666016,
6.38040685653687,42.5543098449707,
3.29129600524902,1.40499615669250,
3.56001114845276,-14.4468669891357,
9.04918193817139,-0.166613563895226,
3.06367540359497,26.3068885803223,
-15.9606904983521,48.6810035705566,
-25.9151496887207,52.7296066284180,
-11.1627531051636,25.5662231445313,
12.4495544433594,-16.4353637695313,
16.0158710479736,-29.1611804962158,
-2.05080556869507,13.9276638031006,
-23.9314365386963,70.6510848999023,
-40.4764060974121,74.2200698852539,
-55.6702957153320,11.0593357086182,
-60.9968338012695,-50.9803276062012,
-39.7070732116699,-42.4020347595215,
5.84147977828980,23.4057540893555,
43.2675666809082,69.6738052368164,
40.2918815612793,51.8374710083008,
2.43140697479248,-3.87647867202759,
-28.3129444122314,-38.0409355163574,
-22.0247726440430,-26.7845916748047,
16.1157321929932,1.26684546470642,
50.4771270751953,13.1141023635864,
51.8136215209961,9.48798084259033,
19.2464122772217,13.1484889984131,
-23.1414642333984,35.0629653930664,
-43.3753547668457,53.8595046997070,
-28.6897659301758,49.7133750915527,
2.78502798080444,25.9619407653809,
21.7357921600342,4.97484397888184,
16.0712108612061,5.41385841369629,
3.91404104232788,17.4691543579102,
6.86985778808594,19.6394176483154,
26.1303787231445,14.3985309600830,
36.3420715332031,17.6014633178711,
13.0458354949951,30.5827198028564,
-31.5109310150147,41.2428436279297,
-62.1269340515137,35.1170043945313,
-55.1299858093262,19.0865154266357,
-20.0659198760986,13.0360784530640,
8.64252090454102,13.1188058853149,
4.96378707885742,-0.0762408971786499,
-17.4578895568848,-31.5411987304688,
-27.1046791076660,-49.7027664184570,
-7.15001583099365,-29.7222862243652,
18.7155380249023,4.78326463699341,
21.7674674987793,5.92516136169434,
4.78866004943848,-29.1008987426758,
-0.282422840595245,-47.7463836669922,
26.0747604370117,-12.5714817047119,
49.7412414550781,40.0725860595703,
27.3679885864258,46.4563598632813,
-28.0312576293945,-2.07076716423035,
-57.4540367126465,-46.5008583068848,
-35.7992553710938,-40.9885749816895,
-4.32183218002319,-0.487305164337158,
-9.26295280456543,37.7279701232910,
-38.4281463623047,59.9629783630371,
-41.7168731689453,65.9457702636719,
-16.1806411743164,48.1156501770020,
-9.28880023956299,5.26806545257568,
-34.4032211303711,-33.3502960205078,
-41.2483024597168,-34.5726661682129,
8.05860328674316,-6.31291961669922,
70.1498336791992,13.8281850814819,
70.2428054809570,13.1371145248413,
6.98129892349243,10.8729295730591,
-47.7544784545898,20.4448833465576,
-47.1737403869629,22.2170429229736,
-24.0337219238281,2.72970223426819,
-24.2082042694092,-8.34125423431397,
-38.7628746032715,14.8500919342041,
-28.9785041809082,48.3803443908691,
4.75737953186035,49.6604804992676,
19.3757152557373,11.3014678955078,
-3.11357498168945,-23.7159233093262,
-29.8454685211182,-16.6913585662842,
-24.5075836181641,18.8948974609375,
-0.663958847522736,42.8426246643066,
12.1573247909546,27.9612274169922,
7.86510181427002,-12.0908803939819,
2.93235611915588,-45.4918594360352,
2.85337138175964,-42.8511886596680,
1.43673753738403,-1.17224633693695,
-6.28618812561035,44.6415214538574,
-6.47541666030884,47.8360214233398,
9.86036491394043,1.41351413726807,
27.2253532409668,-50.5428009033203,
25.2808475494385,-63.0272979736328,
4.23207855224609,-37.3932952880859,
-15.7405948638916,-9.13164234161377,
-17.8027381896973,0.0636593624949455,
2.49014163017273,-1.63073301315308,
33.1690902709961,0.183131277561188,
52.0902786254883,-4.16789197921753,
47.8654022216797,-20.3498668670654,
33.7157821655273,-31.2647361755371,
26.2669086456299,-19.6147060394287,
30.6884765625000,0.0523121356964111,
30.6689910888672,-2.50870990753174,
15.8864583969116,-27.4549598693848,
5.57124900817871,-38.9842758178711,
18.1958141326904,-19.4722747802734,
39.7591819763184,5.93768882751465,
37.5731315612793,7.51346206665039,
6.62659502029419,-9.23755264282227,
-15.9013195037842,-14.1954345703125,
-8.94724082946777,1.25459086894989,
5.73228406906128,6.40553140640259,
-3.54298329353333,-15.6315393447876,
-23.9696235656738,-46.5646438598633,
-12.7262487411499,-53.9604339599609,
37.0093421936035,-32.9010848999023,
76.0137939453125,-0.952544689178467,
58.6004638671875,21.8124923706055,
-2.64868307113647,24.5499343872070,
-52.1407546997070,6.08149385452271,
-56.7532272338867,-19.5328350067139,
-26.1617660522461,-28.8742027282715,
16.5714817047119,-13.3189029693604,
50.8951873779297,10.7386608123779,
60.4750709533691,15.5159730911255,
39.0174102783203,0.848555207252502,
3.60442709922791,-6.63565158843994,
-19.9862613677979,7.29896306991577,
-21.1039714813232,27.6585426330566,
-15.0748004913330,38.6283340454102,
-13.2801866531372,41.8364639282227,
-4.25672435760498,42.0993270874023,
17.3481025695801,34.6114578247070,
21.5158348083496,21.7531795501709,
-14.2670383453369,15.4546566009521,
-57.6433868408203,22.8409786224365,
-50.2406005859375,22.5960140228272,
2.87100219726563,-2.77320909500122,
34.1186256408691,-32.8578910827637,
4.26431798934937,-33.9186477661133,
-37.1711959838867,-4.92319154739380,
-20.3321456909180,14.0122451782227,
37.5593452453613,2.43598270416260,
58.1635513305664,-7.46965885162354,
13.5446109771729,16.3332328796387,
-35.7411460876465,50.9685134887695,
-36.0062675476074,55.8563919067383,
-13.7045669555664,26.4669456481934,
-19.7940635681152,-1.79963815212250,
-47.2708969116211,0.263853192329407,
-49.2632331848145,20.1550750732422,
-18.4385166168213,33.9599266052246,
9.34974575042725,29.6084613800049,
13.4711570739746,5.48418045043945,
13.1715211868286,-31.1377506256104,
30.0268363952637,-54.4256515502930,
43.2111091613770,-31.4154319763184,
23.8183650970459,20.8336143493652,
-14.1882572174072,34.2579612731934,
-30.0117969512939,-21.0558967590332,
-8.66114997863770,-83.5702209472656,
32.1850738525391,-71.2796325683594,
67.5315322875977,6.76873683929443,
68.6109313964844,57.4017791748047,
26.7233657836914,27.0614376068115,
-22.3655433654785,-29.8428802490234,
-25.4294509887695,-34.9635200500488,
27.1269512176514,3.92679882049561,
72.8512573242188,19.6551055908203,
48.7411422729492,3.67400312423706,
-21.7717895507813,7.88424444198608,
-52.7011184692383,45.9896202087402,
-16.0335655212402,64.5073852539063,
21.8613109588623,25.8849334716797,
2.93896698951721,-23.7447357177734,
-28.5506000518799,-24.7420177459717,
-7.92132949829102,8.34401988983154,
42.6103782653809,12.3338060379028,
49.9535522460938,-26.2194290161133,
1.62907361984253,-57.9250106811523,
-37.2255325317383,-44.9429702758789,
-22.2321987152100,-12.7939653396606,
3.97800683975220,9.01018905639648,
-5.94464588165283,33.5330276489258,
-32.0265998840332,67.1491165161133,
-28.5404968261719,75.8805923461914,
-5.76850032806397,39.0851745605469,
-1.76472020149231,-9.98630142211914,
-10.2454710006714,-20.1217021942139,
15.5143566131592,3.34074974060059,
60.9185028076172,12.3479766845703,
61.5291328430176,-10.6227960586548,
-0.926535606384277,-29.0291385650635,
-53.9375762939453,-19.1243553161621,
-32.0527458190918,-6.51634693145752,
28.9759769439697,-13.8123607635498,
43.3983993530273,-19.7096595764160,
-8.15435218811035,-0.582887887954712,
-58.0894393920898,20.7826328277588,
-54.8210983276367,12.2483386993408,
-27.0487155914307,-12.2009696960449,
-21.8245849609375,-6.40439414978027,
-35.8392677307129,33.5804443359375,
-40.8675842285156,61.3963890075684,
-35.8947601318359,44.2336692810059,
-41.6664619445801,2.24273490905762,
-58.0523071289063,-16.8357143402100,
-61.6751060485840,-2.60038638114929,
-41.5200881958008,13.7113943099976,
-9.74218750000000,11.2172231674194,
11.8424768447876,-2.22855401039124,
18.2435722351074,-10.1865158081055,
14.1437253952026,-1.59005308151245,
-1.26119756698608,18.5055541992188,
-16.7791118621826,27.4744033813477,
-8.88127517700195,9.43506145477295,
18.5772914886475,-16.7239685058594,
29.8208026885986,-12.9509716033936,
9.47990226745606,28.6463851928711,
-22.4983062744141,63.6071243286133,
-32.5997467041016,43.7298622131348,
-23.4423274993897,-12.0260410308838,
-19.6048927307129,-34.3975105285645,
-20.9005298614502,6.32279586791992,
-4.24508380889893,48.6847381591797,
24.3308658599854,29.4247341156006,
26.8542289733887,-25.7867374420166,
-9.26401710510254,-37.9107131958008,
-35.7458381652832,11.2174816131592,
-10.3072605133057,53.5636062622070,
35.4048805236816,30.8860054016113,
32.0914993286133,-27.0324707031250,
-26.0756912231445,-47.7003746032715,
-70.9107589721680,-20.7748908996582,
-49.7264633178711,2.51760005950928,
8.57523155212402,-7.08355855941773,
38.4959373474121,-22.4543228149414,
13.2008285522461,-16.5535030364990,
-31.0028114318848,-5.79611778259277,
-47.6605758666992,-15.9853191375732,
-24.4149799346924,-31.0723953247070,
21.6849822998047,-25.5419445037842,
56.3444938659668,-9.55559349060059,
54.6230697631836,-10.7683048248291,
21.2166385650635,-23.7440547943115,
-2.83164334297180,-11.9954490661621,
7.95688867568970,28.0836524963379,
29.9903526306152,51.5658912658691,
28.7453632354736,28.1219444274902,
10.9660081863403,-7.40060806274414,
12.5461063385010,-11.0328149795532,
38.1124382019043,3.58195114135742,
51.8930397033691,1.02509331703186,
24.7472152709961,-16.3557777404785,
-12.5940265655518,-15.4857406616211,
-16.0579051971436,2.93092656135559,
7.47606897354126,2.49180269241333,
19.7546539306641,-29.9915027618408,
19.2195339202881,-52.1244735717773,
31.6350135803223,-27.7017669677734,
54.5026435852051,17.6279525756836,
51.3351440429688,34.1006126403809,
13.4244365692139,22.8454551696777,
-18.3864231109619,14.8665704727173,
-16.3865756988525,13.7558584213257,
-8.12202835083008,-1.63534712791443,
-31.5912361145020,-25.7029457092285,
-66.6853179931641,-31.8851699829102,
-57.0098457336426,-18.3886909484863,
-1.19993281364441,-13.9838476181030,
42.0479469299316,-25.3739185333252,
39.5741958618164,-18.8770275115967,
25.9002780914307,20.2756614685059,
35.1900634765625,47.3834152221680,
44.1442108154297,19.7701606750488,
17.9491882324219,-26.0900611877441,
-22.4922180175781,-20.5785064697266,
-33.4990997314453,36.2751693725586,
-15.4476499557495,67.6875991821289,
-11.8645153045654,37.1110649108887,
-38.0376014709473,-10.3203191757202,
-50.2560729980469,-16.8938331604004,
-16.5828380584717,5.81697607040405,
26.4279003143311,13.5397186279297,
24.8717994689941,-2.22101449966431,
-15.7243099212646,-8.68203926086426,
-42.6660690307617,9.58485794067383,
-30.9762554168701,25.5548820495605,
1.41716265678406,22.6720466613770,
27.2437095642090,16.4811229705811,
28.0788688659668,19.5158863067627,
3.52380776405334,19.5378780364990,
-37.7082824707031,12.2302999496460,
-62.6462135314941,15.3842353820801,
-43.3291015625000,30.7071743011475,
4.29483318328857,36.3596801757813,
28.2537250518799,20.7176628112793,
7.83895492553711,13.1543912887573,
-13.5720586776733,35.9001350402832,
4.85103416442871,61.6504020690918,
35.7773208618164,39.3470230102539,
31.4075336456299,-21.2097187042236,
1.46469354629517,-50.3178863525391,
-0.826409876346588,-15.3260641098022,
35.7644309997559,32.7936859130859,
59.7528076171875,41.3762817382813,
28.8405151367188,27.6904544830322,
-25.7255096435547,32.5848388671875,
-45.8866348266602,47.5413856506348,
-25.2537536621094,25.7909164428711,
-3.18406677246094,-32.5543174743652,
-0.843707323074341,-70.8517227172852,
-0.884576022624970,-58.8737297058106,
9.06100368499756,-37.8361091613770,
13.4633388519287,-44.9675865173340,
4.76114416122437,-55.8793144226074,
-6.50226593017578,-31.0311813354492,
-11.1506776809692,6.54274749755859,
-13.8665008544922,3.14083385467529,
-16.1461944580078,-34.4332237243652,
-14.2930107116699,-44.4941329956055,
-7.71515560150147,-8.04777812957764,
-12.1833820343018,21.7795982360840,
-28.3105545043945,1.14336836338043,
-31.5254783630371,-36.9766616821289,
-2.05190587043762,-31.3306903839111,
25.5784358978272,9.80768775939941,
9.21991920471191,27.2333259582520,
-36.9095535278320,-3.18886041641235,
-50.9879875183106,-37.7870445251465,
-11.1391925811768,-36.8657531738281,
31.0176181793213,-22.5057353973389,
24.5466289520264,-26.0706577301025,
-8.88052558898926,-39.3218727111816,
-8.14313793182373,-34.3139076232910,
34.2495613098145,-8.53508949279785,
66.3158721923828,10.9928541183472,
52.5531425476074,4.95979261398315,
23.8162212371826,-8.07175827026367,
30.6510467529297,-1.47560381889343,
65.7577209472656,22.8767471313477,
74.3097076416016,41.3111267089844,
28.7492637634277,37.5024566650391,
-36.1607856750488,14.3312063217163,
-67.9188079833984,-8.19799041748047,
-52.2216377258301,-5.48125505447388,
-17.7557888031006,23.2967052459717,
0.829013764858246,43.7777099609375,
3.42039489746094,24.5747337341309,
15.1398792266846,-19.9620265960693,
43.0988311767578,-36.7030639648438,
63.8974609375000,0.00838851928710938,
47.1101455688477,58.0494308471680,
-1.39788627624512,76.0171279907227,
-35.7987136840820,41.1579933166504,
-18.8023643493652,0.633945584297180,
24.1904964447022,-1.12862062454224,
32.5135993957520,29.5350856781006,
-11.5521411895752,59.3985595703125,
-59.6866264343262,69.5222549438477,
-61.7192192077637,61.4411048889160,
-26.2793006896973,38.3969841003418,
-7.47240257263184,7.41268920898438,
-27.3847675323486,-18.1707324981689,
-44.3871459960938,-24.3600444793701,
-21.0918273925781,-24.6274738311768,
22.0233039855957,-42.1918029785156,
37.4460144042969,-68.7766418457031,
16.8038005828857,-69.1426696777344,
-5.97873449325562,-31.7700138092041,
-9.52677345275879,8.29919433593750,
-14.9104890823364,10.4479331970215,
-40.6774063110352,-14.6916666030884,
-64.6700744628906,-30.0433139801025,
-58.3005332946777,-31.4415149688721,
-24.1154785156250,-43.9661979675293,
7.20808124542236,-66.5786437988281,
18.7852230072022,-62.7830848693848,
21.7430458068848,-9.29059219360352,
24.0720520019531,56.4388618469238,
14.6073837280273,79.1928482055664,
-9.04785919189453,49.1703147888184,
-25.8178138732910,8.85470867156982,
-20.2312450408936,-3.99337887763977,
-3.11464095115662,7.12347555160523,
7.09841442108154,19.9941291809082,
9.48548793792725,15.1909370422363,
5.86688852310181,-12.6553115844727,
-9.37460231781006,-46.2195930480957,
-39.5168380737305,-53.0125160217285,
-60.6159095764160,-21.9070320129395,
-40.6208610534668,15.1188840866089,
14.6888580322266,20.9289207458496,
53.4772377014160,-1.00248730182648,
43.9142532348633,-5.08727693557739,
7.04382324218750,26.6581420898438,
-20.3168163299561,52.4457435607910,
-29.2086925506592,27.8496513366699,
-34.1478195190430,-17.5144100189209,
-36.9785995483398,-18.6674289703369,
-31.1926364898682,21.7788333892822,
-25.8153915405273,41.2914505004883,
-35.3435287475586,13.2609519958496,
-49.7004814147949,-15.2341156005859,
-38.4351577758789,0.558195948600769,
0.745197534561157,25.9317855834961,
29.9524269104004,3.24455547332764,
20.4515647888184,-46.5263137817383,
-6.65925884246826,-48.8829383850098,
-8.05025100708008,10.8395462036133,
13.8510484695435,55.7262496948242,
27.9366111755371,29.6149330139160,
23.3272590637207,-22.9712848663330,
12.6561079025269,-30.6442565917969,
10.6616973876953,-0.746506690979004,
11.3996286392212,9.02235031127930,
7.41647291183472,-10.0144844055176,
3.55789017677307,-8.73889350891113,
3.55079746246338,29.8494606018066,
0.214782267808914,60.1772804260254,
-4.49125289916992,45.2719535827637,
6.22012710571289,11.6004114151001,
28.3503799438477,4.81333923339844,
23.9428615570068,16.9900455474854,
-23.6367893218994,8.24603843688965,
-67.9597930908203,-17.8825950622559,
-53.3855247497559,-24.9551029205322,
11.2409448623657,-12.2027921676636,
59.7314758300781,-10.5975303649902,
56.6199989318848,-24.4452228546143,
33.7518119812012,-26.5049648284912,
30.5347843170166,1.58419346809387,
28.3809719085693,36.0297508239746,
-7.58136034011841,45.9488792419434,
-56.9895744323731,34.0265045166016,
-62.9068489074707,18.1500244140625,
-22.6638622283936,-1.79349315166473,
5.38927173614502,-23.4131813049316,
-12.6489620208740,-22.0695190429688,
-38.6797294616699,16.0999584197998,
-22.6647357940674,51.0702056884766,
20.7240085601807,32.8720741271973,
38.6870346069336,-17.1776771545410,
21.4134254455566,-31.1475448608398,
4.34415912628174,15.0251235961914,
11.4650058746338,66.5968246459961,
18.9636669158936,65.5061798095703,
5.25789880752564,21.1291332244873,
-5.53086900711060,-16.5500431060791,
5.84225177764893,-26.6520824432373,
19.0469055175781,-30.9411125183105,
2.84017753601074,-39.7951240539551,
-26.6305522918701,-39.9751358032227,
-26.9561462402344,-27.1440296173096,
6.07846212387085,-12.0075254440308,
30.4312191009522,1.49320983886719,
16.2381362915039,26.0378303527832,
-13.2754917144775,56.0404701232910,
-24.7157325744629,63.4789581298828,
-21.2138500213623,42.2744064331055,
-24.0334339141846,19.4552307128906,
-25.6735000610352,19.9861965179443,
-4.58899021148682,31.0464286804199,
28.2573566436768,20.5733699798584,
40.1243095397949,-18.6210727691650,
24.8686027526855,-51.3408164978027,
10.2571649551392,-47.5949935913086,
14.8575553894043,-14.3493556976318,
15.8231420516968,20.0900535583496,
-10.6202602386475,29.3983612060547,
-43.0004043579102,8.17015457153320,
-41.9854660034180,-29.3020992279053,
-8.11864757537842,-49.3200607299805,
19.8634319305420,-34.3853340148926,
19.4814453125000,-2.16383957862854,
8.17094039916992,11.2736759185791,
0.323702812194824,1.58618640899658,
-13.0477914810181,-3.18916511535645,
-38.1706314086914,15.7581071853638,
-48.1365013122559,32.4809112548828,
-20.0500144958496,14.4092607498169,
28.5605564117432,-27.3527832031250,
55.9389305114746,-41.8465728759766,
46.4071884155273,-9.65149688720703,
31.3333835601807,31.3069610595703,
35.7836532592773,41.9783134460449,
43.2271080017090,25.3712329864502,
27.8432140350342,14.4283428192139,
-7.09367179870606,21.0947208404541,
-31.7612476348877,27.5789852142334,
-30.5777797698975,20.7798137664795,
-11.0790319442749,9.74176216125488,
3.87254548072815,3.06571841239929,
0.0338527262210846,0.816664993762970,
-22.0168132781982,-0.161907196044922,
-43.3875312805176,6.27636146545410,
-37.9936599731445,25.7442893981934,
0.152727529406548,40.9228515625000,
39.8706321716309,31.8877792358398,
38.6183929443359,2.86082267761230,
-11.6069755554199,-22.4910392761230,
-61.8430938720703,-29.4642753601074,
-68.9063491821289,-18.1124629974365,
-37.2192649841309,0.596851050853729,
-3.31900334358215,13.6510372161865,
12.3857250213623,15.4176425933838,
16.2782993316650,6.95011425018311,
23.5789184570313,2.17395353317261,
31.2168025970459,14.5354785919189,
33.4436225891113,33.0729255676270,
30.5978507995605,21.5131759643555,
25.0426406860352,-27.8027992248535,
17.1571464538574,-70.9654159545898,
19.6774044036865,-63.3538970947266,
45.6361618041992,-17.4738712310791,
79.5628128051758,8.95702934265137,
78.0433197021484,-9.98946762084961,
24.5726451873779,-34.5096969604492,
-28.8329219818115,-20.9610881805420,
-21.5716247558594,13.5987386703491,
33.4418449401856,22.7398872375488,
63.8798599243164,3.91979217529297,
23.2911014556885,-2.73679471015930,
-45.9017143249512,17.7044601440430,
-74.8349304199219,25.7234725952148,
-57.5216407775879,-8.39098739624023,
-36.7825736999512,-47.3279380798340,
-35.3086547851563,-35.8680305480957,
-30.4165458679199,20.3874435424805,
-8.64938735961914,52.7840843200684,
13.3884944915771,20.9037246704102,
17.4880638122559,-42.0224647521973,
15.3724317550659,-64.6614990234375,
21.9220981597900,-24.8371105194092,
21.8870773315430,28.9160728454590,
-1.56544172763824,42.8647003173828,
-34.6170883178711,12.9335708618164,
-45.2212448120117,-17.3736572265625,
-27.7268314361572,-10.3843021392822,
-15.5727958679199,26.1698284149170,
-28.8266124725342,46.2864532470703,
-45.6717453002930,23.9602680206299,
-38.8937492370606,-18.2485771179199,
-18.9619026184082,-37.9986190795898,
-11.9124402999878,-29.0243263244629,
-24.9209766387939,-18.6616764068604,
-37.9900398254395,-24.3662872314453,
-38.0554504394531,-26.2486228942871,
-27.7084655761719,2.11402893066406,
-20.3209629058838,45.8924827575684,
-17.0541210174561,63.3914146423340,
-16.6225452423096,45.8161010742188,
-23.9661788940430,27.3594474792480,
-39.2474555969238,29.5201930999756,
-48.2408485412598,34.3360786437988,
-35.8122673034668,8.85194969177246,
-8.36292552947998,-36.3897972106934,
21.0667495727539,-58.1472244262695,
36.6293716430664,-39.9917297363281,
30.6230411529541,-14.0678195953369,
2.89347410202026,-14.3109540939331,
-23.9468879699707,-35.1043586730957,
-21.3937835693359,-46.4233970642090,
21.2745647430420,-33.7441749572754,
65.9388961791992,-14.1802310943604,
63.9890403747559,-1.57543611526489,
13.7907314300537,10.9176540374756,
-30.1368579864502,33.7020721435547,
-26.1952972412109,57.1596450805664,
-1.72467994689941,66.7352981567383,
-8.24704933166504,54.8357658386231,
-49.5022010803223,29.9772357940674,
-73.5801696777344,5.01711225509644,
-47.7862854003906,-10.0779647827148,
4.98248100280762,-15.4282360076904,
39.3602218627930,-13.6182851791382,
45.2269668579102,-6.01139688491821,
46.2306060791016,5.90697431564331,
51.5310440063477,20.6274452209473,
50.8658981323242,29.3957424163818,
40.1727294921875,19.1770114898682,
29.8276653289795,-5.15540695190430,
21.6468772888184,-16.9822483062744,
5.35134696960449,-1.56863105297089,
-16.9578285217285,17.8425769805908,
-28.4323844909668,13.7693023681641,
-21.4707756042480,-9.21544075012207,
-7.65325546264648,-20.0904502868652,
-2.39304542541504,1.27107298374176,
-3.36304497718811,31.7773151397705,
-6.91942119598389,44.8931083679199,
-19.5813331604004,45.5288124084473,
-45.8102836608887,50.4180183410645,
-61.9545097351074,46.2397689819336,
-40.0495681762695,9.03431415557861,
0.488854408264160,-42.3914756774902,
13.0312919616699,-57.4505653381348,
-14.8808021545410,-24.5327377319336,
-37.6718177795410,1.93916130065918,
-20.5429782867432,-30.1257667541504,
14.6041631698608,-86.3872528076172,
23.3365688323975,-87.6600799560547,
-0.484818935394287,-20.3912944793701,
-24.4746589660645,38.6887969970703,
-24.0891189575195,26.6200218200684,
-8.23788833618164,-19.0404548645020,
9.01626300811768,-21.3051815032959,
27.9020843505859,23.6167812347412,
44.5461578369141,47.5347442626953,
42.4935569763184,15.5056381225586,
24.2293071746826,-30.7070693969727,
9.96435928344727,-37.0248756408691,
10.0573406219482,-14.4227981567383,
5.07850551605225,-6.25901794433594,
-9.70888519287109,-18.5922927856445,
-11.9280290603638,-23.2249259948730,
11.8398532867432,-9.96907711029053,
32.9674682617188,-4.10924339294434,
16.8527622222900,-10.9965963363647,
-17.9898567199707,-6.57914018630981,
-21.9850254058838,14.7317733764648,
13.0051355361938,27.3779201507568,
32.7800636291504,11.7606935501099,
1.04464888572693,-12.5999526977539,
-47.1687622070313,-18.4086112976074,
-57.5860824584961,-5.78607988357544,
-29.9436206817627,3.98680543899536,
-4.83694458007813,7.91718912124634,
3.84724140167236,21.7239131927490,
12.5810546875000,34.9152259826660,
30.1568126678467,22.7604560852051,
37.4196090698242,-1.43340992927551,
19.5405769348145,4.06909513473511,
-10.8508586883545,39.3898887634277,
-36.7915344238281,52.2902450561523,
-54.3183212280273,12.6895484924316,
-59.4176788330078,-40.9656867980957,
-38.9985122680664,-52.9794006347656,
1.80170929431915,-33.5481719970703,
24.2266178131104,-32.6572151184082,
4.79863309860230,-54.6564178466797,
-25.9354343414307,-46.0441398620606,
-22.5584926605225,8.51350212097168,
9.60012149810791,48.9750328063965,
26.2343235015869,25.6282482147217,
7.88414192199707,-27.2807502746582,
-13.7649965286255,-43.9419784545898,
-5.34115743637085,-22.7680530548096,
18.0602474212647,-17.1527328491211,
24.1519241333008,-41.1623725891113,
10.9272174835205,-45.4247093200684,
4.38901615142822,-1.52020359039307,
9.83945465087891,49.0534896850586,
7.80150127410889,53.1624374389648,
-8.26047325134277,20.0725326538086,
-20.7982578277588,5.47884845733643,
-18.4365139007568,25.5024223327637,
-9.07743263244629,40.9496803283691,
-2.55252456665039,22.4867382049561,
5.84694910049439,-8.58360004425049,
23.5122909545898,-18.5471534729004,
45.6201362609863,-6.66519880294800,
57.3867225646973,5.98427200317383,
56.2210121154785,5.76782560348511,
47.8649482727051,7.62392091751099,
33.6419639587402,25.4182453155518,
12.3375005722046,48.3444862365723,
-5.72208738327026,52.5836029052734,
-6.16219186782837,29.8311042785645,
3.27506732940674,-0.317181825637817,
-0.586095631122589,-13.3389749526978,
-24.7529640197754,2.65234279632568,
-44.3362426757813,30.4073352813721,
-35.2839469909668,41.5214614868164,
-5.05522966384888,27.2751750946045,
11.1721525192261,13.5374307632446,
-5.49268770217896,23.7601871490479,
-37.0256233215332,49.9639358520508,
-52.8389549255371,65.6792755126953,
-41.0780372619629,51.3089294433594,
-19.2498073577881,15.9801712036133,
-3.05192899703980,-20.7412738800049,
-0.0682814568281174,-45.8487625122070,
-4.15898799896240,-53.4215888977051,
-8.50937271118164,-35.6008224487305,
-6.86086845397949,3.74724245071411,
-2.42419934272766,35.4551124572754,
-2.93331480026245,40.5625190734863,
-9.88861846923828,32.6671905517578,
-16.8773174285889,39.7819290161133,
-16.4331607818604,56.5140342712402,
-9.79324436187744,41.0108337402344,
-1.22319173812866,-19.0672302246094,
9.56078338623047,-75.1499862670898,
27.1109542846680,-71.2443237304688,
43.3937950134277,-24.9904479980469,
39.0658798217773,-4.79500961303711,
16.2500114440918,-34.4097137451172,
-5.12844848632813,-55.5968017578125,
-9.54826164245606,-21.1321315765381,
-8.38502979278565,31.4527111053467,
-15.4046907424927,36.5467147827148,
-21.7286052703857,-9.36319160461426,
-9.36965179443359,-37.9655342102051,
13.6411905288696,-15.1301822662354,
21.3818931579590,20.4765739440918,
8.96970939636231,22.6898365020752,
4.41624832153320,3.99169397354126,
23.5477313995361,3.44101524353027,
37.2868080139160,20.2855072021484,
16.0355281829834,19.6635437011719,
-25.9243850708008,-7.12900543212891,
-46.0922927856445,-22.6297626495361,
-30.0847244262695,-13.2707586288452,
-8.80246448516846,-6.34741926193237,
-9.70321846008301,-27.8170528411865,
-22.1660785675049,-57.1140213012695,
-22.5248794555664,-55.6549606323242,
-9.78539752960205,-15.1344795227051,
-1.20083320140839,28.4503364562988,
2.37683939933777,41.8435173034668,
12.6150550842285,30.9744014739990,
25.8266448974609,20.9065799713135,
17.0419692993164,21.3395805358887,
-19.3520011901855,21.1781349182129,
-52.3521919250488,6.07763195037842,
-46.4912910461426,-25.9386749267578,
-13.0600757598877,-56.1176872253418,
9.40515041351318,-56.8932762145996,
-3.09301710128784,-26.0689640045166,
-30.2154884338379,6.26820945739746,
-40.0740699768066,8.51579189300537,
-29.6244144439697,-15.7083921432495,
-18.3298091888428,-34.3694152832031,
-17.6682052612305,-26.1397590637207,
-16.9734096527100,-0.171982884407043,
-9.19019031524658,14.9442958831787,
0.944813609123230,13.4882221221924,
7.82246017456055,6.80719280242920,
12.6181659698486,-4.23495435714722,
23.3141517639160,-18.5688743591309,
41.3952255249023,-23.2924823760986,
59.5381355285645,-5.20645284652710,
65.3138275146484,21.4786224365234,
59.3166618347168,26.0709590911865,
47.4969253540039,6.67205905914307,
37.9963378906250,1.09511744976044,
31.9096698760986,25.3131618499756,
15.6694002151489,44.5196266174316,
-18.6671791076660,14.8074779510498,
-46.3972091674805,-40.5528907775879,
-38.1282081604004,-55.8366661071777,
-3.59715938568115,-12.1569881439209,
10.8728780746460,26.5796298980713,
-17.7485637664795,9.94026184082031,
-49.9447326660156,-32.9963302612305,
-37.1095008850098,-39.5810012817383,
6.67492818832398,-2.39619588851929,
10.8582601547241,31.0889816284180,
-44.4132461547852,31.9333839416504,
-86.9224853515625,19.0690841674805,
-51.1635665893555,11.1475744247437,
25.5981445312500,-1.24204695224762,
49.6163635253906,-30.1264572143555,
2.47833299636841,-52.9382400512695,
-41.2272491455078,-49.5301742553711,
-19.1857395172119,-37.3704299926758,
33.2219848632813,-47.3838577270508,
51.9483947753906,-69.3261947631836,
38.8036346435547,-64.7091140747070,
36.0535697937012,-29.4024772644043,
44.6656799316406,11.3786716461182,
21.5763759613037,35.9344329833984,
-35.4370994567871,40.5881080627441,
-60.9396820068359,30.2485828399658,
-16.5566291809082,7.89271879196167,
43.9163475036621,-12.2783098220825,
47.8385009765625,-3.88450980186462,
2.44039297103882,30.5786590576172,
-25.5014991760254,50.1579208374023,
-1.68739390373230,36.4657592773438,
41.5500259399414,15.5996608734131,
53.8832015991211,14.4573678970337,
32.3119392395020,8.06958866119385,
5.76833534240723,-31.1433029174805,
-9.79696369171143,-74.0643997192383,
-9.80298519134522,-59.1448097229004,
6.87841892242432,7.60212421417236,
16.8873195648193,53.2524337768555,
-5.72096061706543,29.3747806549072,
-47.0359611511231,-20.9757156372070,
-56.4925003051758,-23.8845958709717,
-16.6378517150879,19.4059448242188,
16.6597175598145,43.4979362487793,
-12.1461048126221,14.1608419418335,
-70.1754455566406,-35.8730506896973,
-72.0174255371094,-57.6247253417969,
-1.88569331169128,-45.7673606872559,
49.7483673095703,-19.6919898986816,
17.3438320159912,-3.09080648422241,
-44.1342353820801,-4.64341974258423,
-42.5689392089844,-21.2925491333008,
20.4923572540283,-32.1948051452637,
52.6419944763184,-14.0968484878540,
8.81837654113770,21.4856395721436,
-45.7458801269531,35.5489501953125,
-36.5441780090332,4.65263319015503,
16.4116592407227,-33.8240318298340,
38.5258827209473,-25.0881462097168,
6.39772415161133,27.9965591430664,
-30.6959037780762,65.3363647460938,
-27.6088447570801,54.9189300537109,
-3.58159255981445,31.1863498687744,
-4.07750272750855,36.1229553222656,
-26.9329319000244,62.3794708251953,
-32.7625427246094,67.2431335449219,
-6.25437164306641,36.8265762329102,
27.2936687469482,6.84878969192505,
28.1799240112305,0.739365458488464,
-6.26213932037354,0.699660181999207,
-30.6168632507324,-17.1917304992676,
-12.7907629013062,-46.7801284790039,
24.6739387512207,-60.6039581298828,
33.0265922546387,-52.0538139343262,
-2.09911847114563,-40.0170745849609,
-41.5021858215332,-30.5746021270752,
-43.8873176574707,-12.8721837997437,
-21.1448535919189,8.89403915405273,
-19.9238357543945,11.3236293792725,
-52.9102401733398,-15.6041040420532,
-74.4182586669922,-43.0356979370117,
-47.0069999694824,-27.6551704406738,
6.38090085983276,26.4923763275147,
28.4418144226074,64.8474197387695,
-0.119949340820313,48.5077056884766,
-42.2377624511719,-3.98361420631409,
-53.2436943054199,-37.4665756225586,
-29.2228679656982,-25.2793922424316,
3.37877035140991,9.76972675323486,
26.6913337707520,28.6903438568115,
38.8680305480957,19.8664779663086,
46.0262947082520,5.73631858825684,
51.4215545654297,6.65072441101074,
53.1273040771484,20.7165966033936,
48.5160789489746,29.1045875549316,
39.0326805114746,20.3065452575684,
26.5423221588135,1.94025957584381,
17.2324390411377,-2.73889636993408,
14.7255458831787,14.0347728729248,
15.4401092529297,37.5318069458008,
11.3085689544678,43.6096572875977,
4.23805570602417,30.5861549377441,
-2.59340667724609,17.4104709625244,
-12.1508159637451,16.5443649291992,
-24.3137550354004,21.2892074584961,
-31.6849689483643,16.5716533660889,
-24.2834014892578,11.7355327606201,
-7.72975254058838,23.6698951721191,
-0.488936722278595,44.3783264160156,
-8.07710456848145,46.5996742248535,
-19.3985538482666,21.9024200439453,
-19.2117652893066,1.84651553630829,
-14.5181941986084,16.3769989013672,
-17.4038887023926,53.3797225952148,
-25.1412887573242,68.3571395874023,
-22.6332244873047,44.6762886047363,
-9.50980472564697,11.5825462341309,
0.399491518735886,-3.04003906250000,
-1.63065969944000,-7.25309514999390,
-3.83423948287964,-22.4215488433838,
4.14584779739380,-46.5295982360840,
12.4870567321777,-51.6861763000488,
7.47592449188232,-27.3412628173828,
-2.64888262748718,1.46335089206696,
2.16985797882080,11.8057317733765,
19.4036731719971,9.03308391571045,
21.3144073486328,12.7621049880981,
-4.62663316726685,21.9072360992432,
-32.4470901489258,20.1766281127930,
-25.1807956695557,-0.409903168678284,
11.3438434600830,-20.4085941314697,
33.8892173767090,-11.1551160812378,
13.5247392654419,23.6284065246582,
-22.9933052062988,44.3689918518066,
-31.9056568145752,22.3997650146484,
-8.53048133850098,-27.3338203430176,
12.7721920013428,-54.3325271606445,
12.2329759597778,-29.9190597534180,
8.19566345214844,15.6156101226807,
21.2145996093750,29.5239353179932,
36.7374916076660,8.99272537231445,
25.1684856414795,-5.55955076217651,
-8.40858268737793,8.58636856079102,
-29.4541835784912,19.5234546661377,
-25.9132213592529,-8.59091949462891,
-20.7831516265869,-52.6800308227539,
-27.6598930358887,-58.0900764465332,
-26.1589775085449,-15.8185253143311,
-1.59879517555237,24.5191802978516,
20.7819709777832,20.0247344970703,
8.41985797882080,-5.92029571533203,
-20.3765125274658,-8.34868812561035,
-21.6109600067139,14.9806022644043,
7.30171203613281,27.4779434204102,
20.3490886688232,8.35667324066162,
-7.00529813766480,-21.1605377197266,
-37.9813117980957,-35.0633773803711,
-29.1032104492188,-30.2358570098877,
2.99532461166382,-17.0687580108643,
10.3400688171387,-1.43426239490509,
-10.1705760955811,7.35037326812744,
-16.2739562988281,-4.13025808334351,
12.2342567443848,-35.2939605712891,
43.3419494628906,-58.9850082397461,
35.9229621887207,-47.9516601562500,
0.365180730819702,-5.65348625183106,
-25.5368061065674,29.4934062957764,
-24.4932289123535,35.4177780151367,
-12.0920486450195,23.3531684875488,
-8.29292869567871,9.68818473815918,
-12.8642196655273,-2.57891464233398,
-16.9949226379395,-19.1216583251953,
-23.7015819549561,-33.6899452209473,
-30.6183128356934,-36.1415367126465,
-27.7025108337402,-30.2059898376465,
-9.89517116546631,-26.6752452850342,
12.6656122207642,-24.0175533294678,
18.1448898315430,-14.3431539535522,
-6.03827667236328,-4.43017244338989,
-43.0659751892090,-12.9258480072021,
-55.2895240783691,-40.6444129943848,
-24.7751197814941,-57.2731590270996,
23.0027122497559,-33.7499618530273,
44.0112190246582,7.45072937011719,
20.2028121948242,20.8028507232666,
-14.7098321914673,-10.7609195709229,
-12.9907493591309,-51.2272911071777,
27.9107284545898,-53.7938652038574,
59.9561538696289,-13.3941888809204,
45.2646903991699,30.7521400451660,
5.75986671447754,41.8318214416504,
-10.9517393112183,21.5169372558594,
4.66421413421631,-0.0274784564971924,
18.8531341552734,0.124125450849533,
5.05318593978882,16.4084682464600,
-20.4958000183105,22.6979846954346,
-22.4158554077148,1.67453765869141,
-1.54209661483765,-32.6261482238770,
13.4682903289795,-47.9075393676758,
11.1893053054810,-30.0809364318848,
6.12053966522217,1.76535797119141,
4.71460247039795,23.8674812316895,
-5.70015716552734,33.0489578247070,
-26.4746856689453,38.4814300537109,
-31.6967029571533,39.9019699096680,
-3.82090520858765,26.5452709197998,
27.6356906890869,-0.639247238636017,
21.0137958526611,-10.6556987762451,
-11.0549173355103,9.73552227020264,
-21.9527568817139,34.8410987854004,
11.1909456253052,33.5946273803711,
49.6262512207031,11.8021621704102,
53.3132553100586,1.74529433250427,
37.3523330688477,14.3021221160889,
36.6056213378906,27.8355293273926,
44.3521461486816,28.2005825042725,
28.3170852661133,27.5790863037109,
-9.77346229553223,31.9518756866455,
-31.8974628448486,24.0996894836426,
-15.9992456436157,-4.54554128646851,
16.3531856536865,-23.1351776123047,
30.5160121917725,4.08602237701416,
19.7110881805420,55.9177436828613,
-6.90012645721436,70.5205383300781,
-46.5602569580078,25.9518508911133,
-82.9735870361328,-26.2346992492676,
-83.5594482421875,-36.1529922485352,
-35.9492378234863,-10.9462852478027,
17.7809543609619,7.18575763702393,
24.9836673736572,-0.140794098377228,
-0.973757982254028,-9.32205390930176,
-8.81792736053467,-0.964608728885651,
15.6496114730835,15.4640140533447,
27.2062320709229,24.4003829956055,
-3.30285167694092,26.9299831390381,
-40.5245933532715,22.9007034301758,
-34.2161521911621,14.0373668670654,
5.21696996688843,9.15069389343262,
18.0770263671875,23.6968345642090,
-18.0606918334961,42.2444267272949,
-60.7742919921875,26.5688037872314,
-66.7628326416016,-31.8639030456543,
-37.0214805603027,-78.2225646972656,
3.92373585700989,-61.6137847900391,
38.5177230834961,3.86083698272705,
53.7765655517578,44.0223083496094,
40.4093475341797,20.9935512542725,
6.70099067687988,-20.5181179046631,
-19.6157913208008,-19.9724159240723,
-19.1229496002197,20.7752532958984,
-10.6609745025635,53.0886192321777,
-21.2333469390869,51.2382278442383,
-48.5973548889160,25.0219459533691,
-62.7259216308594,-6.46568489074707,
-52.7377853393555,-36.1503219604492,
-39.7439956665039,-53.7487335205078,
-32.8018951416016,-49.5125427246094,
-15.6437454223633,-33.2841110229492,
14.8709678649902,-36.2946052551270,
29.6018218994141,-59.6239624023438,
12.4797334671021,-62.2842559814453,
-17.9004993438721,-22.7599716186523,
-24.7065620422363,22.9918460845947,
-3.60828685760498,20.4415626525879,
21.8908252716064,-11.8722877502441,
36.9422836303711,-13.4114809036255,
45.1088752746582,28.6742115020752,
43.2911071777344,58.0160255432129,
21.5343780517578,34.3080368041992,
-6.79273891448975,-9.07282161712647,
-8.35588264465332,-12.7778549194336,
23.4870052337647,13.2116861343384,
47.1494483947754,14.1711177825928,
35.4340820312500,-20.4514217376709,
11.4392566680908,-39.9992675781250,
17.1734218597412,-10.8173894882202,
47.3601722717285,33.5038833618164,
56.8163948059082,50.4050292968750,
24.4297962188721,40.5415725708008,
-17.2504711151123,37.0487174987793,
-28.7035007476807,41.1318550109863,
-11.3615236282349,32.9336280822754,
7.01686286926270,10.7934761047363,
14.7207841873169,2.21374034881592,
17.0888614654541,18.4673614501953,
14.3589611053467,38.0613174438477,
-0.485998988151550,35.3892440795898,
-21.2158145904541,14.0540304183960,
-30.9533252716064,-7.23192405700684,
-23.8157691955566,-25.8721218109131,
-15.2625246047974,-45.0977134704590,
-15.0837726593018,-52.7831764221191,
-17.2616004943848,-27.6208248138428,
-6.20659255981445,20.9284019470215,
13.5385398864746,57.4225311279297,
26.6341228485107,51.6208190917969,
23.4035968780518,14.3202552795410,
15.7740783691406,-7.61951684951782,
8.61153697967529,11.9025077819824,
-3.97963237762451,44.7402076721191,
-23.3240013122559,43.8512039184570,
-36.3063316345215,-0.358541488647461,
-25.8942375183105,-45.7848930358887,
3.75366020202637,-50.9526634216309,
31.6904430389404,-24.7825698852539,
43.0786781311035,-15.2979240417480,
44.4698524475098,-35.1895523071289,
45.2702713012695,-43.7368583679199,
39.9042930603027,-6.96321105957031,
19.5302314758301,49.0849266052246,
-11.2309284210205,60.7167091369629,
-36.8781280517578,16.8054733276367,
-49.3335380554199,-27.6930637359619,
-46.9953079223633,-19.1077289581299,
-32.2104682922363,29.2220859527588,
-7.42532920837402,57.2342681884766,
14.8341674804688,36.5182685852051,
18.3204040527344,-0.753198862075806,
8.44391632080078,-10.8894386291504,
4.12097787857056,11.6587104797363,
17.9593677520752,34.6109619140625,
32.5359458923340,32.0671043395996,
29.5934658050537,6.92969465255737,
18.2665252685547,-24.0627822875977,
13.9512472152710,-40.6197509765625,
16.9686183929443,-34.9896583557129,
10.1739473342896,-12.4548835754395,
-0.794891834259033,9.80329799652100,
4.02802705764771,17.3049049377441,
33.2977561950684,17.5659523010254,
60.9765739440918,21.5907974243164,
54.7661399841309,27.7465190887451,
18.4719886779785,18.8301486968994,
-24.1115550994873,-6.59633636474609,
-54.0125122070313,-18.5527534484863,
-64.2136077880859,7.23456382751465,
-48.7474555969238,44.6558151245117,
-11.0240554809570,43.9409980773926,
24.1712703704834,-3.23338174819946,
36.2185821533203,-48.1626396179199,
35.7265357971191,-39.5785408020020,
45.3181304931641,12.1584167480469,
55.4581909179688,51.2904319763184,
33.6795806884766,50.0890007019043,
-21.6685676574707,23.7584724426270,
-61.0404815673828,1.41911017894745,
-40.3187713623047,-14.1141796112061,
14.2939233779907,-24.4880180358887,
40.9188728332520,-22.2076416015625,
20.8005523681641,-4.11860942840576,
-7.05614376068115,11.4414100646973,
-16.7567920684814,8.43091773986816,
-18.4048080444336,-3.59878134727478,
-28.0020446777344,-1.93017256259918,
-32.5721359252930,14.7606964111328,
-25.6791496276855,20.5856723785400,
-29.4440383911133,-1.00298118591309,
-55.0538177490234,-35.3733825683594,
-71.2365646362305,-57.4506492614746,
-36.2064399719238,-62.5198097229004,
33.1057624816895,-48.4220886230469,
73.1366424560547,-10.8456850051880,
51.0292129516602,36.0059318542481,
5.72398185729981,60.9349555969238,
-12.9731454849243,48.7951316833496,
-7.55984258651733,26.9171867370605,
-6.23814201354981,32.5227928161621,
-17.4686679840088,56.6290016174316,
-26.5334815979004,51.2994117736816,
-22.1006507873535,1.35004556179047,
-4.67052459716797,-43.6981773376465,
18.2014980316162,-40.4953460693359,
34.7797470092773,-13.6518545150757,
30.0779571533203,-13.4980182647705,
-1.43300652503967,-40.6115760803223,
-31.3972396850586,-50.1569175720215,
-25.3952999114990,-26.8759899139404,
11.7877607345581,-3.32328796386719,
34.4332885742188,-6.30938863754273,
23.7357311248779,-10.0532617568970,
9.37120437622070,8.55356121063232,
13.2408475875855,23.9460945129395,
18.5769996643066,1.28485536575317,
8.34595870971680,-38.9554901123047,
1.56251740455627,-36.1704711914063,
25.0384235382080,14.4451227188110,
58.1937332153320,47.8719978332520,
49.8408966064453,19.2370357513428,
-1.82580602169037,-31.1671810150147,
-35.1253051757813,-46.4969978332520,
-13.1224431991577,-19.8358325958252,
24.8849411010742,5.13922595977783,
20.3774185180664,2.73623609542847,
-15.3214435577393,-11.9825458526611,
-30.2427406311035,-18.9625320434570,
-10.3403730392456,-24.0783081054688,
13.8563976287842,-30.4515724182129,
26.4966106414795,-31.3267288208008,
41.4749908447266,-25.0130252838135,
62.5590019226074,-19.5680408477783,
56.3403244018555,-13.5502223968506,
6.97689580917358,5.95961380004883,
-41.7376785278320,28.7234020233154,
-40.7695693969727,18.1631870269775,
-7.18864059448242,-29.8752651214600,
9.78746700286865,-67.3923110961914,
6.78702974319458,-51.6659507751465,
20.2252635955811,3.75105977058411,
54.1648635864258,35.2334785461426,
61.8469772338867,10.2748661041260,
25.1903915405273,-36.2494392395020,
-11.4270982742310,-55.6533241271973,
-3.39326667785645,-37.0675544738770,
23.0742683410645,-5.42497444152832,
13.9750852584839,12.7656383514404,
-23.8609580993652,5.43817949295044,
-28.4582099914551,-18.9261035919189,
12.7474803924561,-29.0643157958984,
41.7239189147949,-1.59075164794922,
11.4229345321655,41.0931015014648,
-36.5225296020508,43.9824905395508,
-35.9683990478516,-15.2809286117554,
10.8959102630615,-80.8368835449219,
53.7069358825684,-77.5645751953125,
58.7889785766602,-6.44994020462036,
43.5955657958984,52.8694877624512,
33.1178054809570,50.6697807312012,
31.0598297119141,22.1745853424072,
27.5901927947998,23.1488609313965,
29.9122333526611,43.0155029296875,
39.2800292968750,42.9216194152832,
38.8898353576660,26.4699077606201,
16.9682674407959,36.3174743652344,
-12.9356575012207,70.9731063842773,
-34.6711311340332,71.2331390380859,
-45.3777389526367,6.05743646621704,
-35.8490943908691,-59.5177345275879,
6.56549167633057,-51.9336166381836,
60.8020935058594,7.82144260406494,
82.2697296142578,35.9923057556152,
50.3008422851563,-1.46446037292480,
3.00948286056519,-50.4180374145508,
2.08929371833801,-60.8005867004395,
40.4821739196777,-49.9608688354492,
57.2649879455566,-49.0793876647949,
27.5676078796387,-47.3349685668945,
-0.727801144123077,-19.5385131835938,
8.81616973876953,10.6987905502319,
29.7337131500244,1.70414698123932,
24.0907211303711,-38.6587257385254,
10.3804626464844,-47.9210662841797,
24.9692173004150,2.01690530776978,
45.9701080322266,59.8355636596680,
15.0378408432007,58.7911033630371,
-62.2084045410156,6.75169754028320,
-95.1466369628906,-35.6902885437012,
-33.6304397583008,-33.3260574340820,
53.4039993286133,-0.896636009216309,
67.9565200805664,21.6090068817139,
9.70083045959473,13.0836219787598,
-25.5765209197998,-8.44625568389893,
7.39606237411499,-13.4289855957031,
45.7981567382813,10.7600908279419,
24.9309616088867,40.5735321044922,
-30.6582965850830,36.3270263671875,
-49.2144737243652,-10.9920959472656,
-16.8163642883301,-53.8685417175293,
11.5193910598755,-39.2770690917969,
-6.58017539978027,19.0033550262451,
-40.8050270080566,53.4401321411133,
-39.1594047546387,37.1554107666016,
-2.13049173355103,10.4789342880249,
22.1530246734619,16.4713745117188,
2.48039245605469,34.6236648559570,
-36.8684577941895,16.4200267791748,
-52.5310554504395,-31.6763153076172,
-24.5468215942383,-47.2688255310059,
18.2194995880127,-4.28030014038086,
27.8046340942383,42.4024353027344,
0.425946831703186,36.2055625915527,
-22.1368236541748,-3.60260486602783,
-7.64766979217529,-14.5118036270142,
26.9229946136475,14.0449790954590,
36.7585105895996,29.2664413452148,
12.1115798950195,1.44338226318359,
-5.40699243545532,-30.5720825195313,
15.8512773513794,-17.6684017181397,
49.9012069702148,30.1434326171875,
48.7159957885742,62.8833732604981,
19.1332397460938,52.9353599548340,
4.91827487945557,22.8530426025391,
19.6722946166992,-0.372480332851410,
27.8496646881104,-14.9276819229126,
2.30559897422791,-25.4866924285889,
-32.0784492492676,-26.6314525604248,
-31.7933883666992,-20.4950962066650,
-3.19335246086121,-20.1279716491699,
16.0737075805664,-24.4395160675049,
14.6884584426880,-20.7634868621826,
17.6061325073242,0.512983202934265,
29.2035827636719,28.2342700958252,
15.4901075363159,43.5884590148926,
-35.2183570861816,39.8427085876465,
-73.0587234497070,18.5813484191895,
-49.4647636413574,-18.4333820343018,
9.97125911712647,-57.3770523071289,
32.8487472534180,-64.0701904296875,
1.95587325096130,-20.7468986511230,
-25.6385459899902,32.0016708374023,
-5.40089988708496,37.2034721374512,
31.9121646881104,-8.63786888122559,
34.0883026123047,-45.0760040283203,
7.87781524658203,-25.6756973266602,
1.77899050712585,25.0894393920898,
24.1806182861328,47.0604171752930,
29.9205627441406,22.7053642272949,
-3.97715735435486,-13.5221691131592,
-38.0790252685547,-25.2646522521973,
-25.3122272491455,-14.1851596832275,
19.9671478271484,-5.44500350952148,
48.5791435241699,-9.25780677795410,
43.5465393066406,-22.8715496063232,
32.3775901794434,-34.5573577880859,
41.8081665039063,-36.3071517944336,
54.2949562072754,-25.0693225860596,
42.0284271240234,-6.30636453628540,
12.9132823944092,3.89129328727722,
-1.94672703742981,-1.08133900165558,
9.72838020324707,-13.5182409286499,
27.3609580993652,-23.0464286804199,
24.7681503295898,-25.7278995513916,
3.05308938026428,-21.2197761535645,
-12.8374061584473,-12.1522350311279,
-4.06570291519165,3.66772508621216,
17.4466361999512,20.0331153869629,
25.4532737731934,29.4764213562012,
13.6740217208862,33.9446029663086,
-4.59444379806519,38.8805885314941,
-16.0969696044922,40.3503227233887,
-23.4735660552979,26.3535633087158,
-37.5514106750488,-2.31414747238159,
-55.2094306945801,-27.7964458465576,
-58.7090263366699,-26.7678413391113,
-39.7205276489258,-5.36064243316650,
-12.7498292922974,11.9546318054199,
7.11928176879883,11.9602203369141,
18.7744159698486,8.76781082153320,
28.2451438903809,20.3475074768066,
29.3092765808105,40.5774345397949,
11.7339916229248,42.3378334045410,
-17.9276561737061,19.0785598754883,
-32.9040145874023,-3.19286870956421,
-19.2197704315186,-0.174564719200134,
2.47038698196411,15.2247934341431,
-4.11835813522339,9.98769092559815,
-41.1075363159180,-23.1818637847900,
-69.1964263916016,-52.0415153503418,
-57.3988990783691,-43.0157089233398,
-19.7640991210938,-1.05722117424011,
8.75716400146484,29.9680423736572,
11.1951236724854,21.9445552825928,
4.27292871475220,-5.13675498962402,
-0.0179711580276489,-12.0642623901367,
-7.02999353408814,11.0394964218140,
-17.7567749023438,34.9588394165039,
-13.8033351898193,30.7327327728272,
4.81945991516113,7.95799446105957,
8.41749000549316,-1.37792003154755,
-24.2735767364502,4.67816114425659,
-58.9290809631348,-3.25569868087769,
-45.5636024475098,-35.4208641052246,
7.01761722564697,-53.8200378417969,
37.4686470031738,-29.1311187744141,
16.7567481994629,16.8616828918457,
-8.11503601074219,31.8244953155518,
7.45564746856689,4.97183465957642,
40.2265014648438,-20.6238689422607,
28.1839561462402,-14.6053962707520,
-23.0274353027344,0.504255890846252,
-43.1723518371582,-3.31949949264526,
-2.02637457847595,-14.5779905319214,
51.1456031799316,-5.90996646881104,
62.1749534606934,13.8051128387451,
44.5505218505859,11.2037029266357,
39.9906616210938,-11.0408267974854,
44.0473518371582,-6.69519138336182,
26.2691116333008,38.2209129333496,
-8.44963932037354,82.1898956298828,
-25.9365844726563,80.3605422973633,
-19.3109645843506,44.9030876159668,
-26.1480598449707,22.1422176361084,
-54.3522148132324,30.4422702789307,
-56.0672836303711,44.3962326049805,
-0.451127648353577,36.2152748107910,
63.6252822875977,12.4570846557617,
67.5528869628906,-6.47479534149170,
12.1677083969116,-11.7260780334473,
-37.3451995849609,-2.84318447113037,
-39.0358963012695,13.9388027191162,
-9.42632484436035,18.8798885345459,
15.5120296478271,-5.22940826416016,
25.1850528717041,-42.9773330688477,
25.9604816436768,-58.2850494384766,
11.5771665573120,-34.6383590698242,
-21.3444442749023,2.59238934516907,
-49.1667213439941,21.9182605743408,
-49.0657730102539,20.1425704956055,
-34.6552009582520,21.1586399078369,
-32.0307769775391,28.9990043640137,
-42.4348602294922,28.2219257354736,
-38.7073554992676,18.1856899261475,
-12.3055305480957,17.5074710845947,
18.1011238098145,26.5019664764404,
31.2588787078857,21.4539108276367,
29.5730876922607,-7.27116966247559,
25.3556232452393,-31.1686477661133,
17.2393722534180,-13.8088932037354,
-0.227819800376892,31.7885704040527,
-15.1435108184814,55.5023689270020,
-7.96608352661133,37.4890213012695,
12.4774179458618,8.64291381835938,
16.2017612457275,2.21503782272339,
-8.13126373291016,10.8739852905273,
-33.3526458740234,1.94462251663208,
-30.8729057312012,-28.1688632965088,
-8.25003814697266,-46.7015075683594,
-3.16206526756287,-31.3135375976563,
-28.0388374328613,-4.37808609008789,
-53.8739318847656,3.86325287818909,
-38.8623580932617,-1.95392525196075,
13.3233127593994,9.16036033630371,
54.1500968933106,42.8535041809082,
44.9696388244629,61.6304969787598,
-6.15710735321045,31.9574203491211,
-51.1916580200195,-19.6213493347168,
-57.2876167297363,-36.6592330932617,
-34.0565452575684,-1.67589688301086,
-8.89466667175293,37.8632392883301,
3.74529123306274,32.0669479370117,
12.2637662887573,-7.30135202407837,
16.6282997131348,-29.0092582702637,
6.17039632797241,-8.37007045745850,
-19.2616157531738,23.1278495788574,
-39.3666419982910,21.7975311279297,
-34.6068115234375,-11.7467432022095,
-11.4334230422974,-39.4454727172852,
0.377161055803299,-35.1009902954102,
-16.9609737396240,-11.3084821701050,
-44.3690986633301,1.44982719421387,
-53.7273025512695,-12.9520778656006,
-34.4437522888184,-45.7309455871582,
2.09117650985718,-68.6513900756836,
31.6818714141846,-59.4391098022461,
45.6992645263672,-13.7938480377197,
48.4944458007813,43.4553146362305,
43.8018035888672,70.7269821166992,
32.4866104125977,46.5917778015137,
16.7144432067871,1.98124790191650,
9.09636592864990,-15.5220775604248,
20.1713008880615,10.6510162353516,
41.1406822204590,41.9174003601074,
44.1104202270508,34.4393348693848,
12.1563634872437,-3.58525943756104,
-30.7398681640625,-24.0711250305176,
-48.2433166503906,-4.59635925292969,
-29.8921127319336,25.1787319183350,
-6.40454292297363,25.4276638031006,
-10.3942871093750,2.54433059692383,
-39.8458480834961,-8.25283527374268,
-57.7202682495117,5.17253780364990,
-45.0657119750977,9.56806182861328,
-16.2012348175049,-16.3162841796875,
3.14204597473145,-54.7154045104981,
2.55914878845215,-65.9486160278320,
0.644063115119934,-41.8315544128418,
9.95527839660645,-16.3433170318604,
18.7459545135498,-12.2579898834229,
4.75444364547730,-17.0097885131836,
-30.1011371612549,-9.26966094970703,
-51.8430709838867,9.89588451385498,
-36.4411773681641,16.7629623413086,
-1.59344291687012,2.87933135032654,
17.5367908477783,-7.26466131210327,
14.1919574737549,5.29126548767090,
17.0963001251221,29.3518238067627,
41.1670951843262,42.3271484375000,
59.1397018432617,41.3587150573731,
36.7994956970215,42.7096405029297,
-13.4539299011230,42.2704849243164,
-48.7771873474121,17.8188076019287,
-50.1522521972656,-31.9079132080078,
-34.1208724975586,-61.9480209350586,
-16.9595642089844,-36.4931564331055,
-3.56183910369873,20.2507972717285,
-0.117945656180382,43.6943359375000,
-16.1491317749023,9.98167705535889,
-37.5600051879883,-39.8649444580078,
-29.4642353057861,-58.4330291748047,
12.6473989486694,-42.6344985961914,
47.0374984741211,-17.0339145660400,
36.0281562805176,13.0306148529053,
5.08065319061279,48.5486259460449,
1.53293514251709,66.8986511230469,
20.2685775756836,42.8896636962891,
8.90736770629883,-10.0521240234375,
-41.3013572692871,-47.4027824401856,
-68.0882263183594,-46.7737197875977,
-30.8978385925293,-31.4983501434326,
30.0813827514648,-27.6698417663574,
46.8898200988770,-29.6313953399658,
13.8046131134033,-16.4247283935547,
-13.9770021438599,4.94839525222778,
-3.41621613502502,16.5853862762451,
16.1048469543457,25.0604953765869,
8.05705070495606,39.3096046447754,
-25.2431144714355,41.6317329406738,
-53.9838523864746,13.5644378662109,
-62.8967590332031,-32.8248481750488,
-51.1931762695313,-55.3555068969727,
-16.2545127868652,-36.2898712158203,
26.4748401641846,-5.61591482162476,
40.9930686950684,12.4614572525024,
13.4767742156982,23.5636749267578,
-25.4181213378906,38.2219696044922,
-36.8325157165527,31.6527118682861,
-21.6999874114990,-18.7774353027344,
-10.6327123641968,-69.2530059814453,
-18.7549571990967,-57.2560310363770,
-26.3301982879639,8.47141647338867,
-21.4061412811279,47.1746635437012,
-20.9941139221191,12.7989082336426,
-26.9519844055176,-45.4020423889160,
-18.5385837554932,-52.1690521240234,
8.08719539642334,-3.81536722183228,
15.6218347549438,40.1393165588379,
-15.8777256011963,47.2495651245117,
-47.7024650573731,38.4715423583984,
-27.1044254302979,34.3441047668457,
28.1973571777344,21.3250007629395,
46.3889160156250,-1.11715257167816,
5.30890178680420,-4.02092027664185,
-37.5027618408203,23.0223960876465,
-26.0893821716309,44.3507156372070,
15.4481115341187,27.8442802429199,
18.0036888122559,-1.83796906471252,
-28.7359695434570,-0.440991133451462,
-69.0890731811523,18.9201583862305,
-67.5535430908203,7.87457418441773,
-42.1369476318359,-41.6334915161133,
-22.9323921203613,-76.5391540527344,
-10.8605813980103,-55.4537086486816,
9.14845275878906,-9.87023925781250,
33.5182342529297,7.12301063537598,
45.0325279235840,-0.523872613906860,
36.9171791076660,3.56125855445862,
16.1256885528564,27.6860160827637,
-4.30300426483154,39.0317077636719,
-12.6720161437988,19.5259723663330,
2.23178434371948,-4.68538808822632,
35.2398452758789,-0.931720733642578,
46.5989227294922,28.3206100463867,
9.42510890960693,48.5360717773438,
-46.0743942260742,34.0930290222168,
-55.1665306091309,-5.80507373809814,
-5.58408498764038,-41.5127067565918,
50.4409561157227,-41.7420387268066,
55.1580390930176,-0.290122747421265,
20.9310359954834,55.2073211669922,
-2.40812492370605,72.2911300659180,
-0.920602679252625,39.2305755615234,
-5.19826602935791,-7.88701820373535,
-33.8073348999023,-24.1502532958984,
-56.2361640930176,-5.28633880615234,
-44.3649101257324,16.4429721832275,
-17.3069076538086,22.7410469055176,
-15.2153053283691,25.0035552978516,
-42.5183753967285,34.6486663818359,
-65.0927200317383,38.4779777526856,
-60.8546981811523,18.6882152557373,
-42.0026283264160,-12.1566104888916,
-31.7063617706299,-28.6668148040772,
-32.4313087463379,-31.4396476745605,
-29.7078781127930,-41.9195289611816,
-13.5988569259644,-63.7866096496582,
9.71500396728516,-72.0176544189453,
31.4722518920898,-47.3289833068848,
36.5423088073731,-5.72928905487061,
14.0707092285156,24.0164566040039,
-17.9742317199707,26.1143169403076,
-27.1084384918213,11.8540563583374,
-1.15614497661591,-1.04263210296631,
27.4809761047363,-0.874522328376770,
27.7522563934326,15.8629360198975,
11.4804801940918,39.8802833557129,
16.2415313720703,50.1682167053223,
44.8537902832031,33.5299797058106,
54.8271789550781,10.2021913528442,
20.1909465789795,12.0135965347290,
-18.8370609283447,36.8271980285645,
-14.1493215560913,50.4891319274902,
18.5357761383057,32.2172431945801,
22.4687385559082,2.71884393692017,
-21.4857540130615,-6.41111564636231,
-67.8607406616211,11.0382499694824,
-69.3816223144531,27.7567825317383,
-36.3737335205078,27.2711982727051,
-8.52226638793945,18.7346553802490,
-2.05323696136475,8.92088699340820,
-5.96367216110230,0.997044801712036,
-13.0262775421143,4.78878307342529,
-26.0882644653320,31.2236480712891,
-38.4603576660156,66.1641082763672,
-30.4737968444824,71.1725082397461,
-4.78946495056152,30.4023838043213,
8.98027896881104,-14.1497659683228,
-4.93549489974976,-14.1109333038330,
-25.9615402221680,20.8401145935059,
-28.3684043884277,33.2697219848633,
-13.7059555053711,-2.72322893142700,
-0.671641945838928,-42.4312362670898,
0.0777193605899811,-27.6532154083252,
-3.97389054298401,30.4102439880371,
0.323375880718231,65.5762100219727,
7.18884372711182,40.8359069824219,
14.0936794281006,-9.82412815093994,
17.1373863220215,-26.7376651763916,
9.19715499877930,4.46025276184082,
-12.4535150527954,44.9430694580078,
-27.0241889953613,50.8531341552734,
-12.0868101119995,21.7309513092041,
28.3930549621582,-8.67516040802002,
52.4028434753418,-10.6327304840088,
35.0134811401367,9.51937389373779,
2.53417110443115,21.0837535858154,
-3.66791415214539,7.85296058654785,
15.4842996597290,-18.4562492370605,
15.7747840881348,-30.4216327667236,
-23.7024631500244,-22.2102661132813,
-67.5151901245117,-14.0877008438110,
-66.3639602661133,-17.1165237426758,
-27.9775905609131,-17.8103981018066,
-4.83759880065918,-2.50170946121216,
-24.1059207916260,19.1319923400879,
-55.0889282226563,21.8932533264160,
-50.2299194335938,0.217313885688782,
-2.67796611785889,-19.3068332672119,
44.7099227905273,-10.6845617294312,
49.6542015075684,20.5561218261719,
12.9317407608032,49.6050262451172,
-25.4970149993897,58.7619056701660,
-31.6224803924561,50.0555076599121,
-9.55963706970215,33.9406967163086,
4.96602773666382,16.8669071197510,
-15.4553737640381,4.24041652679443,
-51.4870567321777,-3.65640044212341,
-56.8220062255859,-10.2405242919922,
-18.8213214874268,-17.6590709686279,
18.9753341674805,-20.8255004882813,
12.2011699676514,-15.3516893386841,
-30.8339233398438,-5.72752952575684,
-57.0291976928711,-5.49683856964111,
-44.3062400817871,-15.0867738723755,
-22.4469070434570,-19.9663829803467,
-26.8129901885986,-9.12399482727051,
-37.5536766052246,7.30748319625855,
-13.9724102020264,8.07819747924805,
35.0527992248535,-3.98494005203247,
57.4635124206543,-2.45423698425293,
27.0008468627930,20.5862216949463,
-18.2807178497314,47.2191734313965,
-22.8671779632568,48.4516410827637,
12.1671504974365,27.9432487487793,
37.7959632873535,15.7595939636230,
25.4555377960205,28.5287971496582,
-10.0960531234741,48.0217819213867,
-35.6483802795410,53.1521148681641,
-40.6350479125977,37.1489715576172,
-35.2495422363281,9.30013847351074,
-26.5226535797119,-22.2265148162842,
-11.3988103866577,-48.1888198852539,
5.24654054641724,-51.4292449951172,
11.1741828918457,-25.4656009674072,
0.558194339275360,4.22610330581665,
-10.1635217666626,-1.91016149520874,
-2.99070477485657,-43.7624053955078,
19.5206985473633,-71.9617614746094,
34.9489402770996,-45.5264892578125,
21.6660995483398,11.3695735931396,
-9.28371810913086,31.9928512573242,
-27.8116226196289,-7.54863834381104,
-24.1974105834961,-61.8786697387695,
-13.7906227111816,-70.9501037597656,
-10.3156118392944,-33.3984069824219,
-5.03996562957764,7.93777751922607,
13.2846889495850,19.8093357086182,
29.3528175354004,17.2570362091064,
16.7533798217773,25.8852214813232,
-21.3933811187744,43.8219947814941,
-47.4947357177734,52.1523513793945,
-39.8236503601074,39.5719718933106,
-21.4776916503906,17.8696632385254,
-24.6516304016113,2.52652406692505,
-39.1818428039551,0.484949588775635,
-29.3039150238037,10.5574893951416,
10.1036472320557,26.6686992645264,
40.8237304687500,33.1365318298340,
27.5482406616211,28.3550014495850,
-9.49325656890869,21.5884933471680,
-21.2699432373047,21.9693756103516,
6.51981544494629,29.3903255462647,
38.2451438903809,27.1750869750977,
39.7625427246094,8.36339378356934,
17.6162242889404,-14.1972465515137,
0.678098082542419,-23.4366874694824,
0.447018802165985,-16.3594169616699,
3.52756738662720,-2.31432604789734,
5.90195798873901,6.64454698562622,
18.2646636962891,0.368238985538483,
35.9016075134277,-13.9658737182617,
32.5411605834961,-16.2437267303467,
-4.79924726486206,11.3480453491211,
-42.9062194824219,50.2637710571289,
-38.2232055664063,60.0444488525391,
7.03637886047363,22.3592376708984,
40.2341842651367,-24.0459728240967,
28.4142360687256,-29.4126205444336,
-5.96806097030640,3.45012474060059,
-20.0036983489990,23.1825904846191,
-5.45621395111084,-1.89137411117554,
15.5740671157837,-38.0052375793457,
23.3812980651855,-42.1045074462891,
23.6737709045410,-18.6833572387695,
22.2216606140137,-3.67850303649902,
15.3555021286011,-12.5195703506470,
2.07377862930298,-22.8917655944824,
-6.87747907638550,-20.1625576019287,
-8.75031471252441,-20.4029006958008,
-9.37993335723877,-36.3114585876465,
-7.68228340148926,-53.8196182250977,
8.30793952941895,-52.0736351013184,
35.5132064819336,-35.4379997253418,
49.5864486694336,-21.5109157562256,
36.0136566162109,-12.5588598251343,
13.5599937438965,9.93301773071289,
12.4507598876953,41.0083007812500,
29.8013496398926,51.7251892089844,
36.1476631164551,25.1874027252197,
22.1308860778809,-19.6702518463135,
13.1543149948120,-46.5496978759766,
28.4630603790283,-34.5715599060059,
51.3880119323731,-0.0268039703369141,
54.8911399841309,24.3610439300537,
42.2615661621094,17.5103454589844,
34.2640113830566,-11.1004953384399,
33.3603553771973,-34.1659545898438,
20.7227725982666,-26.1887855529785,
-9.84293365478516,1.77441930770874,
-33.8444976806641,11.9593992233276,
-27.2096214294434,-13.9791193008423,
1.75985383987427,-45.6888313293457,
25.5016613006592,-43.5542984008789,
27.8562602996826,-9.65227127075195,
13.0594253540039,12.6028633117676,
-4.34156560897827,1.08473670482636,
-16.6019248962402,-18.7556152343750,
-17.7410812377930,-13.3355684280396,
-8.06953239440918,5.47384548187256,
0.983284056186676,0.430351972579956,
-5.63874149322510,-26.8710231781006,
-23.3850517272949,-33.1713104248047,
-34.0378036499023,2.97606611251831,
-20.8075351715088,42.1487159729004,
4.59576272964478,34.3598785400391,
18.0121326446533,-15.0018205642700,
4.13714408874512,-47.4221954345703,
-17.3203468322754,-31.8439979553223,
-17.9396667480469,7.06748819351196,
7.98383045196533,24.6734600067139,
39.1269340515137,10.9556264877319,
42.9218711853027,-8.20803642272949,
10.9042034149170,-8.71076107025147,
-24.4584121704102,6.80690383911133,
-25.6344738006592,22.3956260681152,
4.97518157958984,24.4899272918701,
28.3855857849121,6.52447509765625,
23.6804828643799,-20.9243774414063,
13.8808393478394,-33.3397064208984,
28.4847106933594,-18.0615653991699,
50.9372138977051,10.2584562301636,
31.1630058288574,32.9397506713867,
-36.7282714843750,45.7967834472656,
-83.4016571044922,52.2235908508301,
-49.0955200195313,47.8459472656250,
24.3520832061768,22.5599994659424,
44.6241569519043,-10.2843618392944,
-9.03743743896484,-18.9125003814697,
-57.0800056457520,1.82011938095093,
-33.7663116455078,15.6135511398315,
19.4430866241455,-2.71229171752930,
21.6028156280518,-23.5166282653809,
-22.4748058319092,-10.4797925949097,
-33.0703125000000,20.4686260223389,
15.8762502670288,22.7306556701660,
51.4920616149902,-7.88245582580566,
13.4660282135010,-27.1222076416016,
-51.1236152648926,-10.1406669616699,
-63.1613235473633,13.3020935058594,
-24.8401165008545,6.49812412261963,
-5.16376781463623,-19.6338119506836,
-28.6705570220947,-30.8666496276855,
-49.2704238891602,-28.6304225921631,
-37.2002868652344,-31.8939399719238,
-20.5499019622803,-28.9966621398926,
-24.1236000061035,5.30697822570801,
-26.8864288330078,49.3186340332031,
-2.32560253143311,50.9690856933594,
20.9507102966309,5.02368879318237,
7.08304595947266,-28.3203945159912,
-20.0152854919434,-10.2571115493774,
-13.3690071105957,27.6469993591309,
17.3208427429199,29.8517723083496,
21.8560714721680,-1.59077334403992,
-5.49151659011841,-19.2533645629883,
-17.3054809570313,-10.9585990905762,
8.41523170471191,-10.3768186569214,
33.8338317871094,-21.7933826446533,
14.6465568542480,-8.31094551086426,
-30.4571743011475,34.5684890747070,
-51.6649055480957,53.7884712219238,
-43.9600296020508,18.5970706939697,
-40.1290168762207,-31.6669998168945,
-43.1526260375977,-41.7887573242188,
-31.8683376312256,-27.3301391601563,
-5.53194093704224,-37.3718872070313,
10.6610641479492,-69.3752212524414,
8.58308792114258,-62.9799652099609,
4.33422565460205,-6.89322519302368,
-0.0530546903610230,29.9515438079834,
-14.6892223358154,3.25542688369751,
-33.9814834594727,-36.6624870300293,
-27.9652328491211,-23.2222747802734,
7.52556419372559,22.1841640472412,
25.4677429199219,30.5400466918945,
-11.1164045333862,-3.02252435684204,
-62.9937438964844,-15.6657047271729,
-58.4633865356445,17.9767761230469,
3.70823764801025,47.6709671020508,
51.4358978271484,29.3247470855713,
45.2646751403809,-3.90603971481323,
17.2418098449707,6.46359634399414,
4.14024591445923,46.8380508422852,
-4.28232955932617,56.6832046508789,
-34.7156372070313,17.9850788116455,
-69.2805328369141,-26.0820827484131,
-66.1938171386719,-44.1225013732910,
-27.4793357849121,-36.4711112976074,
-0.131380796432495,-15.9654407501221,
-2.79540753364563,10.1389360427856,
-7.32869482040405,23.9824275970459,
5.84784030914307,6.66749620437622,
14.2653236389160,-25.2030868530273,
5.85030746459961,-25.0405941009522,
5.68860292434692,17.4198055267334,
30.7393779754639,49.6726837158203,
43.1612434387207,23.5937938690186,
5.02009773254395,-26.7603130340576,
-51.5777587890625,-30.2568244934082,
-61.0913734436035,13.1635904312134,
-15.3098754882813,33.1984138488770,
17.2545833587647,-9.17450046539307,
-6.33859252929688,-69.4428176879883,
-42.3392181396484,-80.2433700561523,
-31.3811607360840,-35.3452873229981,
4.22157526016235,10.9954652786255,
7.19696617126465,19.8935527801514,
-24.3960208892822,-2.09704709053040,
-30.3692283630371,-24.2205600738525,
14.8948669433594,-25.5613498687744,
61.6124992370606,-6.70322465896606,
53.9720993041992,23.3812332153320,
3.03118610382080,43.6105918884277,
-37.4478607177734,36.2170524597168,
-43.8969383239746,7.14305210113525,
-34.0654449462891,-17.2754955291748,
-23.1223754882813,-27.0491905212402,
-4.76002550125122,-26.5914516448975,
16.0391731262207,-19.5274009704590,
16.1328086853027,-7.59378242492676,
-10.1840400695801,-1.22793662548065,
-39.5372428894043,-9.17580127716065,
-48.2256622314453,-27.6619510650635,
-36.4443740844727,-24.0863304138184,
-19.3759880065918,18.8765296936035,
-7.22615003585815,61.4806938171387,
-0.296406924724579,52.7029724121094,
0.677284777164459,0.619458675384522,
-4.16992092132568,-35.2267990112305,
-6.96911859512329,-23.1105651855469,
1.94156622886658,-2.10746407508850,
13.2047643661499,-22.0567378997803,
13.2628068923950,-60.9046287536621,
7.92921733856201,-60.9934997558594,
11.0335350036621,-18.1220970153809,
21.5988273620605,5.32769012451172,
24.5473918914795,-27.3161640167236,
15.4913997650146,-66.5811996459961,
10.1733522415161,-41.4114685058594,
16.7821331024170,32.2945098876953,
28.2935581207275,70.5994949340820,
27.6379470825195,33.5574722290039,
16.7936611175537,-21.5892505645752,
5.46423864364624,-18.7966518402100,
-4.71830320358276,37.1923637390137,
-16.1098594665527,78.3487472534180,
-21.1212768554688,58.3432121276856,
-8.56875228881836,1.69514441490173,
13.0685815811157,-31.5179233551025,
18.1456050872803,-21.6809120178223,
-2.77863454818726,3.67801856994629,
-28.3434276580811,9.29918003082275,
-39.8784751892090,-11.3869647979736,
-40.9563751220703,-37.3615837097168,
-47.1713638305664,-44.9331207275391,
-57.6049652099609,-27.9015216827393,
-52.6952514648438,-5.60797214508057,
-27.6522312164307,9.71492481231690,
-2.39384365081787,17.2739830017090,
9.65369987487793,17.8116302490234,
23.1408100128174,9.29094982147217,
46.5886650085449,-3.60612154006958,
65.5062179565430,-4.69768095016480,
59.0299758911133,17.5601062774658,
33.5487632751465,51.6367263793945,
12.2005548477173,60.3757438659668,
-1.34512460231781,29.8701820373535,
-24.9074020385742,-12.9025945663452,
-53.4118957519531,-35.4995117187500,
-52.2672691345215,-39.7198295593262,
-11.6137733459473,-45.8630065917969,
25.1715641021729,-56.4143600463867,
12.3992786407471,-54.4173393249512,
-29.0615425109863,-36.7321815490723,
-31.5914497375488,-26.3474388122559,
18.5767707824707,-33.9303054809570,
63.9839630126953,-35.8826026916504,
56.3515396118164,-5.77318954467773,
17.9563713073730,38.9663734436035,
4.79976940155029,57.7312240600586,
22.5488262176514,44.5582008361816,
29.0422554016113,33.7745018005371,
0.803927361965179,42.6068801879883,
-29.1297435760498,43.2524871826172,
-24.4082794189453,3.78317546844482,
7.98238849639893,-47.3017768859863,
31.2931842803955,-54.8882675170898,
23.9924335479736,-8.83066368103027,
-3.63778018951416,41.7243766784668,
-30.9218654632568,51.8860588073731,
-34.2642250061035,30.2541122436523,
-8.96361160278320,13.7243347167969,
26.4306221008301,14.2955465316772,
42.3794021606445,13.3096876144409,
24.3550834655762,-1.64654254913330,
-9.90040969848633,-14.9310932159424,
-24.4026012420654,-17.7824287414551,
-12.2964468002319,-21.6955814361572,
6.30542325973511,-40.4016876220703,
12.8258075714111,-64.6626434326172,
9.90238285064697,-65.3781356811523,
3.49339866638184,-35.5363159179688,
-6.26629972457886,0.539913594722748,
-14.8123130798340,8.22595596313477,
-9.94139671325684,-12.4605350494385,
16.0370197296143,-22.3518905639648,
42.8415908813477,1.73748946189880,
40.3620986938477,39.0665016174316,
6.98277950286865,46.5583267211914,
-20.3905143737793,12.3245801925659,
-12.1530036926270,-33.3042984008789,
19.5709915161133,-57.0694923400879,
34.4218864440918,-57.3424110412598,
20.7827873229980,-46.4097328186035,
4.41329908370972,-24.2095184326172,
10.2130165100098,10.3791618347168,
27.8172836303711,37.6430397033691,
30.5495662689209,30.7486228942871,
16.7604198455811,3.35102653503418,
9.73410224914551,-5.82821607589722,
21.8470420837402,16.7278118133545,
36.8279991149902,38.4290847778320,
39.3720626831055,30.2833557128906,
34.7185783386231,7.90234470367432,
39.6665344238281,5.04556179046631,
46.3265533447266,16.7447299957275,
38.0192070007324,16.7481708526611,
18.6351127624512,2.09290218353272,
8.89391803741455,-0.0713315606117249,
20.3793888092041,16.2659072875977,
32.4237747192383,17.0719165802002,
23.6801071166992,-10.5215148925781,
4.04077196121216,-35.0420303344727,
0.718028247356415,-16.9732799530029,
21.4473171234131,26.2490863800049,
40.5754356384277,34.9470329284668,
36.9943542480469,-5.83750438690186,
20.3177490234375,-44.4294013977051,
18.6545047760010,-30.5237827301025,
42.5200576782227,22.1454086303711,
70.6371612548828,52.8964004516602,
65.2804336547852,34.7623748779297,
20.9687995910645,4.66535139083862,
-30.2376823425293,2.79942035675049,
-57.5553169250488,16.4773559570313,
-57.6110076904297,5.21015691757202,
-46.0573577880859,-37.0843200683594,
-29.4616565704346,-61.3357849121094,
-2.62527418136597,-30.3788013458252,
29.4565277099609,28.7137966156006,
36.7953147888184,55.3432235717773,
10.0502891540527,31.1474876403809,
-15.1902866363525,-3.11398267745972,
-3.10751891136169,-3.94322776794434,
25.3051300048828,26.5336284637451,
16.5537300109863,51.5632781982422,
-35.5909385681152,50.1620750427246,
-66.5790786743164,25.7138023376465,
-32.1828346252441,-5.04498815536499,
27.0187053680420,-18.5360260009766,
34.7213745117188,-0.902193009853363,
-12.9140539169312,39.1461257934570,
-45.6947135925293,59.8948554992676,
-14.5255365371704,35.4173049926758,
42.2718887329102,-4.60248088836670,
57.9437332153320,-6.75550746917725,
22.3804397583008,26.0675392150879,
-20.4341735839844,37.6541252136231,
-30.1518077850342,-1.00887846946716,
-12.1210823059082,-47.5252799987793,
10.2442111968994,-37.5680122375488,
19.1714687347412,19.8335628509522,
8.67716121673584,52.5785636901856,
-14.1823444366455,25.8089370727539,
-27.9246025085449,-25.3385143280029,
-17.1444244384766,-52.0470733642578,
9.59884548187256,-47.2750358581543,
29.6524639129639,-35.2586212158203,
28.9235248565674,-28.6306571960449,
21.1964969635010,-22.1697139739990,
27.2610244750977,-19.3560256958008,
42.8208656311035,-18.6739101409912,
54.0812873840332,-5.41928100585938,
57.4408569335938,28.1138229370117,
47.3737106323242,56.8168754577637,
19.3192081451416,44.1252899169922,
-19.7241668701172,-7.18509292602539,
-49.1650733947754,-41.5286483764648,
-50.3634071350098,-14.1847457885742,
-33.3878898620606,43.9513816833496,
-23.7278156280518,72.0669250488281,
-23.0538635253906,48.1778450012207,
-10.7832307815552,6.24752330780029,
14.3139209747314,-5.65659046173096,
19.3527603149414,21.3224887847900,
-16.6112442016602,49.7495307922363,
-54.9101257324219,43.8258247375488,
-41.4858093261719,2.03226208686829,
15.3976831436157,-34.5583648681641,
51.6104736328125,-27.5669593811035,
27.5051002502441,16.0503768920898,
-24.1771106719971,40.9316978454590,
-43.3654098510742,2.05657243728638,
-18.9363899230957,-70.3057403564453,
16.5934944152832,-96.9619140625000,
37.1403236389160,-48.5234222412109,
43.5581436157227,16.2505798339844,
38.5623588562012,33.3366966247559,
13.4323835372925,6.74531793594360,
-14.4343147277832,-10.4369087219238,
-12.4368619918823,5.60247087478638,
20.9214744567871,21.3461894989014,
40.4086875915527,17.6447315216064,
14.2417507171631,22.9434032440186,
-32.3841514587402,52.6289215087891,
-53.8577880859375,66.8935699462891,
-40.9280853271484,24.3183574676514,
-22.6132774353027,-44.5787200927734,
-14.0011234283447,-69.8138351440430,
1.68126082420349,-39.3729362487793,
28.8051929473877,-14.3602266311646,
39.1704025268555,-32.6814041137695,
27.7323989868164,-53.9456901550293,
23.7572689056397,-33.1463813781738,
42.4896278381348,11.8232498168945,
54.6762428283691,23.3755722045898,
30.7047672271729,-8.13109493255615,
-2.66246914863586,-29.0025043487549,
2.46257042884827,-7.63937854766846,
35.3812599182129,24.8993415832520,
42.1522750854492,32.3183975219727,
5.59260749816895,20.4689826965332,
-28.5382595062256,14.5105743408203,
-17.4581356048584,18.4537849426270,
6.72963285446167,18.4393768310547,
-6.44232559204102,7.23207759857178,
-48.0037956237793,-9.25572109222412,
-66.6084899902344,-17.0733203887939,
-44.7558860778809,-14.2876319885254,
-12.8199119567871,0.105739414691925,
5.33396720886231,10.6651172637939,
14.5950632095337,-5.09906959533691,
29.7447090148926,-51.4359893798828,
43.5264663696289,-81.7252044677734,
50.2924728393555,-49.6878204345703,
52.8719291687012,22.1109371185303,
49.6599540710449,57.4216232299805,
20.6760902404785,28.0836601257324,
-31.8650321960449,-15.4499578475952,
-62.8209419250488,-15.9792079925537,
-31.9007129669189,10.7009267807007,
24.8200912475586,6.11882781982422,
38.3707580566406,-36.3878173828125,
0.313644886016846,-65.5432891845703,
-27.9959831237793,-54.4767494201660,
-0.830251693725586,-39.0347557067871,
51.2864074707031,-47.8618812561035,
63.5007972717285,-48.3976974487305,
26.8858261108398,-2.83890008926392,
-14.8556909561157,63.2748718261719,
-30.4675540924072,88.2973327636719,
-28.9642639160156,60.6816749572754,
-27.5631370544434,33.8878669738770,
-23.5811653137207,38.9410400390625,
-16.3044166564941,49.7870101928711,
-17.7962207794189,30.8541793823242,
-30.1523647308350,-7.46430444717407,
-28.8303947448730,-26.6362838745117,
1.33037281036377,-22.4835128784180,
38.4575653076172,-22.3042888641357,
47.9462699890137,-26.0063591003418,
23.3515644073486,-8.45456504821777,
-9.73529148101807,26.9488048553467,
-21.9288272857666,48.7948532104492,
-14.5445365905762,31.4157638549805,
-5.32316780090332,-2.01650619506836,
-0.185214832425118,-18.4667968750000,
-0.352320343255997,-10.9073476791382,
2.33252263069153,5.70669651031494,
14.6693658828735,15.5990352630615,
34.0672149658203,20.4824790954590,
44.1341476440430,11.2581110000610,
26.6317920684814,-12.1968736648560,
-9.31861305236816,-23.2085151672363,
-34.6527519226074,5.08454084396362,
-38.0677375793457,48.7461738586426,
-35.4921188354492,53.5957603454590,
-45.8023223876953,2.99312877655029,
-62.1237335205078,-57.9067039489746,
-56.1722183227539,-80.0444107055664,
-17.8185672760010,-61.9190025329590,
32.1312065124512,-30.4963378906250,
65.9289093017578,1.30158257484436,
69.0999526977539,39.6341018676758,
41.9245948791504,64.1904602050781,
0.298494815826416,43.1188430786133,
-25.4844646453857,-6.99663448333740,
-13.7677154541016,-27.3796634674072,
16.8185081481934,1.72267961502075,
20.9274692535400,34.9154930114746,
-19.6857547760010,24.3626899719238,
-65.2805023193359,-9.95896530151367,
-65.7502288818359,-18.9003372192383,
-23.2554569244385,-2.86427330970764,
8.57945537567139,1.56825065612793,
2.23059678077698,-11.9973545074463,
-17.0769081115723,-6.60831212997437,
-7.99975824356079,32.6742858886719,
20.2324085235596,55.4938430786133,
29.8892879486084,28.1063461303711,
14.7819366455078,-11.6361417770386,
0.356697380542755,-8.15441131591797,
9.18003273010254,31.4931316375732,
26.4646339416504,44.3291091918945,
30.2735061645508,10.5122966766357,
24.3069858551025,-29.5859909057617,
24.6301593780518,-34.5965919494629,
25.3623580932617,-13.1085271835327,
11.6189279556274,5.14395046234131,
-17.7946319580078,8.34997558593750,
-43.0861206054688,7.01702117919922,
-52.4932823181152,-4.12826681137085,
-51.6382141113281,-30.2075157165527,
-38.5430221557617,-49.7029418945313,
-3.58020305633545,-32.9660224914551,
42.0254478454590,12.9989395141602,
60.9620857238770,49.3141555786133,
30.1304035186768,57.2065505981445,
-22.0529270172119,49.3396949768066,
-46.0731201171875,47.1680870056152,
-31.9012813568115,53.4753265380859,
-19.8764095306397,54.6167221069336,
-38.4428825378418,41.5682907104492,
-68.2111129760742,13.3227157592773,
-73.2980880737305,-27.2390213012695,
-50.2033195495606,-67.1807327270508,
-29.9602108001709,-80.8765945434570,
-27.1409187316895,-57.1083793640137,
-27.3778152465820,-22.2391395568848,
-14.4458265304565,-7.56906414031982,
2.60590028762817,-11.9157295227051,
3.45157313346863,-6.62212610244751,
-15.8955774307251,18.1269245147705,
-35.4288482666016,35.1459960937500,
-38.3018302917481,18.4056415557861,
-39.3739471435547,-22.6882553100586,
-53.0084114074707,-48.7249221801758,
-67.0470581054688,-45.6382217407227,
-50.0225753784180,-28.0051860809326,
3.96746134757996,-16.3177661895752,
51.2424774169922,-8.83823585510254,
44.3990783691406,-3.82051348686218,
-8.00022792816162,-10.1794471740723,
-42.5196990966797,-32.6790199279785,
-23.9942836761475,-53.3848915100098,
15.2255363464355,-42.2623329162598,
21.6793212890625,-3.84940934181213,
-4.03336000442505,31.4879627227783,
-14.7901506423950,36.9786796569824,
10.8642625808716,25.4440422058105,
43.5500068664551,22.4587192535400,
46.8585700988770,33.1901893615723,
31.2107143402100,39.9097328186035,
24.5319786071777,31.1565628051758,
31.9495792388916,16.0687408447266,
28.8111267089844,2.77126979827881,
13.2380352020264,-6.50353574752808,
2.00773715972900,-12.3754911422730,
4.09172534942627,-8.26430702209473,
5.25127792358398,7.60180282592773,
-8.47888946533203,22.5153236389160,
-20.8114032745361,25.5363979339600,
-16.9487991333008,23.8839397430420,
-10.7843103408813,32.3761520385742,
-20.8684158325195,51.4216690063477,
-43.0792198181152,56.5694656372070,
-52.1868515014648,33.8117256164551,
-39.2183113098145,-4.52304601669312,
-25.8281173706055,-32.1602783203125,
-34.7289543151856,-38.6684608459473,
-54.6124534606934,-28.3657760620117,
-59.3512611389160,-12.6027803421021,
-37.7398223876953,4.16687679290772,
-8.16235065460205,21.6258163452148,
5.45134449005127,32.3150444030762,
-6.24327421188355,24.4958019256592,
-31.7718238830566,-1.56750607490540,
-47.4722099304199,-27.0659122467041,
-35.7036590576172,-29.5520477294922,
0.713046550750732,-3.79370999336243,
39.2208518981934,24.8403015136719,
50.0820770263672,22.1056480407715,
28.5146522521973,-7.33264732360840,
-0.725850939750671,-20.9247055053711,
-10.4190845489502,6.90744304656982,
2.78933000564575,40.7276000976563,
18.3789882659912,27.8727035522461,
17.1814098358154,-27.9991989135742,
5.73293685913086,-60.9699974060059,
-4.62678956985474,-31.1420307159424,
-11.9612102508545,22.4655685424805,
-25.4907493591309,34.1804771423340,
-38.9010658264160,4.10224771499634,
-35.4104309082031,-12.2396812438965,
-17.2059478759766,8.01059532165527,
-14.4622268676758,28.2034683227539,
-41.7473831176758,12.8364686965942,
-72.6941986083984,-16.5329399108887,
-60.2683334350586,-15.9733743667603,
-2.38073062896729,7.84626054763794,
46.5225830078125,15.1881980895996,
42.0914154052734,-5.17490911483765,
0.0178995132446289,-20.0657539367676,
-30.9839649200439,-6.01012516021729,
-29.6979312896729,15.6772699356079,
-14.5087518692017,6.72151184082031,
-4.00216484069824,-32.5692062377930,
-0.868140816688538,-56.3827781677246,
-3.56395506858826,-38.0602111816406,
-16.3313179016113,0.647792816162109,
-31.3512058258057,18.4454345703125,
-22.4712333679199,-1.64145147800446,
14.0478410720825,-31.5148468017578,
43.5651855468750,-26.0672092437744,
32.0813713073731,19.9111557006836,
-3.45391130447388,62.9460334777832,
-14.0880041122437,62.7242469787598,
12.5589752197266,30.7896823883057,
33.4308700561523,10.8011503219605,
18.4731502532959,19.6034336090088,
-6.48240756988525,22.7895298004150,
-3.40342259407043,-10.4831180572510,
26.3212833404541,-51.9464263916016,
42.4842987060547,-46.7466430664063,
23.4571094512939,4.06915616989136,
-6.64709663391113,34.2591247558594,
-17.5239353179932,7.68549728393555,
-6.46535539627075,-35.0660858154297,
9.90927219390869,-30.9036960601807,
15.3244590759277,17.1490859985352,
3.31332015991211,46.7031288146973,
-23.7361621856689,25.8768501281738,
-46.6052398681641,-3.92712879180908,
-40.2733879089356,1.22286486625671,
-9.70235347747803,27.3774719238281,
8.49352836608887,34.4740142822266,
-6.60952568054199,16.8788013458252,
-30.4057197570801,7.14389276504517,
-21.3605308532715,12.4803743362427,
19.5907859802246,4.07065820693970,
50.0823097229004,-29.0252723693848,
40.0428962707520,-50.9574394226074,
9.86698722839356,-33.4923973083496,
-8.14079666137695,6.38433361053467,
-11.9630737304688,29.4485816955566,
-17.2898101806641,25.3097419738770,
-26.2093391418457,20.4018707275391,
-25.0822315216064,30.5183601379395,
-11.1069335937500,39.7423019409180,
4.93765735626221,33.0964202880859,
13.0507316589355,17.9897212982178,
17.6369152069092,3.44288635253906,
20.9862461090088,-10.5645418167114,
22.2925968170166,-21.5213489532471,
23.5658683776855,-16.5189800262451,
28.6427688598633,-1.42387962341309,
32.3778839111328,-1.31867265701294,
21.7620048522949,-24.8522377014160,
-5.01964855194092,-42.7406044006348,
-25.1423168182373,-20.2458477020264,
-21.1363105773926,31.1540775299072,
-7.36196279525757,54.5308456420898,
-14.4434251785278,25.2626190185547,
-47.3892478942871,-19.9391422271729,
-76.6520767211914,-36.5137023925781,
-70.0798797607422,-20.3836212158203,
-28.2209529876709,-2.54403877258301,
12.1773433685303,0.280612915754318,
19.4779090881348,-9.86233806610107,
-4.29435396194458,-24.0555915832520,
-27.1404685974121,-37.4780349731445,
-21.7665557861328,-35.1060829162598,
9.14412307739258,-4.33282470703125,
31.2428665161133,35.1147537231445,
17.1237602233887,43.0403594970703,
-19.4864215850830,1.79385876655579,
-33.3070678710938,-48.4553871154785,
-5.40174579620361,-53.8664093017578,
33.1779708862305,-11.8472862243652,
42.9509963989258,32.1820297241211,
24.5913639068604,41.7937431335449,
16.2800102233887,19.8611373901367,
35.5837097167969,-9.55204296112061,
53.5278053283691,-27.0476989746094,
36.3792381286621,-31.2164173126221,
8.62151527404785,-28.2334880828857,
13.1474819183350,-23.5528488159180,
48.2968482971191,-17.4358501434326,
62.2629508972168,-4.70427322387695,
29.4654312133789,24.5309658050537,
-7.27938127517700,57.2647972106934,
0.332311511039734,63.3530502319336,
31.8332176208496,34.0971260070801,
32.2493057250977,1.33551347255707,
-6.20516061782837,-9.54766368865967,
-28.3646793365479,-10.7007379531860,
-2.12426400184631,-25.8771438598633,
34.0702590942383,-44.3795394897461,
28.0030193328857,-34.9824981689453,
-6.62138223648071,-3.48983502388001,
-14.6432094573975,1.76812076568604,
25.0822391510010,-33.8723945617676,
68.4776382446289,-54.2353401184082,
72.4255752563477,-9.64569091796875,
35.1245498657227,61.9940071105957,
-11.1444482803345,71.5853347778320,
-36.9606895446777,7.49271392822266,
-29.5556526184082,-48.0156593322754,
4.70737266540527,-27.2014789581299,
49.4706764221191,40.1660537719727,
72.3535461425781,75.8730010986328,
53.7683029174805,55.9307060241699,
10.9872369766235,19.1979713439941,
-16.7998142242432,-0.0870138406753540,
-9.18402290344238,-10.7059717178345,
23.5990810394287,-17.6222972869873,
51.7989196777344,-7.70913314819336,
46.4498023986816,25.0051002502441,
7.22590446472168,52.0269279479981,
-30.9977684020996,48.3649559020996,
-33.1132431030273,30.4102573394775,
0.591607093811035,31.4621925354004,
30.4604148864746,42.9975395202637,
12.6599607467651,31.6051445007324,
-36.8518257141113,-9.86185359954834,
-62.9681282043457,-47.8617591857910,
-41.5740432739258,-49.2734336853027,
-11.6654014587402,-26.8346729278564,
-17.4528198242188,-22.7928066253662,
-38.0794754028320,-48.9316596984863,
-27.9632263183594,-73.4362792968750,
11.7438077926636,-59.9614944458008,
27.6178760528564,-17.0849494934082,
-7.12275028228760,10.6154098510742,
-43.7875900268555,-3.68139481544495,
-22.8743858337402,-39.8072738647461,
30.7274055480957,-47.4988212585449,
45.6218070983887,-6.71879005432129,
3.76170730590820,41.7406768798828,
-41.3835830688477,53.7302589416504,
-44.1052970886231,30.0980606079102,
-28.4323616027832,9.62118434906006,
-32.7586288452148,10.0148811340332,
-38.5418777465820,9.80462932586670,
-8.83449172973633,-11.6837234497070,
37.8763923645020,-30.3101844787598,
42.3495788574219,-12.8325281143188,
-4.36688852310181,22.2107257843018,
-39.9999923706055,18.3072719573975,
-13.7713003158569,-32.6335372924805,
41.1727638244629,-69.1772689819336,
55.6439056396484,-41.0078506469727,
19.2863445281982,17.2873954772949,
-11.6660585403442,28.6528244018555,
1.47783648967743,-21.0221405029297,
33.8025245666504,-58.4804801940918,
43.8369560241699,-28.2715759277344,
19.6332836151123,29.0934524536133,
-11.7251987457275,37.6111335754395,
-27.4430599212647,-9.07506179809570,
-31.9981784820557,-46.0046958923340,
-37.1952095031738,-33.1949005126953,
-39.0260238647461,-2.36745524406433,
-23.1091461181641,5.07086801528931,
4.07417917251587,5.13966560363770,
18.1742973327637,27.9732303619385,
3.57729005813599,54.8989868164063,
-24.1701965332031,42.3559188842773,
-25.3939285278320,-6.04299020767212,
10.5279283523560,-35.1566429138184,
41.8721351623535,-14.8831977844238,
26.3874816894531,14.1550369262695,
-24.1831417083740,7.09570264816284,
-57.0350914001465,-17.1633872985840,
-48.7358512878418,-12.1712455749512,
-26.5558071136475,23.3364353179932,
-24.8379974365234,46.4052124023438,
-32.9438133239746,34.0211486816406,
-16.4717445373535,2.40184450149536,
19.7185459136963,-22.9352149963379,
30.8137035369873,-32.4589271545410,
-0.461276531219482,-23.7815856933594,
-37.9275932312012,5.15462732315064,
-41.5429992675781,38.2799911499023,
-19.8218898773193,41.7550239562988,
-8.48380661010742,8.07147884368897,
-11.4693136215210,-22.0451774597168,
-0.528676867485046,-13.2973279953003,
29.2361106872559,11.4837789535522,
40.7114486694336,8.59115600585938,
15.3185596466064,-27.8403549194336,
-13.6040811538696,-60.7894668579102,
-3.43142533302307,-61.0864524841309,
35.1395835876465,-35.5496597290039,
41.7041969299316,-9.94911479949951,
-4.62507200241089,3.83874869346619,
-56.0991516113281,3.41563534736633,
-62.0638046264648,-13.8134317398071,
-28.1315441131592,-37.7476806640625,
3.19863986968994,-44.9260559082031,
10.9101514816284,-26.3240013122559,
7.97016668319702,-8.67456150054932,
12.9019498825073,-19.2240638732910,
21.2615051269531,-40.3017234802246,
27.6225299835205,-37.1269912719727,
36.9997787475586,-8.40791702270508,
47.3921508789063,19.4974288940430,
47.9735679626465,29.4785614013672,
40.8789329528809,32.4534683227539,
42.6117744445801,40.8172035217285,
46.1593437194824,46.1892242431641,
21.3580265045166,36.2097358703613,
-33.9789237976074,25.6231212615967,
-70.2314376831055,25.2669506072998,
-47.1499137878418,17.0727310180664,
2.95984172821045,-10.8937911987305,
13.8295936584473,-31.6352462768555,
-26.3611869812012,-11.2871398925781,
-50.1990814208984,27.1472187042236,
-17.4246997833252,23.7006549835205,
27.5059013366699,-30.2367229461670,
25.7411174774170,-67.6932678222656,
-9.53379917144775,-39.1602706909180,
-22.1672439575195,19.8860492706299,
-0.687050580978394,34.2070198059082,
11.0079460144043,-4.93949937820435,
-6.64522552490234,-31.9656391143799,
-21.3177928924561,-13.4330987930298,
-6.94251823425293,9.78054428100586,
14.3487167358398,-5.43550634384155,
13.8380479812622,-39.4964179992676,
6.87081003189087,-48.4329071044922,
26.7287864685059,-24.5721092224121,
59.6052589416504,3.10369253158569,
58.2341728210449,16.8948173522949,
14.5825500488281,19.0355968475342,
-27.6339282989502,7.13689708709717,
-32.7703819274902,-21.4460659027100,
-13.1859788894653,-41.7582550048828,
-2.51449441909790,-19.9789409637451,
-12.5126447677612,31.1910858154297,
-29.7999973297119,51.0915565490723,
-34.6716003417969,17.6318988800049,
-16.1282310485840,-16.8247051239014,
21.3726863861084,0.920361757278442,
57.1084785461426,44.6808700561523,
58.0747451782227,49.4660148620606,
11.8395023345947,6.93417930603027,
-46.9147605895996,-22.8202228546143,
-68.5613250732422,-1.24948227405548,
-43.5342254638672,35.6335487365723,
-3.21678018569946,30.4133739471436,
23.0166511535645,-8.30047130584717,
24.6808719635010,-28.4339199066162,
6.30706119537354,-7.46269273757935,
-20.1472625732422,18.8848590850830,
-38.1864891052246,14.8944797515869,
-22.9734458923340,-14.2115421295166,
21.9447898864746,-39.0047645568848,
58.7104835510254,-39.9981613159180,
54.5601005554199,-14.9761714935303,
25.4319152832031,17.7000122070313,
10.5358428955078,36.9931564331055,
20.9519824981689,30.6679592132568,
24.0836486816406,9.37928771972656,
-3.03743839263916,-2.26431083679199,
-31.3234844207764,8.48157691955566,
-22.5910701751709,25.6672115325928,
15.2321596145630,27.9338035583496,
36.0649452209473,25.1702213287354,
5.33242511749268,35.3831977844238,
-49.8223381042481,49.0978965759277,
-77.3900985717773,41.4715042114258,
-54.1632957458496,16.8283405303955,
-8.79595851898193,9.62347316741943,
12.4061412811279,35.9526138305664,
-6.15038108825684,60.4581375122070,
-39.1194000244141,36.1544837951660,
-46.9722023010254,-29.4532604217529,
-16.8306560516357,-80.0205612182617,
20.1789817810059,-78.8240966796875,
25.2575569152832,-37.9333686828613,
-2.97576689720154,4.52007007598877,
-25.5899276733398,32.8463745117188,
-12.1619901657105,48.1037445068359,
24.3030300140381,49.1975021362305,
46.2165489196777,36.0655174255371,
40.1173477172852,22.0279712677002,
28.0297355651855,21.0889244079590,
30.5569438934326,23.9239368438721,
31.2287158966064,14.1749572753906,
12.4169435501099,-5.21894931793213,
-21.6712093353272,-7.32847166061401,
-44.5517387390137,20.1570167541504,
-44.6913032531738,52.1538124084473,
-35.8633651733398,46.4408645629883,
-31.4065036773682,1.69229006767273,
-25.1123981475830,-43.0533905029297,
-9.86026477813721,-52.2388839721680,
4.43360805511475,-26.5324249267578,
4.05951499938965,-1.60446751117706,
-9.42271709442139,1.16736757755280,
-18.9877319335938,-5.10172176361084,
-22.8418254852295,0.943202853202820,
-32.3421478271484,21.3650703430176,
-49.5370254516602,28.3652667999268,
-57.5250701904297,9.38128757476807,
-42.8687438964844,-14.6467752456665,
-19.3346633911133,-13.0381660461426,
-4.52038955688477,16.0809097290039,
1.39295864105225,40.2166023254395,
10.8685884475708,34.6450233459473,
27.0001316070557,13.7026634216309,
31.7599964141846,13.7176628112793,
22.0651092529297,39.5985908508301,
9.73092555999756,61.2792015075684,
3.78646469116211,56.1224174499512,
-10.2876319885254,26.2658157348633,
-39.2200698852539,-5.57158517837524,
-61.6913108825684,-29.2156066894531,
-51.2108001708984,-46.9202003479004,
-10.0803060531616,-51.7656631469727,
31.2268562316895,-33.6793594360352,
47.8602752685547,-0.861307740211487,
41.1941413879395,17.1773319244385,
23.9251441955566,10.5586118698120,
-1.64644777774811,2.61085700988770,
-30.4353771209717,15.6703758239746,
-49.9796638488770,28.6843185424805,
-51.0806694030762,4.63219738006592,
-39.0693969726563,-48.9239501953125,
-21.4907684326172,-75.9634552001953,
5.83893871307373,-41.9228630065918,
35.5674400329590,11.8576011657715,
42.9640998840332,26.7628574371338,
16.2970466613770,-3.68497967720032,
-21.4553146362305,-29.8682594299316,
-28.4510402679443,-25.6471176147461,
-1.82154107093811,-19.6830196380615,
23.6493949890137,-34.8795776367188,
18.9542808532715,-53.4409523010254,
-1.92519819736481,-41.1532325744629,
-14.4009704589844,-12.5428438186646,
-18.4918251037598,-9.22094917297363,
-23.9341220855713,-39.4120903015137,
-19.2888183593750,-58.6184043884277,
8.12945365905762,-29.8787441253662,
31.7724895477295,29.3324279785156,
16.9716854095459,64.8465881347656,
-31.0032958984375,46.8607177734375,
-57.0421485900879,-0.229543924331665,
-25.9180278778076,-37.2219734191895,
28.5191650390625,-39.5153884887695,
51.0640296936035,-7.80673456192017,
32.2430343627930,34.0014419555664,
9.06791591644287,61.2308197021484,
4.68977117538452,64.6267318725586,
6.08504915237427,48.6026649475098,
1.64286983013153,24.9970436096191,
5.19822883605957,7.94588994979858,
17.0617389678955,6.64195537567139,
14.3775310516357,20.0244789123535,
-17.3007678985596,32.8176155090332,
-50.9156303405762,24.1219406127930,
-45.6433486938477,-12.6007499694824,
-3.87241888046265,-42.3560600280762,
33.5508956909180,-28.7744884490967,
36.3543777465820,10.3210048675537,
18.0561542510986,24.6438789367676,
7.05282783508301,-5.49115705490112,
7.76456308364868,-38.0826568603516,
7.93073987960815,-26.4418449401855,
2.28700852394104,10.0577840805054,
-11.0153188705444,10.2841243743896,
-30.6117839813232,-31.4244403839111,
-49.9513626098633,-53.6182594299316,
-50.9988479614258,-15.6212444305420,
-25.7364120483398,32.6029434204102,
12.8981046676636,19.1687831878662,
38.8255653381348,-40.8800582885742,
39.7636528015137,-63.9577598571777,
26.0393123626709,-15.5700473785400,
18.0169105529785,38.2960662841797,
20.0925903320313,32.2731590270996,
25.7340526580811,-9.41837692260742,
22.1542987823486,-15.9514980316162,
1.56933760643005,23.9441986083984,
-25.0299644470215,48.0379142761231,
-36.5701675415039,16.6133861541748,
-22.6509838104248,-31.7578582763672,
-2.74860119819641,-41.8590011596680,
-5.86057853698731,-10.8513879776001,
-30.9771556854248,21.8202705383301,
-49.7549476623535,33.5623474121094,
-41.0198860168457,29.8986988067627,
-17.3820838928223,17.2721347808838,
-4.62400484085083,8.01051712036133,
-10.6220407485962,16.7795143127441,
-22.4054317474365,41.7439727783203,
-30.8864421844482,57.1172447204590,
-31.4473896026611,32.3603973388672,
-19.9107742309570,-16.8332443237305,
7.80453014373779,-31.8057575225830,
37.0692367553711,4.70088052749634,
43.2745018005371,41.5698471069336,
25.0041122436523,28.4953041076660,
9.36403083801270,-19.3418083190918,
16.5866394042969,-54.1105155944824,
34.0687026977539,-53.0292472839356,
32.2760658264160,-26.6930046081543,
7.27545261383057,7.57357406616211,
-16.3600730895996,35.6127548217773,
-21.0337486267090,35.3628120422363,
-12.6761713027954,-7.48010063171387,
-2.34736299514771,-55.9664878845215,
12.2894096374512,-45.9739761352539,
28.5654659271240,19.0350532531738,
25.5247955322266,64.5865020751953,
-6.89622259140015,39.8878440856934,
-41.3166961669922,-7.18923425674439,
-35.3746643066406,-9.78101253509522,
7.45572614669800,18.4138069152832,
34.3378829956055,14.7697257995605,
9.81463623046875,-22.3110923767090,
-40.4006271362305,-32.7600746154785,
-57.9553718566895,5.43330860137939,
-31.6496639251709,30.3233318328857,
1.44005370140076,-9.83443546295166,
10.8801622390747,-64.6319961547852,
8.38112640380859,-51.5368194580078,
12.7997503280640,21.6532554626465,
19.1053676605225,70.9815521240234,
15.0919113159180,54.0759201049805,
4.57051944732666,15.6592388153076,
-0.272208333015442,7.19779396057129,
-2.29449582099915,21.9648113250732,
-12.8348894119263,30.6163520812988,
-21.2220573425293,28.5694751739502,
-10.6574802398682,28.0167026519775,
9.35739612579346,26.7356033325195,
3.56368136405945,12.5054750442505,
-31.2389965057373,-4.70747756958008,
-53.6451606750488,-4.55518102645874,
-35.6814193725586,4.37647008895874,
-4.26144075393677,-5.11078929901123,
2.52066850662231,-29.4982852935791,
-9.48361110687256,-33.0348434448242,
-2.83644962310791,-2.78190302848816,
24.0641422271729,28.0060997009277,
25.3654174804688,31.8908386230469,
-18.6447830200195,16.1440639495850,
-62.8306961059570,3.18286943435669,
-58.4258880615234,-8.00249195098877,
-22.4326000213623,-28.4272651672363,
-10.4575834274292,-47.2977485656738,
-35.1258430480957,-38.9766921997070,
-48.5456466674805,-7.76640796661377,
-18.5386657714844,9.56934547424316,
25.5438747406006,-11.8244724273682,
39.3247108459473,-48.0563430786133,
21.1259841918945,-58.3442802429199,
4.49337959289551,-31.4239311218262,
5.48008489608765,4.17660760879517,
2.35307836532593,18.2379570007324,
-17.1849613189697,4.53441619873047,
-34.0886993408203,-17.7434711456299,
-26.0939884185791,-24.4170074462891,
0.572412490844727,-11.9795494079590,
15.0486049652100,4.40365314483643,
1.70236575603485,6.49320745468140,
-23.5008850097656,-4.33331966400147,
-28.8387584686279,-11.5300064086914,
-4.41817760467529,-5.58382081985474,
27.7033042907715,7.31280708312988,
32.1919937133789,5.97284269332886,
-2.79545164108276,-12.9406518936157,
-51.2218170166016,-34.7032318115234,
-70.4096069335938,-49.6928062438965,
-39.0938987731934,-55.9295692443848,
16.2795944213867,-51.5754699707031,
43.6027717590332,-35.2556114196777,
20.6249198913574,-10.1874380111694,
-27.4139785766602,8.92145633697510,
-55.6165428161621,12.1048450469971,
-40.4292297363281,10.8523015975952,
1.96676838397980,21.2064609527588,
29.8661289215088,30.9156188964844,
22.0365314483643,7.75531291961670,
-1.05109786987305,-44.9531059265137,
-3.85012531280518,-70.5662841796875,
23.8466415405273,-30.6577835083008,
45.8859481811523,32.8628692626953,
21.4841747283936,44.7489662170410,
-35.7938575744629,-6.27628755569458,
-57.7443656921387,-52.6697463989258,
-5.80189132690430,-41.1537437438965,
70.9585418701172,-0.460423231124878,
82.2029037475586,9.65746688842773,
17.1850643157959,-4.25113773345947,
-38.5162849426270,0.296088576316834,
-18.2393798828125,22.6194438934326,
41.9063301086426,18.5553340911865,
53.6252746582031,-11.5301189422607,
1.80525445938110,-16.8331489562988,
-41.2932281494141,20.6120853424072,
-30.1464080810547,41.5499572753906,
-2.93845486640930,3.34151625633240,
-13.5521039962769,-44.6552276611328,
-45.5469360351563,-31.1663379669189,
-51.9686050415039,28.1647148132324,
-30.1360168457031,49.0947341918945,
-22.4094276428223,5.65407562255859,
-37.7452507019043,-31.6524257659912,
-38.0387649536133,-12.0115165710449,
-9.67703533172607,23.2431240081787,
9.19138240814209,20.0095367431641,
-12.0123815536499,-3.37717247009277,
-48.5574493408203,6.19011068344116,
-53.2360458374023,45.9337387084961,
-23.4656600952148,63.9813003540039,
1.34906268119812,42.2117004394531,
9.44123554229736,18.3207378387451,
20.3912010192871,19.8402576446533,
40.7086143493652,26.8660392761230,
52.2512702941895,11.5448942184448,
42.1663513183594,-6.74298429489136,
23.5132350921631,3.91711950302124,
9.16674137115479,33.7565650939941,
-2.30459737777710,45.0161666870117,
-17.0678215026855,28.0145759582520,
-20.7230854034424,6.90005397796631,
-3.21784830093384,0.427055805921555,
18.9859046936035,5.64428234100342,
21.0495338439941,9.48525142669678,
10.0395765304565,7.65856695175171,
15.5960159301758,7.25179147720337,
38.2380371093750,13.4775438308716,
45.2932014465332,22.9947910308838,
21.1955261230469,33.0980796813965,
-8.22318553924561,39.3002471923828,
-11.4935741424561,37.2101058959961,
1.72066104412079,30.1245841979980,
-0.307138293981552,27.0077247619629,
-21.7534980773926,22.5892543792725,
-32.8399162292481,1.27826619148254,
-20.4616661071777,-34.8088798522949,
-7.41707944869995,-62.5727310180664,
-20.8069820404053,-64.1334838867188,
-48.4837608337402,-48.1976890563965,
-56.5933341979981,-40.4335136413574,
-38.2908706665039,-39.5469512939453,
-22.1256351470947,-23.2869606018066,
-27.0578136444092,17.1062526702881,
-36.9981994628906,55.9442138671875,
-26.0290374755859,60.2140998840332,
1.85810291767120,33.6182746887207,
14.3841896057129,10.5738792419434,
-7.78446292877197,12.1940536499023,
-37.8012504577637,18.1256828308105,
-36.6525764465332,-0.464617013931274,
0.524438381195068,-40.0201530456543,
37.0215110778809,-60.5926628112793,
41.7916069030762,-33.2741317749023,
18.7382907867432,22.0193424224854,
-3.94243955612183,51.7798309326172,
-14.9605302810669,26.5663757324219,
-24.1902198791504,-23.4713478088379,
-35.3542137145996,-46.4762878417969,
-29.1859207153320,-21.9168090820313,
0.877126574516296,19.0554904937744,
31.1445808410645,36.4588928222656,
29.7793502807617,21.8337154388428,
-2.76177930831909,3.91164183616638,
-31.7141265869141,4.00821971893311,
-32.9482460021973,10.1177577972412,
-18.3526325225830,4.35487556457520,
-16.3991832733154,-11.8156948089600,
-27.5996036529541,-17.7514305114746,
-29.7279834747314,0.409777134656906,
-11.9911670684814,27.7596073150635,
7.96855497360230,38.8002738952637,
4.86504602432251,31.7654323577881,
-19.9868659973145,20.1507530212402,
-41.8402900695801,7.46121549606323,
-43.9570541381836,-10.4387245178223,
-31.9629001617432,-25.5954170227051,
-23.3659458160400,-12.6260490417480,
-24.0744190216064,32.0909080505371,
-31.6728591918945,65.4671859741211,
-41.7758102416992,40.3530158996582,
-51.7179489135742,-26.6347236633301,
-52.0020446777344,-65.6768951416016,
-34.8975105285645,-32.5930786132813,
-6.79025268554688,31.6997985839844,
12.5693273544312,55.8630905151367,
9.20018196105957,26.5724296569824,
-8.82538414001465,-11.0014963150024,
-25.5059814453125,-19.8006019592285,
-25.7471160888672,-7.21567964553833,
-8.19264793395996,2.39796209335327,
20.1397819519043,-3.59830379486084,
42.9980964660645,-21.7902889251709,
45.1360054016113,-44.7478370666504,
22.5709571838379,-57.3915176391602,
3.51556015014648,-38.9113502502441,
12.7398242950439,-2.35643863677979,
42.0777854919434,10.3481245040894,
56.6288566589356,-19.9431648254395,
42.0082054138184,-52.1331291198731,
17.8517456054688,-31.3855686187744,
5.93538093566895,25.6813354492188,
-3.11511540412903,49.7713890075684,
-27.9381217956543,14.3765792846680,
-54.5317382812500,-28.8350296020508,
-52.4227066040039,-22.1990985870361,
-26.1286087036133,15.9638681411743,
-19.8852615356445,21.5876235961914,
-50.1981849670410,-24.0271072387695,
-73.8881225585938,-70.3771743774414,
-48.1209564208984,-64.3571090698242,
8.48327159881592,-15.2757930755615,
34.5086669921875,29.8594551086426,
13.6286315917969,41.2500267028809,
-12.1789455413818,28.2243423461914,
-2.71947789192200,13.9654541015625,
22.4847431182861,9.92184925079346,
25.9639186859131,10.6369190216064,
3.00522756576538,6.07126045227051,
-15.5883617401123,-6.35552406311035,
-20.5145759582520,-9.62901973724365,
-21.8135814666748,4.54939222335815,
-18.9732532501221,23.5599822998047,
0.993822097778320,21.2767181396484,
32.3583717346191,-7.43809795379639,
49.5312805175781,-35.4643096923828,
44.2184638977051,-33.3918762207031,
38.8361511230469,-7.73226165771484,
43.8851852416992,6.33435249328613,
37.9392929077148,-6.98941278457642,
-1.63970243930817,-29.9181003570557,
-48.3903846740723,-36.6863822937012,
-56.4436683654785,-20.1466102600098,
-34.3444747924805,3.66122627258301,
-28.5852699279785,20.4751033782959,
-51.4234428405762,24.8780364990234,
-58.6237449645996,22.4073390960693,
-17.1150093078613,21.2856101989746,
41.3025016784668,27.2922039031982,
61.8747863769531,32.8080825805664,
40.9604606628418,23.0257873535156,
19.9965229034424,1.09881150722504,
18.8838958740234,-10.8226737976074,
22.3814449310303,8.35495948791504,
18.1292266845703,46.4989166259766,
23.1503009796143,63.6926116943359,
40.7754821777344,39.8434028625488,
40.7680320739746,-1.85115957260132,
-1.83753967285156,-25.7904396057129,
-55.7194938659668,-21.1448364257813,
-64.5638427734375,-6.99096488952637,
-20.7812232971191,-6.44263076782227,
27.2613925933838,-19.7929286956787,
34.3286743164063,-29.2386493682861,
8.92249584197998,-22.8613071441650,
-4.04479312896729,0.590409159660339,
17.1681041717529,30.7846813201904,
43.4589157104492,46.5357818603516,
43.8611984252930,33.4734153747559,
16.7162551879883,4.88733100891113,
-7.77927684783936,-5.86752033233643,
-11.6432552337646,14.0468225479126,
-7.29307317733765,37.3660469055176,
-15.1001482009888,23.6196193695068,
-28.7716159820557,-20.1392688751221,
-26.2226371765137,-44.8220977783203,
-1.05720341205597,-22.2167606353760,
13.8321971893311,9.14379501342773,
-7.61345911026001,-1.88467383384705,
-47.5708084106445,-41.0351943969727,
-62.8041000366211,-46.4908256530762,
-34.6220741271973,-3.09029722213745,
12.9954566955566,29.5067043304443,
44.7334938049316,2.34246540069580,
48.3223609924316,-44.7092781066895,
33.3665504455566,-34.9539642333984,
10.1533813476563,28.0895767211914,
-8.36423778533936,65.8882522583008,
-11.3755655288696,35.8046951293945,
4.66890144348145,-10.0022106170654,
19.0991821289063,-3.57119727134705,
8.07132053375244,41.7128829956055,
-23.2950801849365,54.9517211914063,
-47.8637504577637,14.7090053558350,
-50.4313163757324,-27.3612117767334,
-42.4178886413574,-29.1532993316650,
-37.8902664184570,-8.01379299163818,
-28.5011329650879,-4.18757104873657,
-4.98093223571777,-19.2437477111816,
17.5050601959229,-21.9938507080078,
17.6112594604492,-0.126964807510376,
-0.332336425781250,21.1805610656738,
0.239110589027405,17.7561359405518,
31.3752079010010,-2.82806563377380,
63.2121047973633,-16.8775959014893,
55.7731704711914,-13.7717590332031,
13.3044862747192,1.37064540386200,
-15.7355365753174,10.8573760986328,
-2.07704234123230,4.16584444046021,
29.5587406158447,-9.58634471893311,
36.6452140808106,-13.4436922073364,
8.10230541229248,-3.44966983795166,
-23.4998512268066,9.46280574798584,
-30.2438030242920,9.51392364501953,
-20.2202053070068,-4.83145570755005,
-12.2519826889038,-16.2206993103027,
-6.51836013793945,-14.5489673614502,
9.40831375122070,-5.09104537963867,
34.7304000854492,5.25747203826904,
46.3982849121094,16.7173500061035,
25.6429347991943,29.0970973968506,
-13.3898639678955,31.2613925933838,
-39.6590156555176,9.31353759765625,
-31.7417945861816,-27.7484817504883,
6.14951896667481,-45.6653404235840,
47.8644180297852,-20.2727699279785,
58.0382614135742,31.2978153228760,
19.0336818695068,66.4717407226563,
-38.7325096130371,58.9198913574219,
-59.5659751892090,26.6166191101074,
-29.8778591156006,10.5203714370728,
1.63702821731567,23.0373172760010,
-15.0259590148926,30.1895847320557,
-60.3892211914063,2.89880967140198,
-62.0602951049805,-38.5190925598145,
-1.59362125396729,-49.1879081726074,
52.0825614929199,-13.2113380432129,
34.8000411987305,25.0068340301514,
-24.5007915496826,20.8694915771484,
-53.0198936462402,-8.21066665649414,
-33.4904365539551,-11.5523605346680,
-13.0773925781250,17.8092041015625,
-21.0462112426758,34.9469490051270,
-30.9205398559570,15.5562171936035,
-17.6613273620605,-7.68922853469849,
-7.22119188308716,5.28727149963379,
-23.0593547821045,36.4134750366211,
-39.4871292114258,25.6560516357422,
-17.0890235900879,-27.9366741180420,
30.1054763793945,-51.7523612976074,
43.6637344360352,3.00442242622376,
9.25452232360840,84.0356063842773,
-24.0517635345459,94.4726333618164,
-14.5612182617188,20.0997085571289,
17.0519065856934,-54.2000999450684,
33.8862876892090,-50.1347885131836,
27.2021141052246,2.84964299201965,
14.8829584121704,23.6840324401855,
10.4786291122437,-5.78307771682739,
10.8098402023315,-23.2808895111084,
15.7435455322266,7.54619073867798,
24.1365661621094,41.5737228393555,
24.1418399810791,23.8426475524902,
6.19863557815552,-24.4548435211182,
-12.8114604949951,-35.1118011474609,
-6.39098978042603,5.53164243698120,
16.8434181213379,42.7700920104981,
20.2566890716553,40.4385375976563,
-1.53772854804993,27.3913745880127,
-15.9985446929932,37.5428733825684,
-1.87189567089081,52.9128456115723,
18.2379856109619,39.9825553894043,
14.1727905273438,14.0485115051270,
-5.80802726745606,17.4011306762695,
-12.4935321807861,43.2919044494629,
-2.39812564849854,43.1606712341309,
3.95168876647949,1.37335836887360,
2.51087117195129,-40.1728591918945,
14.8651094436646,-44.3045501708984,
45.4300613403320,-30.4361667633057,
62.0415954589844,-31.3021392822266,
42.9509849548340,-41.5026016235352,
13.6517696380615,-36.1802902221680,
10.6252021789551,-19.3506622314453,
33.0462265014648,-17.5573444366455,
50.5636825561523,-26.9490909576416,
43.2943496704102,-7.11252880096436,
18.8018665313721,43.0472221374512,
-9.09687900543213,73.7799377441406,
-31.3574085235596,45.2161865234375,
-35.4536666870117,-12.3864507675171,
-13.6860704421997,-38.7709770202637,
13.5262422561646,-9.74828338623047,
8.36786556243897,38.9271125793457,
-29.4082050323486,53.4427757263184,
-54.0644454956055,21.5719223022461,
-32.0466117858887,-22.2635803222656,
4.48008441925049,-39.7236709594727,
2.24027681350708,-16.4877109527588,
-34.2221946716309,17.3830547332764,
-49.5270195007324,17.1626167297363,
-12.4479875564575,-30.9341068267822,
36.4213409423828,-76.4094619750977,
43.8619461059570,-66.6812896728516,
10.6464004516602,-17.7456302642822,
-16.3609924316406,4.97510290145874,
-11.7658538818359,-23.8717422485352,
3.00989174842834,-53.9879302978516,
-3.06311035156250,-32.0333290100098,
-24.4230918884277,20.9673614501953,
-37.8367500305176,32.5499534606934,
-39.0549392700195,-11.6620988845825,
-38.3504066467285,-49.9539756774902,
-37.4524803161621,-40.1131477355957,
-24.4285659790039,-11.3512134552002,
13.7897558212280,-0.523253321647644,
55.8229751586914,7.56113338470459,
60.4979782104492,40.5085563659668,
17.0909881591797,66.1732406616211,
-27.9626140594482,35.2202377319336,
-24.3696174621582,-30.8773021697998,
22.6502513885498,-51.0516586303711,
50.6599655151367,-4.54693412780762,
18.1696434020996,34.1718978881836,
-34.4710578918457,4.16767024993897,
-35.4978942871094,-48.7810440063477,
19.5261669158936,-47.3347396850586,
56.8692588806152,-4.44165706634522,
25.0042934417725,7.25893020629883,
-38.0359230041504,-25.1723880767822,
-59.5533599853516,-43.4965400695801,
-29.4527435302734,-21.4529094696045,
1.62891519069672,-6.43268632888794,
-2.65477490425110,-31.5731201171875,
-16.6504325866699,-55.3576889038086,
-3.31439614295959,-28.2984714508057,
24.0170269012451,15.5311155319214,
31.5938911437988,10.5572490692139,
17.8677444458008,-38.4355392456055,
8.63946342468262,-56.9784088134766,
12.1517410278320,-17.4444980621338,
6.90695858001709,19.1392650604248,
-15.1936368942261,-0.548951625823975,
-23.6794681549072,-41.0333404541016,
3.26527857780457,-44.2377700805664,
36.9836769104004,-1.83667159080505,
32.9265098571777,41.4488449096680,
-7.52586412429810,54.5516662597656,
-37.0898780822754,48.8442382812500,
-22.8415431976318,47.0243492126465,
7.86418008804321,42.8593101501465,
13.4855384826660,25.7420330047607,
-4.28626680374146,0.127480924129486,
-9.95445823669434,-17.9915390014648,
9.87365341186523,-21.8232498168945,
26.6718330383301,-10.5438861846924,
19.8007793426514,6.20703315734863,
0.0988909006118774,3.76594877243042,
-3.11065673828125,-31.3539142608643,
9.62059307098389,-73.5425109863281,
13.5558938980103,-76.0326080322266,
-2.46874427795410,-29.8610534667969,
-21.4215068817139,17.6605415344238,
-22.7523803710938,14.9167890548706,
-13.0416584014893,-28.5793743133545,
-6.06705999374390,-55.9444465637207,
-7.10106134414673,-41.4952888488770,
-4.12062501907349,-12.0698051452637,
13.5912876129150,-2.63567399978638,
40.0244522094727,-3.32335233688355,
51.5759963989258,10.9143314361572,
31.7167778015137,35.3637123107910,
-14.7679738998413,35.9980812072754,
-58.2182235717773,1.49861049652100,
-67.6894912719727,-39.1655006408691,
-38.8294219970703,-50.5805282592773,
-2.86711430549622,-33.6379241943359,
9.18447589874268,-14.0683765411377,
6.87534570693970,-7.85515594482422,
19.0411891937256,-9.63606929779053,
47.0696487426758,-3.83968830108643,
64.1728973388672,8.21722984313965,
52.7510375976563,13.4343767166138,
32.9942321777344,9.83347606658936,
35.5524368286133,2.85312795639038,
50.4894027709961,7.67247438430786,
43.9979248046875,26.0219993591309,
7.71452140808106,41.4833984375000,
-26.7490482330322,35.5954895019531,
-38.2738838195801,8.79404830932617,
-34.1475944519043,-21.3754062652588,
-23.8351745605469,-38.5806694030762,
0.214086920022964,-40.2568969726563,
38.7797622680664,-27.3744201660156,
54.3508605957031,-4.74450683593750,
20.2377376556397,21.4045333862305,
-33.4984512329102,28.5032653808594,
-43.1011314392090,-1.04962790012360,
5.57369899749756,-51.0036163330078,
58.6252059936523,-76.7048797607422,
63.5691528320313,-53.9194602966309,
39.4802398681641,-8.25713443756104,
28.1315155029297,15.9566612243652,
31.8968811035156,4.66527271270752,
18.5687122344971,-21.1782417297363,
-13.1195011138916,-36.3711509704590,
-30.2222232818604,-36.3502731323242,
-19.0797309875488,-22.2327251434326,
1.35399258136749,9.78427219390869,
9.34541988372803,51.1359100341797,
14.4912738800049,69.8139801025391,
27.0737342834473,45.4541969299316,
31.9472332000732,2.71726799011230,
13.8758668899536,-13.7518720626831,
-6.80199337005615,3.54695868492126,
0.663028597831726,14.4373083114624,
26.5074939727783,-7.56599092483521,
36.6259994506836,-30.0738162994385,
25.0647144317627,-16.4825801849365,
8.58858585357666,20.1337242126465,
-7.07585048675537,27.2662200927734,
-32.5106086730957,-10.0796251296997,
-58.7139244079590,-43.3362503051758,
-55.3592681884766,-25.5293197631836,
-17.6501979827881,19.4756603240967,
13.2839412689209,30.4287185668945,
3.60153007507324,-10.8143081665039,
-16.4259490966797,-58.8935661315918,
-0.0623939037322998,-60.6781234741211,
40.9301528930664,-16.9670906066895,
50.0143928527832,26.8440761566162,
16.8160076141357,29.0120525360107,
-9.01278972625732,-5.82955121994019,
1.45877742767334,-36.2507247924805,
15.2203540802002,-32.4438362121582,
-5.60610103607178,-3.20415067672730,
-38.8162422180176,12.9840106964111,
-38.5315055847168,-8.22912597656250,
-6.93360090255737,-36.1599769592285,
6.67390680313110,-22.4104328155518,
-11.6587686538696,33.2421188354492,
-25.8823394775391,71.1623001098633,
-5.93200254440308,53.9053077697754,
25.7615814208984,11.6016855239868,
36.8718376159668,-2.30304455757141,
35.9182472229004,17.2796974182129,
45.4756011962891,27.9101562500000,
54.6744461059570,7.84352636337280,
39.2837028503418,-2.08630824089050,
1.49519371986389,26.9191627502441,
-30.5923423767090,54.5850639343262,
-39.4750061035156,30.1238803863525,
-39.0187568664551,-28.0685729980469,
-48.4092941284180,-57.6933746337891,
-59.1927375793457,-46.0555343627930,
-53.6339836120606,-37.7864379882813,
-28.7790870666504,-54.7207984924316,
7.02154350280762,-56.2882461547852,
41.0845375061035,-12.6907482147217,
57.3190536499023,37.1042060852051,
42.9392547607422,43.0225601196289,
15.5990009307861,22.2726631164551,
11.8603734970093,33.0811882019043,
39.1238479614258,63.0220489501953,
61.3964805603027,49.3022460937500,
40.8679580688477,-11.4754657745361,
-2.86111307144165,-40.7611198425293,
-18.8221092224121,2.50187611579895,
12.0492277145386,49.0841217041016,
51.3231658935547,25.9319496154785,
56.4542961120606,-35.6067733764648,
32.0949707031250,-46.0915145874023,
8.89346885681152,0.500574111938477,
-9.59152603149414,23.3273239135742,
-26.3374958038330,-9.09674835205078,
-31.8494262695313,-33.2896690368652,
-16.0834999084473,4.55010128021240,
7.64951753616333,52.6583938598633,
12.2831954956055,31.1637401580811,
-2.28271317481995,-40.3439254760742,
-12.8989086151123,-73.5753860473633,
-9.65261268615723,-33.8541755676270,
-13.3031816482544,22.2032699584961,
-22.3376159667969,38.1674041748047,
-5.68280410766602,22.5772647857666,
47.8739204406738,24.1239681243897,
80.2704086303711,52.4831619262695,
33.6583061218262,71.1790924072266,
-51.7127990722656,50.6687316894531,
-77.1886672973633,8.49927711486816,
-15.2765560150146,-21.0928115844727,
48.1026535034180,-13.8183422088623,
29.5515670776367,21.1767826080322,
-36.4065666198731,45.9114875793457,
-48.4932746887207,32.6143493652344,
13.0552024841309,-1.93377661705017,
64.4603271484375,-14.1420774459839,
39.7376251220703,5.48771524429321,
-24.3678569793701,20.4661788940430,
-56.3547325134277,-0.720452129840851,
-45.9991035461426,-42.2101211547852,
-30.2481594085693,-56.7298126220703,
-24.0320301055908,-35.5261497497559,
-11.4927110671997,-19.7594108581543,
2.18667411804199,-39.1672096252441,
-3.52250576019287,-66.6196975708008,
-24.8405838012695,-58.3422012329102,
-24.0579986572266,-15.6805114746094,
19.0076503753662,20.8454151153564,
64.4799804687500,27.2180538177490,
66.2849960327148,17.1932888031006,
36.0640220642090,12.2347860336304,
11.3121528625488,13.8368949890137,
1.84979367256165,14.9682950973511,
-4.12543916702271,13.1744651794434,
-6.15893650054932,11.5740928649902,
0.150339603424072,9.31354999542236,
9.32575416564941,8.53579044342041,
8.73652362823486,17.5880298614502,
5.37246894836426,30.9557151794434,
21.2592468261719,22.6377296447754,
42.4030380249023,-18.0008964538574,
30.7881107330322,-56.6085815429688,
-16.3800849914551,-46.3921546936035,
-41.4447517395020,4.49898242950439,
-6.62232112884522,35.9687995910645,
44.7744979858398,14.3428859710693,
51.0583457946777,-23.3146648406982,
18.5454635620117,-21.0826187133789,
0.588660299777985,19.8497295379639,
12.4201984405518,44.2092514038086,
9.21033573150635,24.7096691131592,
-33.0578536987305,-3.99592661857605,
-69.3201065063477,-1.10419344902039,
-50.4308357238770,21.1589527130127,
0.684423446655273,19.2790412902832,
27.1782474517822,-17.8201961517334,
19.9556732177734,-57.8123092651367,
22.3055667877197,-58.7793045043945,
46.4115638732910,-17.8478450775147,
51.4982070922852,32.5149307250977,
9.87314510345459,51.2772979736328,
-41.8582763671875,26.0050964355469,
-54.7704124450684,-23.0222625732422,
-28.9749069213867,-58.7745056152344,
-5.60598659515381,-56.7439041137695,
-11.6836910247803,-31.9235439300537,
-28.5929145812988,-14.9305076599121,
-34.5011711120606,-10.9688367843628,
-31.1174736022949,2.05583310127258,
-32.1174163818359,25.1127452850342,
-38.0925025939941,26.7752475738525,
-39.1154251098633,-12.8792171478271,
-37.8032798767090,-59.9423294067383,
-33.3671188354492,-61.6577110290527,
-23.9756374359131,-15.4406147003174,
-15.8704948425293,20.1234226226807,
-18.5431461334229,4.47907304763794,
-28.3448429107666,-28.9316120147705,
-26.9836273193359,-26.1023445129395,
-7.34962415695190,15.1608581542969,
19.5131950378418,45.7149162292481,
33.5591354370117,36.3164062500000,
35.4011688232422,12.3930473327637,
35.2835464477539,3.15627527236938,
22.8754844665527,10.3172721862793,
-15.5660448074341,20.4786357879639,
-56.7248306274414,31.0690670013428,
-59.5670547485352,43.6844787597656,
-19.1737194061279,42.0946998596191,
15.4607887268066,12.3042945861816,
10.6432590484619,-28.7121391296387,
-9.24669742584229,-44.3829689025879,
-0.0631251931190491,-26.2599887847900,
26.5304660797119,-2.53410601615906,
21.3778915405273,3.91621351242065,
-23.7178268432617,0.390692591667175,
-49.7513580322266,-5.22488021850586,
-13.3623542785645,-15.2057428359985,
47.0811195373535,-23.2927665710449,
61.0686187744141,-13.4390716552734,
17.5137462615967,21.0781898498535,
-26.7414970397949,51.2087745666504,
-23.8194026947022,41.3645706176758,
9.71505451202393,0.0509522147476673,
32.4597473144531,-27.0110969543457,
32.4346847534180,-24.0184230804443,
22.3553581237793,-16.0043106079102,
15.3677635192871,-24.3946437835693,
9.02899074554443,-35.5824928283691,
2.52889466285706,-36.8350639343262,
6.98975753784180,-36.7988128662109,
25.9381561279297,-41.4976692199707,
38.5388526916504,-29.0755062103272,
25.3715686798096,17.2041435241699,
-11.0675086975098,59.7250938415527,
-43.2096939086914,44.4735984802246,
-42.2439880371094,-14.6092376708984,
-9.08528614044190,-42.0279502868652,
20.9693908691406,1.06361627578735,
17.6051349639893,55.1205329895020,
-10.3636322021484,44.5229339599609,
-27.3829135894775,-12.8039398193359,
-14.3245468139648,-44.5903015136719,
6.57104730606079,-27.8371200561523,
3.70191812515259,-11.6575622558594,
-18.1895465850830,-34.5298652648926,
-22.6730613708496,-65.2197341918945,
10.7166042327881,-54.7769012451172,
55.5598411560059,-9.79201412200928,
69.8914489746094,22.9274196624756,
47.5707893371582,23.1577167510986,
13.3167934417725,4.09878206253052,
-10.9722118377686,-18.8975334167480,
-20.4831695556641,-40.6944427490234,
-20.2912788391113,-41.5343742370606,
-9.86584663391113,-5.87200403213501,
0.585101842880249,39.2965850830078,
-5.35027456283569,53.9495315551758,
-29.9621009826660,35.9278717041016,
-47.5381393432617,24.0857429504395,
-36.7719879150391,36.3412284851074,
-10.8045835494995,42.2251701354981,
-1.91288042068481,9.14050292968750,
-10.7481842041016,-36.8345489501953,
-5.20903873443604,-44.5752716064453,
27.5134792327881,-16.3727741241455,
54.3379859924316,1.52435982227325,
38.2687225341797,-2.88147115707397,
-5.15049600601196,-3.20949292182922,
-29.9796161651611,8.06466293334961,
-24.6206684112549,3.30672264099121,
-20.0853519439697,-29.6494235992432,
-37.1391448974609,-59.1438484191895,
-51.7017326354981,-56.4446372985840,
-38.8724822998047,-44.5986976623535,
-13.9917755126953,-51.0334930419922,
-7.72323656082153,-54.9066276550293,
-14.0556688308716,-15.9429330825806,
-1.34572625160217,41.5359764099121,
29.1234703063965,48.6498031616211,
38.0121231079102,-6.64800643920898,
6.45429182052612,-50.4296951293945,
-35.1893920898438,-26.3534545898438,
-41.0726470947266,22.1503009796143,
-10.8116264343262,21.4724407196045,
19.9041748046875,-21.2139148712158,
32.4506187438965,-32.6274948120117,
38.6155700683594,18.5979156494141,
42.6390609741211,78.9451980590820,
39.8897590637207,82.0638427734375,
28.3684120178223,36.7705345153809,
20.9848594665527,1.77844452857971,
20.9674339294434,-0.947356283664703,
24.1247005462647,3.87726116180420,
28.3070011138916,-11.5979795455933,
36.2144889831543,-32.0128974914551,
36.7468681335449,-29.7108764648438,
5.08077669143677,-1.97254312038422,
-53.1886634826660,23.6762466430664,
-83.5394897460938,15.5255165100098,
-40.8775825500488,-24.2424297332764,
33.0335617065430,-55.6988334655762,
54.0822296142578,-43.9906082153320,
3.85134744644165,5.02214336395264,
-54.2575836181641,50.0378265380859,
-58.4156417846680,56.8701057434082,
-29.4541950225830,27.7042007446289,
-18.5464591979980,-4.95071792602539,
-27.3464107513428,-26.9740638732910,
-13.3976001739502,-37.8726577758789,
26.7404937744141,-36.8032493591309,
49.6855125427246,-15.7068109512329,
31.9451675415039,21.9473495483398,
11.0213003158569,50.8752365112305,
15.8135566711426,50.0314140319824,
19.5976543426514,27.0049514770508,
-13.0898303985596,3.38490867614746,
-55.9470939636231,-4.36689090728760,
-49.9118957519531,-0.186471343040466,
8.20227336883545,7.88152599334717,
57.9597091674805,19.7931137084961,
55.7128295898438,30.6737403869629,
19.6799468994141,38.2766799926758,
-1.25751066207886,41.6146507263184,
2.43362522125244,41.9973106384277,
14.3121623992920,31.5217342376709,
27.7114238739014,2.87963700294495,
42.3924560546875,-27.8100490570068,
44.7461013793945,-25.8478546142578,
21.4067153930664,24.2444534301758,
-9.66509342193604,79.6433639526367,
-18.7933921813965,81.1299667358398,
-4.82448053359985,19.4372100830078,
-1.45682728290558,-47.0695457458496,
-22.8081569671631,-51.2273483276367,
-46.8313636779785,2.14161133766174,
-48.0733299255371,52.3662643432617,
-35.8712654113770,54.8328247070313,
-37.6301574707031,22.7644481658936,
-50.5137596130371,-2.28674507141113,
-41.2486419677734,-4.71919393539429,
-1.61936950683594,4.09142255783081,
37.4212112426758,9.65864753723145,
41.5828323364258,7.78916120529175,
11.5403404235840,-9.08042335510254,
-18.5257205963135,-41.4097099304199,
-16.2611007690430,-67.3913116455078,
19.4477119445801,-56.5734786987305,
53.4794731140137,-8.63998985290527,
51.5995445251465,33.1743927001953,
13.5295162200928,25.7938289642334,
-26.7589874267578,-15.2527933120728,
-34.4070434570313,-40.8156585693359,
-14.8927698135376,-24.9963016510010,
-4.42007732391357,13.4906187057495,
-21.3379573822022,37.3116798400879,
-36.8611717224121,32.3190612792969,
-20.8303012847900,13.2611722946167,
12.8419561386108,-0.168586328625679,
17.1628932952881,3.09311866760254,
-13.3459739685059,20.4867515563965,
-38.6590385437012,29.6010475158691,
-23.1995792388916,6.67029237747192,
14.5717220306396,-34.3207435607910,
27.6193828582764,-45.9055747985840,
4.00215435028076,-9.58871650695801,
-22.8282318115234,24.7144298553467,
-27.5476760864258,4.58720922470093,
-15.8655843734741,-48.8586273193359,
-7.29461765289307,-67.5726318359375,
-5.25742292404175,-23.5429420471191,
-5.40514802932739,29.0215110778809,
-7.68814706802368,34.8219604492188,
-3.66630411148071,15.7427768707275,
19.6775112152100,18.5014877319336,
54.8075561523438,29.2067356109619,
64.0188598632813,8.23996353149414,
28.5670509338379,-26.6645336151123,
-21.7825660705566,-20.3658676147461,
-34.1233749389648,27.1519241333008,
2.06542181968689,49.7564086914063,
36.5540237426758,17.5546436309814,
30.1611003875732,-9.28896427154541,
-0.253742098808289,19.5389995574951,
-22.7624053955078,61.4639968872070,
-34.7029304504395,42.4359741210938,
-42.3931350708008,-18.8240947723389,
-37.0714225769043,-36.9432182312012,
-11.7412538528442,4.65538692474365,
13.2594881057739,28.1348419189453,
11.6667032241821,-8.31528186798096,
-2.51216030120850,-42.0877456665039,
11.7281179428101,-10.5750436782837,
47.0948867797852,46.8988189697266,
45.1231155395508,46.7710876464844,
-10.7722587585449,-9.30483245849609,
-56.3202514648438,-49.2675056457520,
-33.0315513610840,-35.5288467407227,
19.0681610107422,-13.9446229934692,
21.5084743499756,-28.5694770812988,
-23.2878227233887,-49.1403503417969,
-43.0156059265137,-27.2978744506836,
-12.1016969680786,22.9225330352783,
9.47117805480957,45.4737052917481,
-26.4344520568848,22.5558052062988,
-68.1065292358398,-10.4976119995117,
-41.2929878234863,-20.9431877136230,
29.9204597473145,-6.18692398071289,
56.9669990539551,9.68091773986816,
17.1841392517090,7.38476228713989,
-22.4824275970459,-15.0428905487061,
-14.0608549118042,-42.4781608581543,
8.66866970062256,-56.7085189819336,
2.09238386154175,-45.6329574584961,
-12.4618949890137,-19.0865364074707,
-0.816018581390381,-0.684135079383850,
16.0355300903320,0.583938360214233,
-6.40492486953735,-11.0144433975220,
-49.6009178161621,-25.5631179809570,
-46.8112258911133,-38.3481254577637,
13.9031276702881,-37.7419776916504,
56.0966987609863,-9.73775196075440,
21.1111412048340,33.8987770080566,
-47.2575759887695,63.3276290893555,
-60.1583251953125,57.6536941528320,
-8.14557552337647,28.6783866882324,
38.8358917236328,6.11078739166260,
25.6632099151611,5.94732904434204,
-22.1989898681641,19.8174858093262,
-43.8549652099609,29.7215843200684,
-22.1821517944336,22.1442337036133,
4.57921123504639,-3.07819223403931,
1.58126568794250,-35.6900634765625,
-20.5153350830078,-47.3095817565918,
-26.7406539916992,-20.3613834381104,
-8.69391632080078,30.7736167907715,
10.5472927093506,65.3768997192383,
5.95835304260254,53.6558074951172,
-23.2086143493652,7.98228645324707,
-49.7189483642578,-33.3408660888672,
-48.9135208129883,-48.0924224853516,
-25.7364044189453,-43.0735664367676,
3.38685250282288,-32.1331138610840,
28.9037570953369,-20.9616355895996,
43.2443389892578,-1.29251480102539,
37.2577857971191,20.1784515380859,
12.5447540283203,22.1472148895264,
-13.1484632492065,-7.21298456192017,
-11.0881252288818,-48.2742500305176,
23.2825260162354,-67.4132766723633,
54.3120117187500,-43.3704795837402,
43.2127532958984,7.69583034515381,
2.45329046249390,47.9567565917969,
-19.6789627075195,52.4214859008789,
-0.190777182579041,27.6491985321045,
26.3415241241455,1.02033460140228,
15.0064830780029,-8.41640853881836,
-25.6542434692383,-6.01573133468628,
-43.8289375305176,-11.9478683471680,
-22.0529575347900,-32.5716361999512,
-0.932512044906616,-41.1480484008789,
-16.9231319427490,-19.0579242706299,
-47.8208465576172,12.4570045471191,
-43.9754600524902,7.44284439086914,
-5.42407894134522,-37.0491409301758,
17.4890403747559,-66.7172393798828,
-8.23827934265137,-34.4154090881348,
-45.5793876647949,34.3601989746094,
-41.8432693481445,57.8585777282715,
-3.63851451873779,9.22001171112061,
21.3847293853760,-50.7864494323731,
8.21215057373047,-59.6894607543945,
-18.0724353790283,-21.4509277343750,
-18.7187194824219,15.1466636657715,
0.854665994644165,29.2536468505859,
0.653922796249390,38.6855735778809,
-30.5854816436768,45.6268539428711,
-57.4870300292969,33.2598152160645,
-44.2719383239746,7.26849937438965,
-0.816054105758667,7.03700733184814,
22.7597599029541,39.5925598144531,
-4.66890811920166,51.4142837524414,
-48.8775100708008,4.31547880172730,
-49.3029747009277,-57.8826942443848,
2.32575893402100,-55.7220230102539,
44.0299987792969,11.4527769088745,
20.6099681854248,62.1205139160156,
-45.7737236022949,40.0285568237305,
-74.3897628784180,-20.9663162231445,
-26.7070255279541,-59.0906448364258,
42.5632324218750,-55.4084625244141,
55.6440849304199,-36.2793464660645,
6.33733510971069,-16.4144134521484,
-37.8289146423340,11.1169824600220,
-32.0703048706055,33.1072654724121,
-6.75868320465088,23.3359127044678,
-10.1845388412476,-16.2351970672607,
-42.7893524169922,-44.5202407836914,
-59.3353118896484,-42.7541923522949,
-37.8915405273438,-32.1620903015137,
-7.39470577239990,-33.3696289062500,
0.560064077377319,-37.7761268615723,
-8.05218315124512,-40.6364364624023,
-14.0200386047363,-46.0492172241211,
-8.79918193817139,-51.7906913757324,
4.36268424987793,-42.2866210937500,
30.0588703155518,-6.45100164413452,
59.5937995910645,30.5781440734863,
56.6131439208984,38.0609588623047,
4.73651885986328,35.5997543334961,
-48.5543785095215,50.3549842834473,
-44.9449157714844,60.9358901977539,
5.76421594619751,21.6144065856934,
34.6969108581543,-46.1983108520508,
3.48378229141235,-63.4372825622559,
-37.9022560119629,-5.93016481399536,
-25.5756034851074,44.4381980895996,
24.5017490386963,14.5730304718018,
50.5813331604004,-49.6699104309082,
43.2859954833984,-47.2926406860352,
39.7872810363770,28.9979476928711,
53.7266387939453,75.5065002441406,
52.8383941650391,30.2798156738281,
23.5734252929688,-45.7992591857910,
2.31680750846863,-61.5674934387207,
13.3176784515381,-22.1082267761230,
20.1954059600830,-3.04059767723084,
-10.0842494964600,-26.0109939575195,
-47.8808250427246,-41.2994804382324,
-38.7673301696777,-7.60183763504028,
5.92791128158569,40.7854194641113,
11.6127243041992,54.4917259216309,
-41.2057991027832,28.3661594390869,
-79.2364883422852,-6.55292844772339,
-42.3042449951172,-26.3253860473633,
34.7275886535645,-37.9100341796875,
72.4395370483398,-48.9153633117676,
46.1534690856934,-46.1195449829102,
1.44829440116882,-19.6289024353027,
-19.8424453735352,12.9675855636597,
-14.2274951934814,31.5350608825684,
1.81106925010681,30.2809028625488,
21.6462802886963,26.3052177429199,
30.7457160949707,38.7785034179688,
7.74483489990234,57.5762481689453,
-34.4692001342773,50.0794486999512,
-49.1514625549316,8.07678031921387,
-18.2870540618897,-30.4906692504883,
11.5567808151245,-24.7593345642090,
-0.572913885116577,16.2871799468994,
-35.8718490600586,40.4666442871094,
-39.5553703308106,19.1251010894775,
-5.65658712387085,-12.9411983489990,
22.5023708343506,-4.65294027328491,
20.1580543518066,37.8579559326172,
12.5607500076294,62.9608078002930,
23.4010219573975,43.2238883972168,
28.3673553466797,9.73798370361328,
1.27462029457092,4.97115468978882,
-33.4116477966309,31.0649566650391,
-33.9736289978027,51.5437240600586,
-9.79490661621094,44.2364616394043,
-8.35894012451172,15.5646047592163,
-38.9793090820313,-14.9369955062866,
-50.7204170227051,-35.2352828979492,
-8.49693107604981,-38.4000091552734,
55.3519554138184,-21.2368164062500,
75.0397872924805,8.49509906768799,
33.1233825683594,33.2366828918457,
-22.4739723205566,39.4688034057617,
-41.4353561401367,22.8994483947754,
-21.6818199157715,-3.15224647521973,
8.86205101013184,-21.4753742218018,
26.5786075592041,-20.1127891540527,
25.5250549316406,4.09590339660645,
7.78603887557983,29.6256561279297,
-16.8131828308105,31.5985031127930,
-33.5117950439453,5.73623514175415,
-35.5620346069336,-26.4332675933838,
-29.0058879852295,-42.2490806579590,
-25.7826347351074,-38.2704315185547,
-31.2063102722168,-33.9295501708984,
-37.8257942199707,-40.8501510620117,
-35.6704216003418,-46.6395874023438,
-27.7494087219238,-42.0616645812988,
-21.9435997009277,-33.3822631835938,
-16.2872238159180,-35.5018463134766,
-6.99020862579346,-44.7263221740723,
8.62594795227051,-31.7887382507324,
26.4925727844238,12.5500240325928,
30.1500110626221,57.4982910156250,
10.3470439910889,55.7440452575684,
-17.9278450012207,8.13566875457764,
-24.2376003265381,-33.9475479125977,
4.29778051376343,-26.0867214202881,
42.0243835449219,13.8278617858887,
52.0199050903320,27.9952259063721,
25.7731933593750,-8.33427524566650,
-2.00026774406433,-56.2910728454590,
-2.97169589996338,-66.6275558471680,
8.16428661346436,-38.1766128540039,
-1.14869832992554,-13.1199064254761,
-21.1589603424072,-17.1245098114014,
-14.6063480377197,-37.9832992553711,
26.9655284881592,-44.7508354187012,
55.2488784790039,-34.1002540588379,
29.2002391815186,-24.8257560729980,
-25.9243640899658,-28.7930068969727,
-46.9239234924316,-38.6134567260742,
-21.1153697967529,-39.7659568786621,
3.87861323356628,-29.9357852935791,
-9.46132087707520,-15.9735574722290,
-33.0363807678223,-4.90171527862549,
-22.4571685791016,9.59002971649170,
12.1702690124512,29.7594261169434,
20.0515804290772,37.8488616943359,
-12.8499774932861,17.4833602905273,
-44.4482192993164,-19.0582160949707,
-37.0927963256836,-39.2615966796875,
-4.67558002471924,-16.3028030395508,
14.1368570327759,27.1618270874023,
8.34549999237061,38.3691482543945,
1.58471333980560,-2.99985384941101,
11.8961105346680,-52.8034248352051,
36.0637016296387,-60.0310707092285,
57.2734985351563,-33.0968208312988,
65.4279251098633,-21.5623073577881,
53.7322959899902,-42.3238372802734,
21.1011810302734,-50.1629066467285,
-14.2601623535156,-8.08897304534912,
-31.2528266906738,43.8577957153320,
-27.2088928222656,38.1779632568359,
-18.5554027557373,-21.5945816040039,
-15.0166568756104,-57.2401847839356,
-14.5392894744873,-25.1555404663086,
-10.2419185638428,27.1133213043213,
-7.19983148574829,34.8723144531250,
-16.6654624938965,5.18535614013672,
-34.2330360412598,-8.99365520477295,
-45.7070350646973,2.29708480834961,
-42.5487060546875,-5.74567461013794,
-24.9800987243652,-44.3982696533203,
7.51197052001953,-63.7465820312500,
44.7264289855957,-28.4234275817871,
62.9254989624023,30.3216342926025,
49.0578041076660,52.3892288208008,
21.9076404571533,32.4675865173340,
19.5700988769531,11.0231151580811,
47.2637252807617,6.51252794265747,
67.6799163818359,-3.28928494453430,
48.5320281982422,-20.7269420623779,
10.5320997238159,-20.1663150787354,
-0.962005496025085,5.12884521484375,
28.1264495849609,26.6480140686035,
57.8330345153809,13.0454607009888,
54.5098762512207,-24.9280300140381,
33.6981391906738,-44.1490516662598,
27.9509582519531,-27.7767333984375,
38.8448143005371,4.39949131011963,
42.0209770202637,30.1421127319336,
18.3989048004150,39.2549591064453,
-20.6073303222656,33.5339012145996,
-45.7893524169922,20.2601127624512,
-38.0805435180664,23.3377361297607,
-5.84689140319824,47.6039161682129,
22.7866973876953,64.1269989013672,
12.4967966079712,37.4854011535645,
-40.7480773925781,-18.6874122619629,
-87.0986633300781,-49.3822860717773,
-68.9764175415039,-27.9665107727051,
-3.02217674255371,6.26861143112183,
32.9066390991211,1.12246584892273,
0.363946914672852,-33.8963508605957,
-42.7727127075195,-43.6387481689453,
-28.2019290924072,-6.13499069213867,
24.4433593750000,36.2528152465820,
29.4339694976807,44.7300300598145,
-29.0005226135254,27.8132934570313,
-67.7783279418945,16.8861312866211,
-24.0892601013184,18.3921756744385,
44.8423995971680,18.6042861938477,
42.7889175415039,12.4657363891602,
-27.3953437805176,11.6943302154541,
-70.4543151855469,15.3564596176147,
-37.8987503051758,14.4899301528931,
16.2465591430664,3.33988404273987,
22.3370742797852,-10.4755945205688,
-4.31753110885620,-23.8583126068115,
-13.0401773452759,-42.9295043945313,
8.31671810150147,-58.6509628295898,
20.6851177215576,-50.7259140014648,
3.29320359230042,-17.0225086212158,
-17.9025535583496,9.30587673187256,
-16.4752788543701,10.8599348068237,
-1.49956846237183,5.95315885543823,
6.32527923583984,20.2327079772949,
6.28975248336792,50.5158805847168,
1.77186274528503,64.4342575073242,
-12.1533927917480,49.3284568786621,
-30.3121509552002,28.7033329010010,
-39.8689498901367,23.9766387939453,
-41.0283164978027,25.5508365631104,
-45.9122886657715,19.0004997253418,
-61.4676742553711,7.20344066619873,
-69.5047988891602,-7.53015899658203,
-45.7033843994141,-30.5368881225586,
-2.68559217453003,-55.1875724792481,
20.0989589691162,-52.8977241516113,
11.6970624923706,-4.15938901901245,
-5.50499820709229,50.3499603271484,
-13.2997322082520,49.8137207031250,
-18.6387634277344,-5.23759078979492,
-27.3026485443115,-46.7356986999512,
-29.2066535949707,-22.3600387573242,
-19.0743331909180,28.0018577575684,
-14.5931825637817,28.0638141632080,
-29.8220863342285,-27.8253974914551,
-40.5841484069824,-63.2440681457520,
-15.4794445037842,-27.3109760284424,
34.6543693542481,39.7367897033691,
52.8635520935059,62.5475616455078,
11.5574016571045,21.1130828857422,
-52.6699256896973,-33.8160095214844,
-74.3144607543945,-45.3400268554688,
-43.8784408569336,-14.1238136291504,
0.902838349342346,18.8458690643311,
25.3351478576660,16.3512153625488,
25.7315387725830,-19.9507598876953,
19.1419067382813,-57.4262237548828,
11.8540468215942,-60.8598861694336,
3.50613498687744,-25.5604190826416,
-6.06541347503662,11.1261072158813,
-14.2266426086426,14.0622053146362,
-21.2411670684814,-7.23351764678955,
-22.8149967193604,-12.0732288360596,
-16.5316066741943,4.50147533416748,
-11.0140399932861,12.1954154968262,
-23.4617862701416,-15.1092462539673,
-54.6429252624512,-49.6355590820313,
-67.6689605712891,-44.6473922729492,
-36.5969543457031,-4.42452001571655,
13.6736955642700,26.0233230590820,
36.8342666625977,24.6359920501709,
11.6039247512817,18.7519359588623,
-29.3588256835938,31.8770332336426,
-49.0039482116699,43.8194961547852,
-45.5780563354492,23.0818214416504,
-42.6486854553223,-19.7678127288818,
-47.6509323120117,-46.6049270629883,
-49.3408050537109,-46.0510940551758,
-41.0910873413086,-43.6747016906738,
-24.1183738708496,-57.4283103942871,
5.89647006988525,-73.1932601928711,
43.8816108703613,-66.0455245971680,
63.9476776123047,-34.8382339477539,
39.9208679199219,5.13951683044434,
-15.3673620223999,44.2780342102051,
-52.6814956665039,68.3064422607422,
-50.6207542419434,59.7563133239746,
-37.1862983703613,26.8942928314209,
-46.2335472106934,6.34816312789917,
-61.9063491821289,21.0129051208496,
-40.8570938110352,42.8082389831543,
10.4038887023926,22.6888465881348,
37.6865234375000,-31.5522384643555,
17.0858535766602,-65.0957260131836,
-8.11759662628174,-45.5743980407715,
7.89536762237549,-9.30220031738281,
46.4033813476563,-8.76181411743164,
58.2728271484375,-30.6567287445068,
29.7201271057129,-20.1979045867920,
-0.392773270606995,34.0537872314453,
-5.39069938659668,78.5051498413086,
1.30146765708923,59.0938072204590,
-3.54105210304260,-6.62902975082398,
-8.32221126556397,-50.5870742797852,
8.62258148193359,-35.4725837707520,
36.3908424377441,15.9518766403198,
51.4152526855469,45.9379615783691,
40.5157241821289,27.9912509918213,
11.2453632354736,-15.1175384521484,
-28.1836662292480,-40.1426086425781,
-60.7973442077637,-29.4611434936523,
-59.6526756286621,0.673692643642426,
-16.3053493499756,22.0000762939453,
33.9082183837891,20.8248882293701,
40.8379440307617,10.2478275299072,
6.21469497680664,3.77628040313721,
-12.8522272109985,-5.70951366424561,
14.4085140228271,-20.5076942443848,
49.8789482116699,-24.3313121795654,
37.0371475219727,-4.99300861358643,
-15.7888154983521,27.4609966278076,
-51.0317993164063,41.4295158386231,
-42.6439933776856,18.1742687225342,
-25.9814262390137,-20.3396434783936,
-33.6912307739258,-42.4358406066895,
-50.4514732360840,-42.6258926391602,
-36.7416915893555,-31.6285762786865,
3.70932435989380,-15.5305500030518,
27.6390018463135,5.76869201660156,
11.4777536392212,20.0063457489014,
-21.0627079010010,4.80356693267822,
-25.3200130462647,-36.4862098693848,
4.54431390762329,-62.5805015563965,
39.1659584045410,-41.4224472045898,
52.6880378723145,6.40193653106689,
39.9311485290527,26.4294853210449,
19.9611186981201,1.01953744888306,
15.6120500564575,-32.8785095214844,
25.4841403961182,-30.8466415405273,
34.4161872863770,3.28969812393188,
29.9185733795166,26.5306682586670,
9.82636070251465,19.8090400695801,
-13.6196260452271,1.94692933559418,
-31.4947471618652,-6.71548175811768,
-37.3404426574707,-5.48596906661987,
-26.2374763488770,-9.13863277435303,
6.86140823364258,-16.8194236755371,
46.7035865783691,-16.5593185424805,
55.4995574951172,-6.32371950149536,
14.7966432571411,2.15062165260315,
-41.3824882507324,-3.43871498107910,
-55.9560737609863,-21.3030834197998,
-10.1938610076904,-36.0744705200195,
48.2509880065918,-31.9061927795410,
60.4246482849121,-1.93359375000000,
23.3398704528809,32.6668739318848,
-17.8157463073730,37.4205017089844,
-27.4687767028809,6.11544084548950,
-14.0471305847168,-30.3738632202148,
-3.38877820968628,-31.6202449798584,
-0.0761609971523285,2.00452709197998,
3.97759866714478,28.1621589660645,
6.32585716247559,19.2136249542236,
-1.20809864997864,-6.93596076965332,
-12.9836568832397,-15.9877262115479,
-12.7416210174561,-6.24018192291260,
2.18953990936279,-2.12934374809265,
10.8721284866333,-7.74142408370972,
-1.01246643066406,-1.10572040081024,
-24.8552265167236,27.6927394866943,
-42.4293212890625,50.0964851379395,
-45.6057968139648,31.1724319458008,
-41.7051239013672,-19.8410758972168,
-32.9553375244141,-59.1709060668945,
-18.7150268554688,-57.0428276062012,
-0.224198579788208,-21.9559745788574,
15.4181585311890,17.2735176086426,
23.2934741973877,41.1521530151367,
24.4312648773193,50.4965209960938,
15.9277057647705,45.1524085998535,
-2.10535120964050,24.4626903533936,
-22.6803131103516,0.0281802415847778,
-31.5449981689453,-10.3563642501831,
-18.4126663208008,0.702982485294342,
6.55020236968994,20.9422950744629,
22.0335903167725,24.7034893035889,
18.1655788421631,5.37113094329834,
3.59927654266357,-18.8472900390625,
-7.46162700653076,-21.3695640563965,
2.19535017013550,-5.01259517669678,
27.3761787414551,6.68577003479004,
43.8912811279297,-6.10889244079590,
25.6137390136719,-34.5319366455078,
-24.0337524414063,-47.5010795593262,
-64.9627532958984,-34.4589843750000,
-56.0787849426270,-15.0916223526001,
-6.88846063613892,-14.4117612838745,
24.1314353942871,-29.2108879089355,
2.60375499725342,-29.5941276550293,
-41.2138023376465,-1.70377683639526,
-46.5857276916504,34.1944427490234,
-2.96191525459290,48.4166526794434,
29.5561752319336,34.8930244445801,
0.725875854492188,21.4460906982422,
-60.7967376708984,28.0379791259766,
-81.2503738403320,44.3963508605957,
-32.7230606079102,47.4959869384766,
32.4190063476563,29.0565109252930,
43.2732200622559,2.92527222633362,
-1.78954458236694,-18.1027297973633,
-41.3176765441895,-32.0534210205078,
-24.0075778961182,-40.6911544799805,
32.3271484375000,-34.3757591247559,
68.0995788574219,-12.4104766845703,
54.2845001220703,11.3361740112305,
13.5821075439453,23.3832054138184,
-6.56791353225708,25.8492717742920,
7.43040180206299,35.1118469238281,
24.2132148742676,55.5799179077148,
10.5526514053345,69.3247070312500,
-16.5051536560059,54.7459907531738,
-17.1582298278809,19.3459873199463,
17.3924598693848,-12.7629747390747,
49.1420898437500,-22.0699176788330,
38.0170440673828,-13.5909061431885,
3.32132244110107,-11.5676012039185,
-0.246729254722595,-26.9293689727783,
28.0323829650879,-39.2961692810059,
35.1268539428711,-22.2452430725098,
-7.14396047592163,26.3482379913330,
-54.9303817749023,69.0956954956055,
-51.5483474731445,68.5570831298828,
-6.26976108551025,28.8228607177734,
18.3534297943115,-10.0559072494507,
8.40960502624512,-17.3317222595215,
7.87463712692261,-10.4563159942627,
40.6396980285645,-20.7584934234619,
61.0896987915039,-43.0177650451660,
24.7595329284668,-42.2642364501953,
-32.4728736877441,-11.0575084686279,
-35.5739784240723,16.7730484008789,
21.9793319702148,5.29483127593994,
70.6102828979492,-30.8149719238281,
62.9381103515625,-52.5420989990234,
22.2740058898926,-40.2352867126465,
-0.574677348136902,-12.1544065475464,
4.51879692077637,14.9483718872070,
19.4283523559570,42.9767303466797,
35.3366546630859,65.9173431396484,
46.3639030456543,65.6913986206055,
38.8517112731934,40.5615005493164,
7.39189338684082,23.5403556823730,
-20.4028110504150,34.8474617004395,
-7.55356597900391,53.0393524169922,
24.5721530914307,44.2139511108398,
19.2808322906494,14.2090015411377,
-31.5465965270996,-4.92030334472656,
-66.9968109130859,-11.6034679412842,
-36.4130516052246,-32.0590972900391,
32.6494865417481,-66.1966018676758,
72.7921371459961,-65.5034255981445,
50.8195991516113,-5.67634820938110,
-1.31062674522400,53.6644363403320,
-38.8093376159668,45.9352340698242,
-39.8274078369141,-13.0026397705078,
-6.08988571166992,-43.2715911865234,
39.8292999267578,-8.85675525665283,
57.4721031188965,38.3358726501465,
19.4869441986084,41.9651451110840,
-46.1593284606934,6.84222221374512,
-68.5562057495117,-22.1519832611084,
-21.6252975463867,-27.1820507049561,
43.1672935485840,-20.7580928802490,
62.8041877746582,-7.16469383239746,
34.1334953308106,18.8205966949463,
2.34752130508423,36.7996025085449,
-2.67350006103516,18.4420375823975,
5.55244922637939,-24.8584537506104,
8.63279151916504,-46.5785064697266,
8.34243774414063,-30.8270587921143,
1.32518231868744,-8.75672054290772,
-24.6745109558105,-5.59415531158447,
-51.4352035522461,-9.93509769439697,
-41.9839591979981,-2.94764709472656,
8.57054328918457,4.78890180587769,
45.6356582641602,-11.6030063629150,
19.2074146270752,-36.9928550720215,
-35.9583091735840,-32.2693786621094,
-42.8055801391602,1.82427430152893,
6.77092885971069,22.5125408172607,
44.1643638610840,11.7447080612183,
14.2559852600098,-4.07532501220703,
-48.9907188415527,2.04799532890320,
-66.9786987304688,15.7561674118042,
-31.6588973999023,11.4278383255005,
-3.88271951675415,1.03696155548096,
-22.8473186492920,3.60679841041565,
-59.9900817871094,10.4098844528198,
-64.6709213256836,-6.03290557861328,
-29.2124252319336,-41.8699798583984,
8.18829154968262,-57.1600875854492,
16.8510189056397,-36.2969093322754,
0.499042391777039,-18.0119495391846,
-11.5958585739136,-34.4725112915039,
4.03684806823731,-59.5682868957520,
35.8182868957520,-47.9199409484863,
51.3386383056641,-0.0425820350646973,
25.3977737426758,38.3386077880859,
-29.9018611907959,33.1563873291016,
-64.8862838745117,-4.41981315612793,
-44.4431304931641,-41.1465873718262,
3.66777276992798,-54.5108108520508,
27.5098037719727,-36.3580932617188,
12.9625902175903,7.20285081863403,
-10.9808616638184,45.6741180419922,
-16.6842670440674,39.5043525695801,
-7.80739212036133,-8.23665142059326,
2.07875061035156,-43.5971565246582,
16.0083160400391,-21.9469890594482,
34.5356903076172,30.7934265136719,
35.3172836303711,51.6141433715820,
0.283967375755310,20.9819297790527,
-39.9062690734863,-13.9932346343994,
-36.2393836975098,-14.7116174697876,
4.53773736953735,8.82788085937500,
23.0490036010742,14.7837314605713,
-11.9797182083130,-1.74123334884644,
-55.1602249145508,-11.1111993789673,
-48.9330329895020,-0.448510706424713,
-2.63466882705688,9.23018360137940,
32.4224090576172,-4.19141006469727,
36.0791816711426,-30.3988380432129,
35.2399368286133,-34.6037216186523,
38.6455001831055,-7.02141952514648,
19.1454963684082,31.1997165679932,
-29.0594520568848,41.1765670776367,
-56.1897010803223,7.37390804290772,
-25.0722503662109,-48.0947036743164,
28.9545860290527,-82.0161972045898,
46.5559806823731,-71.3093566894531,
26.9828987121582,-25.9230041503906,
16.7572021484375,23.7044181823730,
28.8770523071289,47.6706123352051,
28.4718589782715,39.2774543762207,
-2.86753320693970,9.34770011901856,
-28.7071933746338,-20.4528160095215,
-13.5914592742920,-29.6118450164795,
23.8953189849854,-5.96666336059570,
39.1196899414063,33.8603591918945,
32.8218574523926,60.0124130249023,
33.6357307434082,58.6612243652344,
38.0352554321289,46.8727607727051,
16.9600753784180,44.4954414367676,
-25.9524593353272,45.2935714721680,
-47.2274475097656,22.6667480468750,
-23.8904113769531,-27.4082508087158,
14.4598913192749,-67.7225189208984,
28.7762222290039,-64.7993774414063,
18.0263862609863,-25.4008522033691,
10.2945709228516,9.31560897827148,
13.2015686035156,20.8834533691406,
13.5894298553467,28.2063598632813,
11.8911285400391,47.8221626281738,
18.5472850799561,64.6318206787109,
21.0120811462402,59.6260337829590,
-2.71055746078491,39.8521003723145,
-44.5917434692383,32.2823410034180,
-61.0521163940430,38.8633613586426,
-31.1574020385742,30.8523941040039,
12.6705379486084,-3.90773773193359,
32.8677368164063,-34.3064270019531,
27.3248291015625,-29.5009956359863,
20.3812732696533,0.0962589308619499,
19.8043251037598,14.9837217330933,
8.90530776977539,-0.605577230453491,
-12.7447566986084,-24.1045036315918,
-15.6717586517334,-33.6991004943848,
10.2860984802246,-22.2202529907227,
35.9783554077148,4.68909645080566,
26.7189292907715,43.9769706726074,
-14.1373558044434,76.4449234008789,
-54.4141311645508,66.9755935668945,
-64.8181991577148,10.1865806579590,
-40.7022171020508,-52.6055526733398,
4.06754589080811,-67.3588409423828,
41.0644874572754,-33.3614387512207,
47.8158950805664,1.21551156044006,
20.1844882965088,4.69300508499146,
-8.85331916809082,-4.75936079025269,
-0.999466896057129,-5.68347549438477,
35.8658714294434,1.33999109268188,
58.6987915039063,2.06041002273560,
44.7535552978516,3.79124283790588,
20.0848407745361,25.1131019592285,
15.5862255096436,61.3035697937012,
18.2116107940674,76.1106796264648,
1.34111142158508,48.6906127929688,
-25.8833332061768,0.0176427364349365,
-26.6509494781494,-35.1094474792481,
2.41482710838318,-36.9895782470703,
19.7781734466553,-10.8560867309570,
-7.44034242630005,16.2328910827637,
-50.6443672180176,9.04782390594482,
-58.6147918701172,-38.0879058837891,
-23.2058982849121,-85.5425567626953,
14.2948074340820,-84.2217407226563,
23.9929466247559,-36.8227691650391,
7.35105371475220,-5.24664258956909,
-18.6857128143311,-27.0076198577881,
-36.4499244689941,-57.8493957519531,
-31.3879833221436,-34.8857841491699,
-2.25441527366638,25.6266536712647,
31.5273265838623,42.2665443420410,
45.0159759521484,-6.90044784545898,
40.1180610656738,-42.0536918640137,
40.7243804931641,-2.08150529861450,
50.1788825988770,68.5030822753906,
34.2699661254883,72.5165023803711,
-19.2920265197754,1.53050041198730,
-59.4272766113281,-54.0600700378418,
-30.9884262084961,-34.1431617736816,
36.7745933532715,21.2021102905273,
61.1814613342285,44.1311073303223,
13.2103385925293,23.0287532806397,
-48.1471328735352,-2.89405369758606,
-57.9223785400391,-20.6542110443115,
-29.0505237579346,-42.1226844787598,
-17.3923015594482,-55.0074195861816,
-31.4743385314941,-27.9573001861572,
-36.1765785217285,25.3589305877686,
-18.4071159362793,47.7731857299805,
-11.6444301605225,6.36721801757813,
-32.8497619628906,-60.5065956115723,
-47.5251464843750,-85.6156387329102,
-30.9474601745605,-48.9627304077148,
-0.542348623275757,6.31067657470703,
10.8214864730835,27.9545707702637,
10.0611619949341,12.4084577560425,
19.7196083068848,-16.4358482360840,
31.7466602325439,-27.4010715484619,
22.0675277709961,-9.38227367401123,
-7.54333972930908,17.3219184875488,
-24.0580215454102,25.2667732238770,
-18.5007095336914,3.36357259750366,
-22.8627834320068,-27.1332283020020,
-44.5452651977539,-36.3558540344238,
-47.7894134521484,-19.3567199707031,
-6.92323493957520,3.53254652023315,
34.8891983032227,13.7428760528564,
23.3262329101563,11.9759359359741,
-32.7042388916016,6.70568943023682,
-65.6054611206055,-0.994703173637390,
-39.9231033325195,-20.2871093750000,
13.2290039062500,-41.5049133300781,
41.7701148986816,-47.0619087219238,
38.1785240173340,-26.2653865814209,
27.4165172576904,10.3355216979980,
20.4257717132568,38.0349006652832,
7.17447471618652,43.1942634582520,
-10.0843610763550,34.1769332885742,
-24.3319778442383,31.2794532775879,
-37.9182319641113,41.5821838378906,
-52.9190483093262,44.0283050537109,
-53.9114990234375,15.4523401260376,
-24.6141433715820,-29.3431262969971,
17.8762817382813,-48.9947929382324,
40.8888549804688,-18.8907604217529,
33.7352752685547,36.2523345947266,
22.0815048217773,62.9490585327148,
24.8454246520996,42.5305671691895,
23.7782096862793,9.60974502563477,
0.925805985927582,-0.367312818765640,
-18.1392230987549,8.32383155822754,
1.07469415664673,8.23234176635742,
41.0709495544434,-6.33795547485352,
55.1715698242188,-12.4854621887207,
33.7605705261231,2.89177989959717,
14.5089120864868,13.9816274642944,
19.5382041931152,-2.80512452125549,
23.3892726898193,-32.8756523132324,
0.468543410301209,-37.2264595031738,
-20.8786334991455,-18.0546035766602,
-3.07151579856873,-13.9200096130371,
37.3443412780762,-41.7329559326172,
45.6041641235352,-59.5979461669922,
7.02628898620606,-24.3730869293213,
-29.1419849395752,38.2602882385254,
-30.0979652404785,57.0172004699707,
-19.2751178741455,12.4374246597290,
-32.7415771484375,-39.9962654113770,
-54.6081390380859,-41.7145767211914,
-46.7265739440918,-5.78851890563965,
-11.3143224716187,18.4750633239746,
13.5498685836792,18.8285636901855,
5.45427703857422,20.6809215545654,
-12.2305889129639,32.7560348510742,
-9.61257457733154,40.0145492553711,
11.5905570983887,38.0037384033203,
27.3581829071045,44.7621498107910,
32.5485610961914,55.4558982849121,
32.9201393127441,43.7256622314453,
27.5609111785889,4.11370277404785,
11.1597204208374,-22.9208297729492,
-10.0627574920654,-7.70341777801514,
-28.6336765289307,19.8587894439697,
-37.7027816772461,10.7992925643921,
-31.2394294738770,-25.2571525573730,
-10.4590845108032,-31.8036251068115,
12.1993017196655,1.67837619781494,
12.7225313186646,24.7894401550293,
-14.1572818756104,3.61699438095093,
-32.4941596984863,-36.6679916381836,
-5.23375129699707,-51.2353782653809,
49.8381958007813,-41.4902153015137,
73.8306808471680,-36.4350280761719,
45.8889923095703,-39.9307746887207,
13.0598583221436,-31.2327556610107,
21.0861835479736,-16.0070686340332,
50.3285751342773,-18.2442855834961,
43.7423744201660,-39.5356864929199,
-3.46786355972290,-42.1761093139648,
-34.0880432128906,-12.2289419174194,
-9.67953014373779,12.5235967636108,
34.9720840454102,-2.18225193023682,
39.7820777893066,-31.4090671539307,
-0.353192329406738,-26.9180526733398,
-35.4167633056641,14.9350452423096,
-32.5256958007813,46.0663032531738,
-9.40703487396240,32.2556915283203,
1.15370297431946,-9.21376132965088,
-1.36079037189484,-30.3816623687744,
2.95109820365906,-17.5830421447754,
13.7665605545044,12.1548395156860,
17.1235294342041,36.5345611572266,
1.31732273101807,46.3203620910645,
-19.9827213287354,39.4387130737305,
-26.1287288665772,22.6478519439697,
-13.2247400283813,8.58301448822022,
0.588315606117249,2.66868448257446,
1.03727054595947,-2.10224676132202,
-12.6353225708008,-12.9634313583374,
-31.3763504028320,-24.3771781921387,
-39.1671943664551,-26.5496253967285,
-31.2749404907227,-27.9347858428955,
-20.1678848266602,-42.9912757873535,
-9.26661014556885,-67.6928482055664,
7.43584346771240,-71.6306610107422,
34.7220726013184,-37.0163078308106,
53.2033157348633,8.49615287780762,
39.2738914489746,26.4254016876221,
-0.207664489746094,11.8966293334961,
-25.8953456878662,2.09745860099793,
-9.36431884765625,25.1298599243164,
20.6593036651611,57.4024658203125,
20.6038246154785,59.0841026306152,
-3.13130187988281,19.9896354675293,
-3.43793678283691,-21.6521415710449,
33.1917839050293,-22.7718505859375,
56.6432037353516,13.7849197387695,
23.7879543304443,46.2875785827637,
-37.7331275939941,38.9448165893555,
-67.5323181152344,-0.0752789974212647,
-52.4845657348633,-36.2498245239258,
-34.1038894653320,-44.9600028991699,
-36.9117965698242,-37.5161972045898,
-29.7087478637695,-36.2264099121094,
11.3653297424316,-34.7266540527344,
57.2166023254395,-10.3040428161621,
63.3502731323242,30.2820510864258,
35.5835227966309,51.7520523071289,
13.4239091873169,32.4579010009766,
12.9104700088501,3.54474973678589,
18.4072399139404,11.1977500915527,
23.2237777709961,57.3663177490234,
32.7604141235352,84.1246795654297,
36.1721801757813,54.9067115783691,
6.71936702728272,7.06901264190674,
-46.5568084716797,1.88056063652039,
-69.5453491210938,33.8180503845215,
-31.0940189361572,43.9044227600098,
25.9152107238770,6.00862789154053,
35.2964935302734,-30.2090644836426,
-2.77432489395142,-13.7031688690186,
-26.1233367919922,35.2674598693848,
-2.98075819015503,50.9775810241699,
30.4544811248779,24.0969409942627,
33.0493011474609,6.58598804473877,
12.6548824310303,24.8666477203369,
6.86096763610840,44.0610694885254,
20.8107509613037,25.2707328796387,
22.5940303802490,-7.63178157806397,
0.512819766998291,-16.6007061004639,
-16.2410736083984,-12.7284908294678,
0.146882057189941,-29.6234741210938,
35.9678726196289,-54.0740089416504,
47.7301177978516,-42.5799980163574,
17.0496883392334,5.44295692443848,
-24.7902755737305,28.4110698699951,
-40.6458015441895,-4.24461936950684,
-20.9135837554932,-48.1390419006348,
7.02567100524902,-45.7753219604492,
14.6408243179321,-8.22376823425293,
1.00027775764465,17.1746177673340,
-18.2239227294922,23.6731777191162,
-39.2130432128906,35.3086929321289,
-57.5940284729004,45.5397720336914,
-58.6409416198731,16.9686431884766,
-25.9067344665527,-40.9914321899414,
24.8293952941895,-66.7969284057617,
52.5014686584473,-28.7695770263672,
39.0531425476074,24.3104648590088,
13.4109001159668,20.0209331512451,
16.7638015747070,-34.0787086486816,
40.9493560791016,-68.6830902099609,
38.6843872070313,-47.2310371398926,
-0.642761707305908,-8.78326320648193,
-32.8884201049805,-0.569998860359192,
-16.7121791839600,-19.9460430145264,
31.3028869628906,-35.0434913635254,
57.1693458557129,-23.8424720764160,
43.2712097167969,7.19526386260986,
21.7341957092285,33.9303779602051,
19.9412803649902,36.1846923828125,
19.4289474487305,3.99862813949585,
-10.6446475982666,-40.7579574584961,
-51.5162124633789,-55.4902000427246,
-52.6422958374023,-20.6861572265625,
-4.92651796340942,30.6359100341797,
38.9187088012695,45.6149826049805,
26.7109146118164,16.9998416900635,
-21.4395446777344,-9.28514385223389,
-40.4153404235840,-1.69686222076416,
-7.15140533447266,18.1132564544678,
32.3519630432129,15.0976572036743,
34.3831214904785,-7.69693040847778,
13.7783927917480,-9.29036521911621,
8.75435638427734,24.5518779754639,
18.7692489624023,56.7927017211914,
18.5182151794434,46.5394287109375,
12.5781650543213,1.70136404037476,
22.6000633239746,-27.5232772827148,
39.2816810607910,-10.6551494598389,
23.8036708831787,24.8172149658203,
-23.5376434326172,30.3277263641357,
-45.5845832824707,0.285285234451294,
-11.0283355712891,-33.2354125976563,
33.8910255432129,-39.2263259887695,
30.2039031982422,-22.2758865356445,
-3.58525562286377,-10.8213596343994,
-0.216372251510620,-7.95424604415894,
40.7377700805664,7.03858661651611,
48.0622863769531,34.7310600280762,
-5.11126518249512,46.0696945190430,
-54.1444931030273,18.6296958923340,
-36.8684921264648,-24.7220172882080,
16.2934265136719,-39.3643531799316,
31.3376884460449,-13.1993598937988,
0.385361194610596,7.61734485626221,
-18.9746894836426,-16.8353214263916,
2.66055321693420,-60.0699234008789,
28.1267242431641,-62.9979934692383,
21.0327167510986,-15.0509233474731,
-1.06695652008057,24.0408916473389,
-7.07957410812378,6.53209304809570,
-6.57930898666382,-38.0584907531738,
-19.8549346923828,-40.8977088928223,
-33.7676010131836,9.91748619079590,
-21.3779182434082,53.2239799499512,
9.89770603179932,42.7204666137695,
26.6636657714844,10.7642660140991,
13.6616859436035,10.1299457550049,
-13.4293098449707,33.1516876220703,
-30.4519672393799,33.4401359558106,
-38.8989868164063,4.56939697265625,
-43.1068611145020,-16.4933242797852,
-35.8425674438477,-19.1837158203125,
-17.4409008026123,-30.3004665374756,
-7.11725568771362,-58.7122116088867,
-16.6788558959961,-65.4076919555664,
-30.6922550201416,-30.4759807586670,
-28.5485343933105,1.51777625083923,
-10.2673349380493,-18.4518451690674,
9.06020832061768,-54.4312133789063,
24.3244380950928,-40.6110763549805,
37.8056488037109,14.2001514434814,
41.9952964782715,28.3499240875244,
22.0270557403564,-16.6024723052979,
-18.1731815338135,-41.6372489929199,
-48.3038330078125,1.68006134033203,
-45.4226951599121,46.8158264160156,
-22.8494262695313,14.9209403991699,
-6.24656677246094,-58.0869979858398,
-2.49618291854858,-63.9728507995606,
-1.88991367816925,11.4402132034302,
-4.33550119400024,59.1808929443359,
-5.34094810485840,7.36719608306885,
10.3939647674561,-76.7071533203125,
47.6765899658203,-82.9569854736328,
75.9940643310547,-9.45122337341309,
59.7781448364258,57.1506500244141,
3.88736009597778,65.9454879760742,
-36.0960464477539,43.7065124511719,
-26.7704524993897,28.1755695343018,
0.778298974037170,22.6482620239258,
5.75518178939819,15.8645887374878,
-4.24151802062988,14.9027605056763,
7.19965171813965,24.7554512023926,
27.4738159179688,31.4906826019287,
15.6411218643188,20.1369762420654,
-27.1930046081543,1.50248336791992,
-46.0909004211426,-1.23293304443359,
-10.7015953063965,6.20551824569702,
27.2243156433105,10.3709354400635,
6.34611606597900,15.5756502151489,
-50.3549079895020,26.1266479492188,
-65.4419326782227,26.1261444091797,
-17.9944763183594,6.47367382049561,
34.7346305847168,-19.8192462921143,
36.0049171447754,-25.6590881347656,
4.53474426269531,-0.228121042251587,
-13.5836467742920,28.5268821716309,
-15.6473226547241,39.1129341125488,
-29.1595382690430,31.9411659240723,
-49.5261077880859,13.7359027862549,
-37.3299980163574,-18.5625267028809,
15.1856164932251,-54.4885253906250,
62.2878952026367,-60.6490592956543,
57.4019241333008,-23.8509044647217,
11.9816360473633,14.5703849792480,
-17.7751102447510,5.56777858734131,
-3.25732779502869,-38.3177604675293,
25.4613761901855,-50.3450012207031,
30.0355281829834,-1.22872543334961,
15.6051769256592,58.0995483398438,
9.01795578002930,59.7855987548828,
16.9082756042480,4.53667163848877,
14.0399751663208,-41.7908134460449,
-14.7804918289185,-38.0287857055664,
-37.5635375976563,-8.32968997955322,
-16.9883518218994,8.69233417510986,
28.0052757263184,4.63347291946411,
39.4948463439941,-4.12450504302979,
0.993684053421021,-9.78534412384033,
-35.1126098632813,-17.1302452087402,
-16.1628341674805,-22.8082771301270,
37.1640052795410,-25.3193492889404,
50.7765121459961,-30.9392433166504,
3.19248723983765,-42.7675170898438,
-46.9113349914551,-46.2131538391113,
-42.3022308349609,-24.4757690429688,
-1.60806763172150,9.27936649322510,
15.6004619598389,17.1478118896484,
-10.2255411148071,-11.3236141204834,
-34.2073974609375,-34.7130317687988,
-17.8388919830322,-14.1153469085693,
20.1365356445313,36.4482803344727,
29.7875671386719,69.2492523193359,
-3.49597716331482,56.7208061218262,
-41.9484901428223,18.5287704467773,
-43.9624099731445,-6.53772211074829,
-9.16150188446045,-8.16227531433106,
26.6088180541992,1.40639078617096,
31.9471836090088,7.99119758605957,
10.3854846954346,11.3948125839233,
-9.53137779235840,14.3832015991211,
-5.66864109039307,16.8840961456299,
17.4176902770996,16.8180713653564,
37.7166328430176,12.3233900070190,
31.6886940002441,4.59854507446289,
-1.20709908008575,1.65795063972473,
-35.5496330261231,13.0814533233643,
-42.9825057983398,32.0047111511231,
-20.4623165130615,35.2629241943359,
3.31994533538818,9.12551689147949,
-1.11538386344910,-32.2988739013672,
-24.6286487579346,-59.4192504882813,
-29.9077148437500,-54.9628944396973,
-5.10243177413940,-36.0717124938965,
17.5011081695557,-20.5657691955566,
5.55099010467529,-7.12696456909180,
-32.3570175170898,15.5041389465332,
-52.5359268188477,38.6981773376465,
-34.8834266662598,46.1717262268066,
-4.03800106048584,38.0549316406250,
12.5701799392700,26.3830070495605,
11.6150894165039,18.4789257049561,
0.574141383171082,8.38662815093994,
-17.0659313201904,-5.00644731521606,
-33.3536109924316,-7.59050750732422,
-29.8268585205078,3.68455481529236,
-2.27787399291992,6.87415742874146,
18.4052505493164,-9.72451686859131,
7.50447177886963,-29.0058727264404,
-18.1066608428955,-25.9973888397217,
-14.2189512252808,-10.3606309890747,
20.3011150360107,-18.2733058929443,
39.4471206665039,-50.6136016845703,
12.8413820266724,-61.5533752441406,
-31.7038669586182,-19.3308429718018,
-44.0517692565918,38.1032142639160,
-24.5350055694580,45.7824668884277,
-8.21820259094238,-7.03581666946411,
-11.7026176452637,-58.2253608703613,
-15.0977449417114,-51.9601745605469,
-0.665355086326599,-1.79166293144226,
18.4358921051025,29.0497989654541,
23.5751743316650,9.02692699432373,
22.5017185211182,-26.6860389709473,
34.6645851135254,-33.2234878540039,
58.4189300537109,-7.45876979827881,
68.1754760742188,14.6179885864258,
47.9658317565918,11.5778026580811,
7.94393253326416,1.08868145942688,
-27.8226070404053,8.33064460754395,
-46.3762016296387,21.4910411834717,
-44.9054908752441,12.7133197784424,
-29.1907386779785,-13.4496765136719,
-10.1587619781494,-20.7418384552002,
2.72073984146118,5.02521181106567,
5.60092878341675,32.2442512512207,
3.55707716941834,18.8654479980469,
-0.795868992805481,-28.9710922241211,
-7.62607908248901,-50.8429374694824,
-20.3274745941162,-13.0454921722412,
-32.4269943237305,45.5318717956543,
-27.9883060455322,61.1438598632813,
-4.84131908416748,22.6039104461670,
22.2472858428955,-17.6097335815430,
36.0323410034180,-10.5498437881470,
30.5360355377197,28.5660457611084,
13.4135293960571,47.3966140747070,
0.184419825673103,31.2027072906494,
3.00501728057861,15.6591463088989,
17.1486759185791,24.3696804046631,
20.5788726806641,30.2073745727539,
-1.78181576728821,3.69787526130676,
-38.1060523986816,-36.4540634155273,
-56.1337585449219,-43.5058021545410,
-42.8653602600098,-14.7375364303589,
-27.1759109497070,6.01239013671875,
-42.4316024780273,-7.58398008346558,
-69.5981292724609,-24.6228637695313,
-57.4927062988281,-14.7354087829590,
1.12401986122131,4.96761369705200,
53.4272079467773,1.20347833633423,
59.2138671875000,-19.2324619293213,
42.4528083801270,-18.5788784027100,
46.6997146606445,4.64562940597534,
63.5437927246094,12.0576753616333,
49.4453468322754,-12.6297369003296,
3.23346877098084,-36.0106124877930,
-20.0144634246826,-32.4675559997559,
1.28869283199310,-23.4852809906006,
18.7234325408936,-36.5218200683594,
-9.13897418975830,-59.0362739562988,
-44.7684974670410,-57.1659660339356,
-25.0973129272461,-29.4949932098389,
39.3544921875000,-11.3465166091919,
78.3956146240234,-16.7238368988037,
58.9575462341309,-20.2052288055420,
23.8207664489746,-5.07720184326172,
14.2713775634766,8.86649894714356,
18.8042678833008,0.141331732273102,
12.8266592025757,-17.8087291717529,
8.33778190612793,-22.2569217681885,
33.6240425109863,-14.2119026184082,
64.3173599243164,-7.15719270706177,
54.8472137451172,-1.61297965049744,
10.1847457885742,10.4227085113525,
-15.2469406127930,24.7305679321289,
6.70295286178589,20.5711059570313,
41.0938987731934,1.64979338645935,
47.5133895874023,-6.46006965637207,
26.6939735412598,7.44029235839844,
2.65574145317078,18.3583354949951,
-12.4900236129761,4.22773838043213,
-24.3693275451660,-23.7685718536377,
-33.0300865173340,-39.3591651916504,
-26.9795417785645,-39.7714996337891,
-19.7727050781250,-37.4522399902344,
-28.0507717132568,-31.0049133300781,
-43.7460937500000,-10.3430337905884,
-39.5312843322754,17.6400470733643,
-12.4513120651245,23.7103309631348,
10.0196056365967,-5.98809576034546,
17.5540904998779,-42.9702453613281,
29.2287712097168,-50.2652893066406,
45.8715095520020,-22.6702804565430,
41.0084228515625,12.0782299041748,
-0.157569766044617,30.9946460723877,
-40.1215209960938,27.2104282379150,
-27.0750579833984,6.70612335205078,
28.2779312133789,-11.1244258880615,
56.1384811401367,-1.76213598251343,
19.7134552001953,36.9724006652832,
-42.9120407104492,67.4673385620117,
-71.3568496704102,51.1471405029297,
-53.9426765441895,-4.70638561248779,
-13.0001382827759,-42.6794281005859,
28.5180320739746,-27.6586456298828,
53.1153793334961,11.2251424789429,
40.6057052612305,24.7277088165283,
-6.90131139755249,10.6120891571045,
-50.3441238403320,7.53778457641602,
-47.7708816528320,21.2800960540772,
-13.7110252380371,24.6584129333496,
-2.81524515151978,2.77674937248230,
-33.6251983642578,-19.0822811126709,
-58.5359039306641,-19.1155700683594,
-42.0426521301270,-14.0032453536987,
-15.8076286315918,-28.0582313537598,
-17.6145973205566,-51.0735473632813,
-25.5756931304932,-50.7539482116699,
-4.92454338073731,-27.6044158935547,
25.7080669403076,-10.4117116928101,
20.3677253723145,-11.7922735214233,
-22.2310562133789,-12.0776176452637,
-38.4806747436523,-6.42376232147217,
-4.47683238983154,-16.1192302703857,
22.5966129302979,-41.9804916381836,
2.35876893997192,-52.9577064514160,
-25.5138854980469,-34.4144821166992,
-3.04116296768188,-16.8726615905762,
40.2260437011719,-27.5959892272949,
35.2052459716797,-42.4993934631348,
-12.6367864608765,-15.5672645568848,
-26.1357288360596,40.4750747680664,
15.1266231536865,58.7601776123047,
42.6920890808106,20.6363468170166,
5.28940534591675,-19.9555263519287,
-43.0010986328125,-14.0065240859985,
-22.5822963714600,12.2242250442505,
47.1922111511231,10.8596105575562,
72.5447387695313,-11.8923511505127,
18.9977436065674,-12.7966365814209,
-44.6620407104492,9.60948085784912,
-53.2853660583496,15.4010887145996,
-24.8043804168701,-6.83788919448853,
-10.7976970672607,-14.9698228836060,
-16.8432865142822,19.8732528686523,
-19.6531276702881,53.8646354675293,
-12.6708202362061,30.7454528808594,
-9.91144084930420,-38.0982856750488,
-13.7517929077148,-78.5366058349609,
-7.34281063079834,-50.5064315795898,
14.7336988449097,7.29073143005371,
29.2322387695313,34.0922164916992,
20.1403827667236,11.7124137878418,
0.474465608596802,-25.6734523773193,
-11.5444135665894,-35.8161239624023,
-15.8676700592041,-12.8228626251221,
-17.5950622558594,18.8384742736816,
-15.7211284637451,29.7175045013428,
-16.0421714782715,10.5685577392578,
-26.0112705230713,-24.3070316314697,
-39.5909309387207,-52.9476509094238,
-37.0864601135254,-59.5808219909668,
-12.5977325439453,-48.1773872375488,
10.2571220397949,-29.6392650604248,
3.32698583602905,-10.7022628784180,
-28.6777877807617,4.45624971389771,
-48.9001693725586,10.2221651077271,
-35.1131057739258,4.77898216247559,
-7.45074796676636,-14.4470615386963,
4.46906280517578,-38.4500122070313,
-0.232222884893417,-50.7895812988281,
-8.99589729309082,-38.6583557128906,
-11.4950113296509,-8.09834861755371,
-7.10952425003052,16.4406433105469,
0.889460623264313,11.6271638870239,
4.80709981918335,-14.7157669067383,
-5.81341791152954,-36.7226600646973,
-30.5001678466797,-39.7512893676758,
-40.5129203796387,-31.4563846588135,
-8.14430236816406,-26.1909503936768,
42.0599555969238,-21.0939483642578,
53.5576438903809,-9.32108402252197,
8.42240810394287,0.982003569602966,
-35.9814338684082,-8.20924186706543,
-17.1281986236572,-30.1906070709229,
44.4301834106445,-38.4628906250000,
76.0295028686523,-21.2197113037109,
47.1060180664063,1.62545275688171,
6.35052394866943,3.76145935058594,
3.74101567268372,-8.25278949737549,
18.7302093505859,-0.423681646585465,
-0.749269723892212,32.6433601379395,
-50.1431884765625,56.6081886291504,
-72.3290023803711,35.2189979553223,
-36.6609535217285,-17.1551361083984,
19.2135715484619,-52.1921615600586,
41.0736999511719,-41.2030830383301,
24.8466529846191,-14.8711042404175,
6.08353233337402,-18.0050392150879,
-0.806093573570252,-46.8376235961914,
-4.29939413070679,-55.2110023498535,
-15.4642267227173,-15.2623243331909,
-24.6721611022949,42.8035812377930,
-16.7679271697998,63.8389472961426,
5.19778490066528,32.1679344177246,
20.5961837768555,-8.37135696411133,
22.9180107116699,-12.6199026107788,
22.0312690734863,15.3469343185425,
26.0686893463135,40.1494255065918,
32.4652900695801,42.6288757324219,
27.9391250610352,39.9259300231934,
1.52872550487518,47.2726097106934,
-31.6693801879883,53.5529785156250,
-31.2038764953613,32.4188385009766,
14.7639646530151,-11.5521497726440,
66.9049301147461,-36.8243446350098,
74.4660644531250,-20.5639362335205,
30.8828639984131,15.2748594284058,
-6.63346576690674,27.8233261108398,
1.44484424591064,2.48111891746521,
21.8808002471924,-22.1875476837158,
-3.32466340065002,-6.92026138305664,
-60.7847366333008,31.2186164855957,
-75.5498352050781,44.8690795898438,
-17.8366489410400,13.7436666488647,
43.7311325073242,-31.3697586059570,
35.9639244079590,-48.8408164978027,
-17.7809734344482,-34.3703422546387,
-31.4147224426270,-21.5504798889160,
15.7346544265747,-19.8539867401123,
48.5241889953613,-3.21283698081970,
5.37099266052246,39.9375762939453,
-72.7072067260742,67.1507644653320,
-102.519279479980,36.1003456115723,
-61.9150009155273,-31.7559452056885,
-9.80652999877930,-60.4389228820801,
6.17068719863892,-19.1806049346924,
-5.20919036865234,34.2807655334473,
-21.7227497100830,31.2676963806152,
-37.8651657104492,-12.2918357849121,
-48.1096115112305,-27.3211193084717,
-37.5772895812988,3.57748150825501,
-4.64929914474487,25.2637176513672,
33.6156387329102,-3.21606683731079,
53.5904312133789,-40.9650154113770,
49.5017776489258,-29.0168037414551,
33.6884040832520,18.5657634735107,
11.9780645370483,38.6639671325684,
-8.00456905364990,9.43517112731934,
-2.28773212432861,-27.5198917388916,
27.8298454284668,-34.8232536315918,
35.2182083129883,-23.6039676666260,
-9.91080474853516,-21.1948127746582,
-58.7135772705078,-26.9727878570557,
-41.6973991394043,-22.5689144134522,
27.4504451751709,-10.8622751235962,
55.9571762084961,-4.12931299209595,
3.80351781845093,4.57583141326904,
-52.9024543762207,18.4268741607666,
-31.6686096191406,21.0300102233887,
38.0453605651856,-3.92802071571350,
56.8282012939453,-37.6896171569824,
11.3860883712769,-48.4184989929199,
-12.1281747817993,-34.6836090087891,
27.3893127441406,-21.8019351959229,
66.5347290039063,-19.0129299163818,
42.9487838745117,-1.93532657623291,
-7.74932765960693,38.0966186523438,
-16.5063533782959,64.0520248413086,
14.9352121353149,39.9423675537109,
32.0324058532715,-6.61264419555664,
21.7031803131104,-17.6411628723145,
18.6532878875732,20.4134578704834,
31.2842121124268,62.5249099731445,
17.6548385620117,65.5738296508789,
-32.3630065917969,39.7742042541504,
-58.2763633728027,22.4435367584229,
-22.7455921173096,23.8303833007813,
25.1042633056641,27.3257637023926,
31.3276443481445,21.2830924987793,
15.3112325668335,12.8915548324585,
20.0556812286377,16.1940116882324,
34.3643035888672,23.6601448059082,
14.1455459594727,26.0250988006592,
-29.2092304229736,25.4898395538330,
-36.2146072387695,30.6855068206787,
1.31291675567627,38.6777610778809,
19.3824424743652,36.5404624938965,
-17.9826297760010,17.1524124145508,
-48.3456802368164,-9.75354290008545,
-14.5217800140381,-16.7183380126953,
41.1838989257813,6.52309417724609,
35.0868568420410,32.9986572265625,
-25.1558284759522,26.9888820648193,
-58.9296264648438,-18.8872699737549,
-35.7168426513672,-62.8071708679199,
-9.85489463806152,-58.4767684936523,
-26.7133274078369,-8.71475791931152,
-53.5102005004883,31.1836795806885,
-35.2105178833008,22.4976272583008,
14.9022016525269,-12.7390699386597,
44.5882720947266,-19.5070438385010,
41.9635848999023,13.3058729171753,
42.1316528320313,40.7600860595703,
54.9307518005371,23.9082088470459,
52.6937713623047,-20.2353000640869,
28.8395271301270,-41.6962318420410,
16.7934951782227,-22.6226329803467,
33.8732185363770,6.30901861190796,
51.9814300537109,11.7915372848511,
40.4330749511719,1.19766640663147,
11.9065504074097,-0.861852109432221,
4.71619749069214,16.3546199798584,
25.9253978729248,37.7118415832520,
39.2111396789551,42.0242958068848,
23.8477134704590,24.6573009490967,
-3.37515211105347,-5.68879604339600,
-14.7341756820679,-28.5413169860840,
-13.0399322509766,-22.2022895812988,
-17.4371471405029,11.7793560028076,
-30.3074188232422,41.7731208801270,
-36.8327827453613,37.5214691162109,
-25.9701213836670,5.70434427261353,
-6.66105365753174,-10.6769733428955,
4.33973789215088,13.9335203170776,
2.91982507705688,52.9237060546875,
1.25499975681305,61.0502586364746,
5.62814235687256,30.9778804779053,
2.77219176292419,0.346735954284668,
-17.1560516357422,-1.71208477020264,
-40.7569046020508,14.8239154815674,
-42.3028335571289,18.6561012268066,
-17.1247444152832,-0.203350663185120,
8.91099262237549,-20.3926410675049,
5.50863552093506,-22.1816635131836,
-17.6716632843018,-7.47312116622925,
-26.8940181732178,10.8118495941162,
-10.8817758560181,21.6474761962891,
3.96493816375732,26.7049236297607,
-9.50058078765869,28.4872074127197,
-39.2563247680664,27.3181438446045,
-49.4565582275391,22.8450870513916,
-28.9354171752930,5.51096248626709,
-4.73639488220215,-24.2771816253662,
-5.74209070205689,-47.8208770751953,
-24.9404773712158,-49.8082733154297,
-29.4097080230713,-31.1276779174805,
-4.61481332778931,-11.4511241912842,
25.6959800720215,-7.62132215499878,
31.6837692260742,-10.4763059616089,
9.75309085845947,-3.42939901351929,
-14.1303548812866,11.2173070907593,
-18.2539215087891,21.5544414520264,
-7.36597537994385,29.6686801910400,
0.846608877182007,42.1160545349121,
-3.23057389259338,42.9300384521484,
-15.7282686233521,9.69571304321289,
-26.9317111968994,-45.4721069335938,
-27.8373146057129,-67.6324691772461,
-15.5656719207764,-26.6480941772461,
3.12406492233276,32.1338996887207,
8.53290653228760,37.7689933776856,
-3.80157470703125,-13.8593502044678,
-15.6827917098999,-59.0123481750488,
-10.3482856750488,-48.4269905090332,
0.648303210735321,-13.6978559494019,
-9.60282707214356,-7.28074550628662,
-39.7055282592773,-28.3270988464355,
-55.7176055908203,-36.5704536437988,
-35.3943862915039,-20.6776027679443,
-6.75970268249512,-10.5026569366455,
-6.68387794494629,-24.8940181732178,
-23.1438350677490,-42.5641250610352,
-16.8950405120850,-36.2486038208008,
12.6986227035522,-13.4065246582031,
18.7678623199463,3.53399848937988,
-18.1941490173340,5.55360412597656,
-51.9882431030273,1.83027112483978,
-31.7890205383301,-8.22370243072510,
22.6931438446045,-29.1711883544922,
48.4805984497070,-40.7377433776856,
27.4533920288086,-22.2695426940918,
3.60509634017944,9.65112495422363,
11.4380779266357,20.6003284454346,
26.1656894683838,-2.89438295364380,
7.31867074966431,-37.6030540466309,
-33.5315132141113,-54.9429130554199,
-47.9984588623047,-44.7862663269043,
-20.1546802520752,-18.7928180694580,
17.2929286956787,11.0242309570313,
29.1209049224854,23.9084014892578,
15.4626255035400,-3.46123695373535,
-0.285625457763672,-56.9885520935059,
-1.70739567279816,-73.1010589599609,
4.91227245330811,-22.1770992279053,
4.12923288345337,42.0482215881348,
-5.52849960327148,44.8138008117676,
-15.4086608886719,-7.11313438415527,
-10.2283391952515,-34.4893302917481,
18.4111194610596,-4.48134708404541,
45.6375083923340,25.4026489257813,
40.7792549133301,0.570818662643433,
0.715303897857666,-39.7143058776856,
-40.8303871154785,-24.3476676940918,
-54.5403900146484,30.3478755950928,
-45.2662277221680,38.3262939453125,
-33.6461486816406,-17.2496528625488,
-23.4667339324951,-55.2236022949219,
-1.63820397853851,-13.6727371215820,
25.5874500274658,56.2309799194336,
26.4514980316162,65.4720153808594,
-8.54080677032471,15.0249862670898,
-43.4970626831055,-20.8109035491943,
-31.2869262695313,-6.73601341247559,
23.8160476684570,15.9383287429810,
68.2642211914063,4.34456825256348,
64.7970046997070,-22.2640438079834,
30.3839149475098,-19.9941577911377,
6.30658435821533,6.09814405441284,
6.13466072082520,16.1672325134277,
9.90682888031006,-1.52807092666626,
-4.31046915054321,-20.6801128387451,
-27.4358177185059,-19.1995334625244,
-35.3344345092773,-5.63275432586670,
-19.9772090911865,4.41698455810547,
2.49476289749146,1.24379801750183,
5.27962875366211,-12.8960094451904,
-16.1598873138428,-30.7586631774902,
-38.9736862182617,-46.2594299316406,
-36.5294609069824,-54.1940383911133,
-3.54137825965881,-48.7039031982422,
30.4582633972168,-37.0633964538574,
30.5804767608643,-27.2311458587647,
-2.28041338920593,-17.7639579772949,
-30.8726978302002,-7.79243230819702,
-18.0695056915283,4.53690481185913,
30.1319599151611,21.9137744903564,
65.9191207885742,41.8701477050781,
47.7083702087402,48.6836357116699,
-9.09412860870361,26.5945835113525,
-47.1045455932617,-14.5951786041260,
-29.1109199523926,-42.9018478393555,
16.3805236816406,-33.2275886535645,
28.4161682128906,-4.05120992660523,
-6.68053865432739,6.35298490524292,
-39.0345573425293,-14.1569032669067,
-19.8835601806641,-33.3263549804688,
31.2217960357666,-18.0744342803955,
47.9143257141113,25.0490226745605,
3.94440126419067,54.2430648803711,
-53.0556106567383,47.7660255432129,
-63.1013374328613,23.6866397857666,
-23.6342449188232,8.86727428436279,
21.5114154815674,5.31806993484497,
39.0499420166016,-3.47272706031799,
37.8740043640137,-25.1560287475586,
42.0533866882324,-39.9057731628418,
48.0852050781250,-27.9030094146729,
45.6930847167969,7.99507427215576,
35.8700218200684,41.9031982421875,
28.4872303009033,49.5646095275879,
24.1487789154053,31.9463500976563,
9.63884353637695,9.80842018127441,
-18.1855964660645,4.35553121566773,
-43.9401321411133,16.2960243225098,
-46.1424522399902,27.6534519195557,
-29.2093467712402,19.0978126525879,
-13.7868041992188,2.32084417343140,
-14.8925590515137,-0.368579089641571,
-25.1570301055908,20.5596733093262,
-16.2179622650147,39.0959701538086,
18.7511425018311,29.1108303070068,
55.3790473937988,-1.87201249599457,
60.5218467712402,-16.0447521209717,
23.3127155303955,7.35461282730103,
-27.0572204589844,42.5499496459961,
-49.3956451416016,50.6101074218750,
-26.8625259399414,20.5423851013184,
16.7115840911865,-14.8246164321899,
46.7188568115234,-18.0865859985352,
50.0964202880859,8.52678108215332,
39.6193466186523,36.5122108459473,
32.1625747680664,46.6998443603516,
23.9242534637451,43.4797019958496,
-1.92846608161926,41.8645095825195,
-38.0975074768066,42.5505790710449,
-54.7320060729981,36.3282775878906,
-33.1146697998047,25.2206153869629,
5.10203027725220,20.0532932281494,
16.5555953979492,13.2676048278809,
-8.26626205444336,-11.5593328475952,
-33.9819221496582,-47.0429306030273,
-21.8817653656006,-58.7899017333984,
16.8958950042725,-29.9038467407227,
42.3837623596191,8.03056049346924,
43.2882499694824,10.3447446823120,
42.9211769104004,-13.1887664794922,
52.5056877136231,-11.9548931121826,
45.7779083251953,26.7881031036377,
3.97613096237183,52.8872337341309,
-43.4463119506836,25.7520656585693,
-52.0418968200684,-22.0006103515625,
-13.9931182861328,-26.1267127990723,
29.8810291290283,12.1556873321533,
43.9220199584961,31.4142074584961,
32.3492012023926,3.76398515701294,
14.5650806427002,-29.6120586395264,
-3.18992543220520,-20.0295867919922,
-15.8935852050781,15.2539043426514,
-12.4328880310059,28.0259571075439,
1.05361139774323,9.99255943298340,
-0.917717814445496,-3.80781984329224,
-20.9764080047607,6.91590404510498,
-20.5388736724854,21.8371582031250,
19.5603218078613,16.2089633941650,
58.4839859008789,0.559278666973114,
37.6556243896484,-9.14733791351318,
-25.1929893493652,-15.4275169372559,
-47.8536911010742,-25.6434898376465,
6.82542610168457,-29.7998580932617,
67.5742797851563,-16.2309265136719,
56.9511146545410,10.2926979064941,
-4.61949110031128,30.2532711029053,
-33.1500205993652,35.0689392089844,
-1.94215893745422,34.8802909851074,
34.9047698974609,39.5533447265625,
29.1792392730713,42.3772392272949,
-4.71354103088379,36.2006072998047,
-29.7356605529785,19.3830947875977,
-39.5048065185547,-7.89070367813110,
-45.2367477416992,-43.3592987060547,
-35.7236785888672,-71.2996215820313,
-2.52876853942871,-68.8777465820313,
26.7582817077637,-30.6580505371094,
15.6771373748779,15.3381347656250,
-28.1021556854248,31.1029453277588,
-55.1799278259277,10.4668645858765,
-46.3578567504883,-17.2628402709961,
-39.1508026123047,-22.2553710937500,
-50.1243171691895,-6.31324386596680,
-52.1927909851074,0.0545630753040314,
-17.1235275268555,-18.3124961853027,
29.9705123901367,-42.4867477416992,
33.5521469116211,-45.1926155090332,
-11.8727664947510,-29.3828372955322,
-44.5378646850586,-21.8692512512207,
-19.9996299743652,-38.4437522888184,
34.7836265563965,-53.3191795349121,
58.9864997863770,-35.2306594848633,
29.3176689147949,4.65558958053589,
-17.8209304809570,24.2543277740479,
-33.9211730957031,-0.608369827270508,
-7.48651361465454,-35.8285293579102,
38.5419502258301,-33.2327194213867,
70.3060989379883,5.74748420715332,
64.8355255126953,36.6642150878906,
26.9367179870605,22.8919601440430,
-15.9539422988892,-17.5472850799561,
-34.4434204101563,-41.0506973266602,
-12.0598907470703,-25.5270061492920,
30.9562644958496,7.89172315597534,
51.8337364196777,29.8766651153564,
29.4542751312256,27.2469177246094,
-17.5916366577148,15.2061996459961,
-52.7102165222168,13.1429080963135,
-55.2232704162598,26.2073707580566,
-42.0837326049805,36.6086311340332,
-43.3401565551758,26.6730155944824,
-50.2096328735352,-6.63999986648560,
-32.1546630859375,-41.8574066162109,
17.9577789306641,-54.1235809326172,
61.2445030212402,-40.6614990234375,
50.1992721557617,-24.4909744262695,
-10.8297176361084,-21.5750293731689,
-56.0889434814453,-32.3319816589356,
-38.9908638000488,-45.3379402160645,
15.9008541107178,-47.3802337646484,
40.5412521362305,-35.7684440612793,
5.91931343078613,-15.3347549438477,
-38.1355056762695,2.54854536056519,
-30.0457763671875,-0.367597162723541,
28.6280460357666,-23.8872966766357,
73.3797302246094,-47.0806427001953,
56.3311767578125,-46.2569427490234,
2.39247608184814,-25.1399574279785,
-27.9594631195068,-3.98819518089294,
-12.5895576477051,6.90130853652954,
10.9881200790405,20.8031711578369,
2.33184719085693,43.5445938110352,
-34.5545463562012,51.7027702331543,
-57.4823837280273,22.9044551849365,
-36.5142707824707,-23.3797264099121,
13.2323036193848,-37.9356155395508,
51.5726890563965,-1.89998292922974,
48.7646942138672,46.9616928100586,
14.9505949020386,61.0274276733398,
-8.59724330902100,35.6569061279297,
1.86225640773773,9.59572505950928,
27.5276069641113,6.32217884063721,
31.8313903808594,7.53412628173828,
2.60814380645752,-9.42602825164795,
-31.1495265960693,-31.2399787902832,
-35.7600402832031,-30.6175270080566,
-18.1114234924316,-4.80896282196045,
-7.49930810928345,11.4588479995728,
-4.37043094635010,-7.95814418792725,
9.05684757232666,-39.6933937072754,
30.7633800506592,-40.0670967102051,
33.3128662109375,-0.623198032379150,
10.8036489486694,38.5837211608887,
-5.93050003051758,35.4656639099121,
8.86746215820313,-2.72638893127441,
30.9526157379150,-28.8992080688477,
18.8658943176270,-11.3976640701294,
-20.8176422119141,20.6943035125732,
-41.5805740356445,20.1555480957031,
-29.3854370117188,-12.0416908264160,
-21.4802227020264,-25.0817623138428,
-37.6262855529785,11.3154830932617,
-44.2241058349609,58.4457359313965,
-8.34071063995361,56.9764671325684,
38.2407035827637,0.110062599182129,
45.9707946777344,-43.0819396972656,
19.1112270355225,-21.9569396972656,
5.48964500427246,30.4365520477295,
18.6559696197510,52.4050407409668,
13.6574859619141,40.8782997131348,
-32.9657707214356,35.1317672729492,
-71.7580108642578,42.4218788146973,
-51.1763076782227,24.9996032714844,
3.45241546630859,-21.9855499267578,
18.5212821960449,-47.5036659240723,
-23.1724681854248,-19.8094139099121,
-65.9851989746094,10.6224222183228,
-60.7970809936523,-14.6364860534668,
-15.6908969879150,-61.2730102539063,
28.8567008972168,-46.9241714477539,
51.9041900634766,28.0553436279297,
47.5656509399414,70.5205612182617,
15.8827695846558,30.2088718414307,
-29.7638931274414,-24.2320995330811,
-54.9627342224121,-21.0966529846191,
-30.6536102294922,12.5925521850586,
20.9050655364990,7.56746101379395,
49.8095626831055,-25.6141929626465,
42.9260711669922,-15.4750595092773,
27.6390647888184,44.4780807495117,
19.6909980773926,76.4438552856445,
14.1702127456665,37.2818222045898,
2.09373807907105,-19.9444255828857,
-10.3575735092163,-27.5000286102295,
-17.0298557281494,-5.35797119140625,
-20.7657012939453,-4.96447801589966,
-27.8305130004883,-20.3431072235107,
-25.3528308868408,-6.63507080078125,
-11.2911243438721,24.6575298309326,
-10.3088331222534,17.1226558685303,
-32.9493980407715,-39.7474098205566,
-46.5933074951172,-83.7284851074219,
-13.2425994873047,-61.5597381591797,
46.4086837768555,-2.60143518447876,
61.0516777038574,24.3827819824219,
7.48897457122803,0.668257772922516,
-53.5919342041016,-33.3439598083496,
-56.2399559020996,-45.4994621276856,
-12.7949409484863,-45.7744522094727,
8.89155292510986,-45.6726799011231,
-19.2005443572998,-43.3828659057617,
-54.7710418701172,-35.5182838439941,
-48.5283203125000,-23.7228126525879,
-13.1928024291992,-11.1412181854248,
9.69187259674072,4.76792669296265,
4.37389230728149,23.3268985748291,
-2.88400053977966,36.4437179565430,
7.45086145401001,36.5854148864746,
28.8495521545410,24.0751056671143,
37.9655227661133,7.08056640625000,
26.3415470123291,-11.8485393524170,
-0.659428477287293,-25.6975536346436,
-23.4677085876465,-14.5984563827515,
-28.1455516815186,19.8153686523438,
-18.0544776916504,43.0814666748047,
-9.80790042877197,25.8435688018799,
-20.5022506713867,-17.0081233978272,
-45.8208427429199,-35.3923225402832,
-61.9032287597656,-16.3204212188721,
-56.5085487365723,8.20960617065430,
-46.5038719177246,6.57217979431152,
-48.7188644409180,-4.90760135650635,
-60.4588088989258,3.04881739616394,
-62.9360771179199,21.3932456970215,
-44.9320602416992,10.1207838058472,
-12.4905185699463,-34.4310646057129,
20.6141567230225,-62.9793205261231,
44.4963798522949,-41.5551757812500,
52.1245574951172,5.97309017181397,
39.4583206176758,33.8622817993164,
18.4092445373535,26.6245651245117,
12.2209596633911,-0.459830611944199,
24.8623828887939,-31.6676025390625,
32.2062339782715,-53.1904487609863,
16.1002655029297,-49.4407691955566,
-11.8553638458252,-19.7992210388184,
-20.5090065002441,5.30206394195557,
-5.19031620025635,-12.2674942016602,
10.6148376464844,-53.0816116333008,
10.6909685134888,-54.1578445434570,
12.3123130798340,0.357310175895691,
29.4483070373535,50.7538604736328,
46.9026603698731,48.9360046386719,
35.6798515319824,19.3626594543457,
5.11862277984619,13.0578422546387,
-4.19032526016235,22.7706317901611,
22.1606502532959,10.1035985946655,
45.9966354370117,-21.5233402252197,
24.0885467529297,-22.7970695495605,
-30.3616695404053,12.4087114334106,
-60.9593811035156,20.0099906921387,
-36.6732254028320,-27.3705501556397,
14.7740631103516,-67.4412307739258,
42.5808067321777,-38.4852714538574,
27.4120521545410,19.3930950164795,
-0.372425079345703,21.9567890167236,
-10.7809247970581,-27.9902667999268,
-1.18213796615601,-43.5031700134277,
7.18109989166260,10.5018386840820,
0.372767329216003,67.3549423217773,
-12.9710874557495,61.8598785400391,
-13.4563474655151,20.3034210205078,
7.93140554428101,11.8135986328125,
30.9026603698730,32.2996215820313,
32.7200584411621,24.8331661224365,
18.2534599304199,-21.3571681976318,
7.58165502548218,-47.0581054687500,
5.12635087966919,-15.1632146835327,
-5.77069711685181,31.2528457641602,
-38.2955818176270,38.3548851013184,
-70.8490142822266,13.8645763397217,
-71.2031860351563,-0.948237836360931,
-48.1733627319336,9.24217033386231,
-37.5178680419922,22.6901397705078,
-41.0282325744629,20.4191493988037,
-26.8946056365967,14.5255022048950,
15.8016490936279,21.1721897125244,
43.5581283569336,25.6406497955322,
21.2435855865479,8.33286094665527,
-17.6217422485352,-22.3850784301758,
-9.98563575744629,-42.4681282043457,
40.8813705444336,-34.9597434997559,
61.4231338500977,-2.87253618240356,
19.6593074798584,31.1455116271973,
-25.7227973937988,31.9331684112549,
-8.04961013793945,-4.30972051620483,
44.9907798767090,-34.9914207458496,
47.4821929931641,-17.8353652954102,
-19.0532913208008,35.8272552490234,
-80.4642715454102,61.4473037719727,
-81.5359268188477,18.4784355163574,
-43.8658561706543,-47.2216873168945,
-20.5874710083008,-56.8538246154785,
-19.0036354064941,-5.38282203674316,
-11.0279493331909,40.9916076660156,
8.11529254913330,43.7299957275391,
13.0697193145752,35.7428550720215,
-8.37953090667725,43.4886512756348,
-33.8352584838867,34.8649978637695,
-41.8112907409668,-18.2297935485840,
-30.8103733062744,-72.2642822265625,
-2.15281462669373,-55.9224586486816,
37.9898300170898,14.9312400817871,
58.5026664733887,44.9486351013184,
27.9799270629883,-1.74444007873535,
-27.9925289154053,-50.4949989318848,
-46.6814880371094,-31.5389003753662,
-6.05301761627197,19.9287204742432,
45.8390579223633,23.1759262084961,
44.5540733337402,-15.1584434509277,
7.16270399093628,-23.2296504974365,
-2.23556923866272,11.3099937438965,
31.7175731658936,33.0532341003418,
56.4046211242676,13.5792579650879,
39.0657844543457,-2.69086480140686,
10.2565469741821,24.0936908721924,
10.0881872177124,50.8705558776856,
24.9235553741455,23.4954910278320,
25.5283412933350,-32.4747314453125,
14.4580717086792,-44.4807167053223,
18.1908569335938,2.24232625961304,
26.3445529937744,46.3647918701172,
3.58867788314819,50.4440956115723,
-48.4926033020020,37.4802970886231,
-78.4180297851563,27.4637050628662,
-51.3263893127441,7.03112792968750,
-1.95269012451172,-31.9963703155518,
12.9330949783325,-59.0209236145020,
-9.17644882202148,-44.1464462280273,
-23.9033737182617,-5.31049013137817,
-6.39794921875000,8.95857810974121,
24.5285243988037,-10.6680269241333,
43.6899795532227,-26.3961219787598,
48.1972351074219,-16.8429737091064,
49.9014701843262,2.71615862846375,
47.3125190734863,14.2661352157593,
31.4016666412354,19.8867549896240,
4.90767288208008,15.2903089523315,
-12.4936122894287,-9.83297157287598,
-11.1500520706177,-38.9212303161621,
1.11650395393372,-39.0456848144531,
7.00723123550415,-6.76694583892822,
-0.877310156822205,12.0202121734619,
-18.5186920166016,-18.0486927032471,
-33.0518341064453,-61.9893264770508,
-33.8989257812500,-58.2250900268555,
-23.9701251983643,-3.08156585693359,
-12.5238656997681,38.8771171569824,
-5.88508272171021,25.4479541778564,
-3.23380351066589,-10.4717683792114,
-1.05429315567017,-20.8516731262207,
1.43781745433807,-8.18266487121582,
-1.46218442916870,-2.60492229461670,
-9.81790828704834,-8.12282848358154,
-22.3482913970947,-0.738293707370758,
-30.6474494934082,22.1197052001953,
-26.0935192108154,28.7642135620117,
-5.85538196563721,1.24771881103516,
20.6075973510742,-36.2488937377930,
40.8793067932129,-47.1893310546875,
45.4378356933594,-27.6796474456787,
37.1389694213867,1.06329345703125,
25.3131332397461,24.8142375946045,
15.7751884460449,41.2285537719727,
10.6925230026245,41.4195976257324,
16.2252635955811,22.5951557159424,
28.2789306640625,1.93272900581360,
30.4366111755371,-0.524560868740082,
10.2477169036865,13.8940925598145,
-19.1833610534668,20.8969020843506,
-27.5013370513916,8.52542781829834,
-0.890081882476807,-5.39847469329834,
28.0345230102539,-0.285632848739624,
17.5023975372314,15.0574836730957,
-30.7179718017578,16.8300304412842,
-64.3438796997070,3.81642460823059,
-40.8192520141602,-3.40236282348633,
17.0213851928711,4.12516975402832,
42.9155921936035,15.3368768692017,
10.8569192886353,13.6439495086670,
-33.2576255798340,5.33854341506958,
-30.3616371154785,5.62393474578857,
7.30924987792969,15.8542633056641,
16.9359130859375,27.1051807403564,
-26.9677467346191,28.6604385375977,
-69.4574584960938,21.2659244537354,
-47.4552764892578,9.04252243041992,
22.0671806335449,-6.82935714721680,
66.2981948852539,-18.6319942474365,
47.1016578674316,-17.9546775817871,
2.60697960853577,-2.92431974411011,
-15.5945329666138,12.8715610504150,
-8.02854347229004,11.8038396835327,
-7.58265876770020,-8.76726055145264,
-19.6713981628418,-36.2725830078125,
-18.4214515686035,-49.8600196838379,
8.18450832366943,-38.8072357177734,
35.4285507202148,-8.48566913604736,
38.8233070373535,21.3118991851807,
16.7237949371338,29.9871654510498,
-15.7957725524902,13.2125253677368,
-34.3159103393555,-12.8567104339600,
-19.7257366180420,-18.5927238464355,
21.4846668243408,5.90898990631104,
52.8893737792969,46.3159523010254,
40.6867523193359,68.7360229492188,
-4.45600080490112,53.8213729858398,
-24.9303112030029,15.5491056442261,
10.1586999893188,-17.6053009033203,
54.9087181091309,-28.8540229797363,
54.6531715393066,-25.5759506225586,
24.1336059570313,-22.2721004486084,
16.5687675476074,-23.6144561767578,
34.8967208862305,-23.3450889587402,
31.2765731811523,-13.4199466705322,
-9.86145782470703,4.17491006851196,
-37.3416862487793,29.4794120788574,
-10.8201017379761,54.0582008361816,
29.0620918273926,58.3971099853516,
22.2826213836670,28.7588863372803,
-15.8435544967651,-16.0989532470703,
-18.8520298004150,-36.3137893676758,
21.8262901306152,-13.2771596908569,
43.0845718383789,22.3947067260742,
12.4686613082886,27.0007495880127,
-19.9855327606201,3.28804063796997,
-6.67524909973145,-8.30993652343750,
23.4563293457031,12.9813184738159,
17.9445571899414,35.7665405273438,
-16.8427200317383,19.3536911010742,
-31.8224449157715,-28.3806819915772,
-15.5024223327637,-58.9510078430176,
-2.89363718032837,-52.3438186645508,
-8.47009277343750,-33.2368125915527,
-0.894273996353149,-29.4001407623291,
35.0816383361816,-34.5963439941406,
60.0508003234863,-19.2370052337647,
46.6575088500977,19.2688674926758,
26.2092437744141,54.0557975769043,
32.6424674987793,61.0218048095703,
45.4751129150391,42.5999565124512,
28.8267784118652,20.2481937408447,
-5.25609827041626,11.1375646591187,
-9.32975959777832,12.4493722915649,
20.1705760955811,11.2997703552246,
36.3629837036133,-2.92132091522217,
15.5667209625244,-29.1767482757568,
-8.23407649993897,-46.8903923034668,
-1.91741085052490,-34.9408035278320,
7.58480930328369,0.597443580627441,
-13.6634187698364,33.3293418884277,
-41.0336837768555,33.1094245910645,
-32.4195747375488,0.0314354896545410,
2.34095382690430,-36.5403518676758,
9.17470169067383,-48.4741859436035,
-21.5910205841064,-36.8265419006348,
-38.9740295410156,-25.5854511260986,
-2.38622093200684,-32.6754379272461,
55.1584663391113,-47.8433532714844,
77.0620040893555,-40.9663810729981,
51.1497573852539,-5.46344041824341,
14.7739562988281,31.8590507507324,
-11.0808019638062,36.3032989501953,
-32.0435638427734,4.53433895111084,
-44.1345367431641,-35.4497451782227,
-22.0438137054443,-50.5157432556152,
30.3022460937500,-32.4109954833984,
71.6712493896484,5.81808757781982,
65.8564376831055,41.5702590942383,
27.8017425537109,47.6489601135254,
-4.72381162643433,16.8430061340332,
-8.17292976379395,-26.5781764984131,
3.50018835067749,-42.0250167846680,
7.70644617080689,-16.7852382659912,
-0.404138445854187,13.9459838867188,
-15.3627634048462,16.1154708862305,
-31.0902481079102,-2.39164566993713,
-38.8015632629395,-10.7692728042603,
-32.4815483093262,-2.55011534690857,
-25.5454959869385,-1.90130114555359,
-28.6603546142578,-18.6946277618408,
-36.1943855285645,-25.2058467864990,
-32.7060432434082,-0.341241240501404,
-26.4782199859619,30.7186603546143,
-39.5718727111816,36.9676437377930,
-70.2228393554688,22.2303676605225,
-81.4267501831055,13.9879455566406,
-39.4335021972656,19.2722511291504,
25.7904262542725,14.8968200683594,
53.1293525695801,-4.42853927612305,
24.7775783538818,-15.7035684585571,
-14.4887609481812,-11.8608207702637,
-20.9087543487549,-18.4942626953125,
-4.21651649475098,-52.0007934570313,
0.730925977230072,-80.6760177612305,
-11.7743368148804,-57.5523185729981,
-18.5852069854736,7.74770116806030,
-13.2610359191895,49.7032470703125,
-14.4799499511719,30.6790103912354,
-30.3306980133057,-15.2207584381104,
-36.8455848693848,-31.4910774230957,
-15.6303920745850,-5.73636484146118,
19.6612663269043,25.4848537445068,
37.1301803588867,25.9218521118164,
28.1632556915283,2.25644516944885,
14.6773843765259,-15.1758060455322,
6.71079349517822,-6.99248886108398,
-0.481546044349670,13.8663024902344,
-8.34572219848633,17.7612743377686,
-13.2857770919800,-10.5282382965088,
-13.6197528839111,-52.4257888793945,
-13.9708700180054,-64.3304977416992,
-19.1372566223145,-26.2508602142334,
-23.1712894439697,28.8771686553955,
-19.9302730560303,43.1707763671875,
-9.61044502258301,3.69558691978455,
7.54902791976929,-44.4478187561035,
36.2112464904785,-52.8673553466797,
61.7872619628906,-20.5535736083984,
52.7134857177734,13.9165296554565,
3.97130298614502,23.6430816650391,
-38.8704185485840,19.1126937866211,
-35.1436157226563,11.8803167343140,
-0.120684623718262,0.298309683799744,
16.6733951568604,-16.5471153259277,
4.24534702301025,-27.0646133422852,
1.97280526161194,-19.4875106811523,
32.5885086059570,-5.87085914611816,
57.4945678710938,-7.65670967102051,
35.8183898925781,-25.3684864044189,
-5.97391891479492,-35.2753257751465,
-9.07309341430664,-25.6606044769287,
25.5873146057129,-6.82882499694824,
40.5073165893555,5.01709938049316,
15.9920444488525,11.1451396942139,
-5.11236286163330,24.3486843109131,
13.5066280364990,45.9749603271484,
38.2999076843262,55.9309158325195,
20.9386615753174,40.4200859069824,
-19.1723346710205,4.97343492507935,
-24.5199680328369,-30.4430961608887,
12.7891349792480,-47.1088562011719,
41.0121459960938,-36.2635231018066,
30.9294567108154,-8.23400497436523,
12.8065013885498,18.4524497985840,
18.7356700897217,32.3692436218262,
24.4560832977295,34.6209754943848,
-3.69898080825806,32.3520393371582,
-37.9327011108398,27.1934661865234,
-24.7133064270020,18.9314918518066,
31.3972854614258,16.4364833831787,
62.8126640319824,34.6637344360352,
24.6130523681641,62.6376495361328,
-44.8463211059570,63.5346603393555,
-68.4690628051758,22.8254718780518,
-25.1410846710205,-19.3658447265625,
28.2831974029541,-17.3973712921143,
33.6103515625000,27.1086959838867,
-10.2738895416260,61.0740585327148,
-57.2323493957520,48.5620040893555,
-68.2261199951172,10.6120471954346,
-45.9639549255371,-22.1529541015625,
-23.0260639190674,-46.2451705932617,
-19.5769195556641,-74.1309814453125,
-22.3392562866211,-88.2493438720703,
-9.87048053741455,-57.5613822937012,
15.0899648666382,0.905944824218750,
27.3264389038086,29.8600997924805,
12.5952959060669,6.01410579681397,
-9.94895839691162,-25.2888393402100,
-10.1988706588745,-15.1898651123047,
16.9395313262939,29.2974376678467,
38.4948806762695,60.3948516845703,
34.7934722900391,52.7405204772949,
15.2335319519043,21.6462421417236,
0.0756206512451172,-10.3991279602051,
-7.93522739410400,-40.5465736389160,
-19.9526824951172,-65.4748840332031,
-32.7980804443359,-69.0564422607422,
-19.5186252593994,-56.4598579406738,
22.4932479858398,-51.1661071777344,
58.4939765930176,-50.3120765686035,
48.7396697998047,-28.7409687042236,
1.42510819435120,18.7668838500977,
-36.6077117919922,41.5061645507813,
-31.8569374084473,5.30551147460938,
-7.02925252914429,-49.6979560852051,
-3.46036982536316,-52.3558158874512,
-26.1820087432861,-3.44377994537354,
-42.3393058776856,25.8757801055908,
-27.4134502410889,-8.97006797790527,
1.98900961875916,-53.6501274108887,
9.18240356445313,-39.0387954711914,
-11.5930490493774,16.1352958679199,
-32.2209129333496,35.5510711669922,
-26.2738838195801,-6.33408117294312,
-6.05841588973999,-54.7339057922363,
-3.18092679977417,-56.6103935241699,
-23.6953296661377,-18.0623035430908,
-39.5002326965332,16.4948787689209,
-19.8326301574707,24.8297290802002,
30.6898536682129,19.1050739288330,
65.5124435424805,15.9410228729248,
51.1652221679688,26.0994434356689,
5.99284219741821,51.3490219116211,
-28.6134185791016,73.1425552368164,
-28.1040115356445,59.1199226379395,
-7.77294206619263,2.72784662246704,
8.75671768188477,-46.1838378906250,
23.2600193023682,-36.5076179504395,
44.6997947692871,14.4835329055786,
59.8543319702148,43.4611320495606,
40.3037719726563,27.2009525299072,
-9.60964012145996,8.05986309051514,
-48.5183639526367,21.7034912109375,
-49.1585273742676,41.0708923339844,
-33.7549934387207,12.9232225418091,
-37.2778053283691,-47.3666076660156,
-51.6676101684570,-72.0124511718750,
-37.6530952453613,-31.8324127197266,
12.9133691787720,22.3655300140381,
58.0592994689941,33.7912864685059,
61.4627380371094,8.34099864959717,
30.4084453582764,-14.4003267288208,
-0.00258708000183105,-11.9847450256348,
-18.0784893035889,4.20918178558350,
-31.4100894927979,20.7469081878662,
-31.9837932586670,22.9293441772461,
-10.6498336791992,4.03633880615234,
17.8631439208984,-30.1387786865234,
25.5332584381104,-54.8418235778809,
13.7642621994019,-48.3804931640625,
15.4983549118042,-29.3551368713379,
45.0086784362793,-31.9718856811523,
75.4966812133789,-45.9300613403320,
74.8557434082031,-26.0268306732178,
53.5532989501953,22.7026100158691,
34.1019744873047,39.1022567749023,
18.2435379028320,-1.37152791023254,
-13.1000480651855,-44.6038284301758,
-45.2682838439941,-31.8122863769531,
-39.0652427673340,7.95527505874634,
7.42945241928101,4.53244686126709,
43.1229553222656,-41.6381530761719,
19.5003604888916,-51.2932701110840,
-38.7825164794922,-1.92272806167603,
-65.1480865478516,33.7164421081543,
-32.0455017089844,0.408576846122742,
17.7247505187988,-49.2921600341797,
27.7654018402100,-29.1016445159912,
-1.41963529586792,39.0049057006836,
-23.6439895629883,60.4415245056152,
-6.31864547729492,4.06078720092773,
30.1735992431641,-50.1431236267090,
55.2640914916992,-33.5316352844238,
60.4089202880859,23.1097126007080,
59.0248260498047,48.6394042968750,
52.1717185974121,34.0651016235352,
28.6539592742920,32.2688293457031,
-10.6408405303955,63.3279647827148,
-40.0977172851563,84.2861862182617,
-33.3618545532227,58.8646240234375,
-6.02091312408447,6.96388387680054,
8.13382816314697,-32.5101737976074,
2.23694157600403,-47.6159820556641,
-1.86998081207275,-45.6853065490723,
16.3929538726807,-38.5128021240234,
39.7823448181152,-31.9006900787354,
35.9236450195313,-23.4303207397461,
4.31719732284546,-9.54331016540527,
-17.2220401763916,9.58781909942627,
-2.95717287063599,25.5121059417725,
21.2186565399170,21.3751525878906,
15.7369813919067,-8.78914070129395,
-19.2816314697266,-33.6118431091309,
-33.0133171081543,-27.2927989959717,
2.19418048858643,-7.89942789077759,
53.7813148498535,-4.20329570770264,
61.8978118896484,-6.66720247268677,
18.3981742858887,15.6980180740356,
-24.6640052795410,57.2174186706543,
-29.0078182220459,66.3655853271484,
-18.6184082031250,19.3468341827393,
-25.0139026641846,-31.1893482208252,
-33.0034561157227,-31.0617179870605,
-8.47402858734131,4.23963165283203,
38.1880645751953,7.95030260086060,
58.0137863159180,-26.1827335357666,
35.7430686950684,-35.5666809082031,
7.23504066467285,12.0130195617676,
0.761706173419952,63.2296104431152,
-4.12931919097900,52.2737350463867,
-26.5614280700684,-0.361169457435608,
-37.7253379821777,-15.6785678863525,
-7.39270401000977,28.1382446289063,
30.4323024749756,75.0052032470703,
16.0051422119141,67.1607055664063,
-39.7784614562988,17.8983020782471,
-66.1782379150391,-25.1234340667725,
-33.5480346679688,-45.4880752563477,
4.18967390060425,-61.8018379211426,
-3.36059474945068,-72.9380111694336,
-26.7613735198975,-56.1748657226563,
-10.7412786483765,-10.0796813964844,
39.3333663940430,29.1649570465088,
65.2573471069336,29.7441787719727,
47.1539573669434,2.73021316528320,
27.8265285491943,-17.1499652862549,
31.2829532623291,-7.60230064392090,
27.6525211334229,21.9581298828125,
-3.94795608520508,45.4262390136719,
-32.8152618408203,51.3190650939941,
-19.2975730895996,40.7995452880859,
22.0407638549805,20.4396820068359,
45.7509384155273,-0.761961102485657,
40.2051086425781,-8.52270889282227,
26.4367008209229,1.20829892158508,
16.7345943450928,22.7634353637695,
-3.89275693893433,40.8029937744141,
-34.6568183898926,37.6092453002930,
-46.9769668579102,4.43766355514526,
-25.8750953674316,-33.8195571899414,
2.06291627883911,-45.5498962402344,
2.66530609130859,-25.7418937683105,
-10.4706029891968,-1.99254679679871,
-4.25838613510132,-3.38631367683411,
25.4768486022949,-20.7168178558350,
43.5917549133301,-19.9894695281982,
24.6127262115479,1.11521852016449,
-13.7977466583252,6.93540763854981,
-30.0841197967529,-20.1280269622803,
-13.5282306671143,-40.9529037475586,
8.63077163696289,-10.5735597610474,
6.88588476181030,44.3822021484375,
-16.2569637298584,55.3277511596680,
-28.0434150695801,1.30927324295044,
-5.15178537368774,-54.7521553039551,
38.8282051086426,-46.1749954223633,
66.7919616699219,5.41935253143311,
50.3012199401856,30.1066875457764,
4.46755504608154,8.73660850524902,
-27.0381870269775,-12.3971347808838,
-19.0885791778564,4.94204807281494,
12.3924932479858,39.5025520324707,
28.5976696014404,51.9126663208008,
6.45505285263062,46.8171043395996,
-38.7476310729981,47.8786048889160,
-68.4271011352539,47.3413162231445,
-60.8004646301270,17.2862129211426,
-26.5475749969482,-36.0177268981934,
6.80769777297974,-63.4158020019531,
14.8781938552856,-36.4172477722168,
-5.41039991378784,16.9404392242432,
-30.8407192230225,37.8319473266602,
-33.1527557373047,12.4491720199585,
-1.20560765266418,-16.9138469696045,
39.9112777709961,-12.2937126159668,
48.3035926818848,22.5493354797363,
16.8637580871582,51.9114990234375,
-23.0227241516113,41.4938583374023,
-35.2770881652832,-4.81756734848023,
-16.9982414245605,-48.3387298583984,
0.673878431320190,-52.3361015319824,
2.98030185699463,-20.5734081268311,
3.50451040267944,10.9007825851440,
11.0024518966675,15.3609504699707,
14.2466468811035,6.31134510040283,
3.00153160095215,13.3899660110474,
-18.4628028869629,36.1403236389160,
-34.5838584899902,36.3382301330566,
-39.0197944641113,0.209789395332336,
-30.9968223571777,-31.3208427429199,
-5.26788949966431,-17.4391269683838,
26.6630821228027,27.6712207794189,
33.7509117126465,50.3565444946289,
-3.26608872413635,25.6835155487061,
-50.5344276428223,-17.9715995788574,
-48.3153610229492,-40.2046623229981,
6.02110052108765,-36.1293640136719,
44.5189056396484,-18.4992256164551,
21.2004432678223,10.3567571640015,
-27.4173259735107,44.2609939575195,
-40.1279487609863,58.9888687133789,
-11.0763731002808,32.4307937622070,
10.8423662185669,-10.6470403671265,
0.491533637046814,-21.0695457458496,
-15.2673740386963,7.68723773956299,
-15.3465242385864,29.6364765167236,
-19.5628643035889,17.2773761749268,
-40.4346885681152,-3.20126962661743,
-48.6156539916992,1.04509294033051,
-24.2668685913086,20.2940464019775,
1.79745435714722,19.1099166870117,
-6.72523307800293,-4.82202529907227,
-24.6305236816406,-12.3654689788818,
-9.79621791839600,11.1462316513062,
17.9492073059082,34.2173957824707,
3.22513341903687,35.2134437561035,
-53.4211807250977,27.9973239898682,
-79.2221145629883,25.6554946899414,
-31.2274208068848,19.4833850860596,
30.9321022033691,4.83691406250000,
35.3439140319824,3.79679846763611,
2.61213684082031,26.3591880798340,
4.66287040710449,37.9719886779785,
40.1785011291504,4.99385070800781,
50.4084777832031,-41.3263549804688,
21.0022239685059,-39.2975463867188,
8.08447837829590,11.6712007522583,
36.2993698120117,39.3837432861328,
56.2640419006348,7.22790193557739,
22.7254161834717,-32.3632621765137,
-23.5598983764648,-20.2454128265381,
-19.9733638763428,16.4194126129150,
17.8642311096191,9.32467269897461,
21.0716438293457,-39.8621978759766,
-24.5910873413086,-58.0188369750977,
-59.5547676086426,-9.29464817047119,
-48.6030845642090,51.6937065124512,
-34.0690002441406,53.6627311706543,
-52.0217742919922,0.745662689208984,
-69.9071807861328,-43.0015792846680,
-48.3256530761719,-46.2831726074219,
-5.53440189361572,-34.3479728698731,
8.24760532379150,-36.3098640441895,
-18.2700920104980,-44.4255180358887,
-42.2914047241211,-39.3383064270020,
-33.6085357666016,-18.9931297302246,
-5.77384948730469,0.454294323921204,
16.9517288208008,5.10915374755859,
37.7116241455078,-5.17649173736572,
59.0350837707520,-12.5866098403931,
65.0651473999023,0.684975981712341,
50.1330184936523,33.7857437133789,
29.3284454345703,60.7283554077148,
13.5225343704224,52.6080932617188,
-9.83052635192871,7.95558547973633,
-43.4219207763672,-32.0654296875000,
-60.2492942810059,-31.9011650085449,
-35.6630287170410,-2.85653185844421,
9.26117229461670,16.0577106475830,
26.1593036651611,7.28097581863403,
7.14181566238403,-11.8110904693604,
-7.27874660491943,-25.6769771575928,
10.6694202423096,-31.1274929046631,
32.0199890136719,-35.2490348815918,
20.2614803314209,-30.4038944244385,
-8.37528610229492,-12.7078275680542,
-8.43351650238037,4.69704008102417,
29.1203899383545,5.27725410461426,
62.8210868835449,-3.17044472694397,
58.3889579772949,2.28851842880249,
22.6058940887451,24.2363357543945,
-10.2781047821045,43.1085662841797,
-26.2930488586426,42.7873458862305,
-32.7072029113770,36.6504211425781,
-36.1109733581543,32.4571914672852,
-38.0220298767090,17.0026721954346,
-37.1833114624023,-19.8392448425293,
-30.8132286071777,-59.8014793395996,
-8.85593318939209,-72.1021423339844,
25.8046321868897,-53.0499038696289,
44.8695144653320,-29.8479099273682,
23.1463356018066,-20.8126850128174,
-20.9382610321045,-15.3154315948486,
-42.5591697692871,0.153535962104797,
-20.1311588287354,13.3648748397827,
15.8013820648193,10.6131153106689,
24.7774753570557,-0.435352087020874,
3.97666072845459,-11.6786403656006,
-9.81255149841309,-24.4005413055420,
-1.74149870872498,-41.1974639892578,
13.5110225677490,-44.3993949890137,
18.6069965362549,-24.6962337493897,
14.6239166259766,1.04416465759277,
9.74178791046143,1.61830484867096,
2.17905926704407,-13.6422948837280,
-8.06098747253418,-4.71491622924805,
-7.09937095642090,32.3111228942871,
11.6397142410278,43.8836250305176,
33.4617881774902,4.99279975891113,
38.0827102661133,-35.9717788696289,
28.6146564483643,-15.1670541763306,
25.8719768524170,49.5771980285645,
34.2023010253906,77.0231018066406,
29.9647617340088,36.1559638977051,
0.308229923248291,-19.9154376983643,
-32.3560600280762,-35.4711074829102,
-36.6423339843750,-27.2740745544434,
-16.0963897705078,-40.1949043273926,
3.81109571456909,-63.2638473510742,
4.15804529190064,-46.1303520202637,
-6.49526691436768,14.3342266082764,
-14.5212287902832,54.3119812011719,
-20.0055904388428,30.4820270538330,
-30.0688800811768,-25.0316905975342,
-37.4775161743164,-51.1851196289063,
-32.2836799621582,-30.8394145965576,
-14.2503767013550,12.4492778778076,
4.36751222610474,44.6841201782227,
11.6795835494995,51.7843704223633,
-1.29888737201691,34.0141944885254,
-30.0375614166260,-0.201342433691025,
-52.6137619018555,-31.0691108703613,
-39.7395629882813,-40.6536788940430,
12.8919572830200,-34.9871635437012,
67.1161346435547,-35.0513420104981,
75.8139419555664,-33.9272651672363,
38.2827262878418,-14.4328718185425,
3.78589868545532,12.4289665222168,
14.2127237319946,15.1879005432129,
51.9198112487793,-1.60812079906464,
63.2334976196289,1.09713137149811,
30.2982749938965,40.4527282714844,
-6.74202108383179,76.6849899291992,
-11.2918624877930,60.1511688232422,
6.23852252960205,3.72797250747681,
5.70718288421631,-38.1708526611328,
-20.4078884124756,-48.0786628723145,
-33.1229476928711,-52.2526321411133,
-4.95582580566406,-56.9514389038086,
39.1061325073242,-30.4642982482910,
46.9328460693359,24.9697227478027,
3.59491419792175,50.2507286071777,
-47.5773162841797,10.8049945831299,
-55.9174575805664,-43.2596397399902,
-18.2021713256836,-36.6990928649902,
24.9032020568848,19.7080726623535,
29.6165390014648,46.9339408874512,
-3.35965490341187,15.3911275863647,
-34.4435958862305,-17.9881668090820,
-36.1708106994629,-5.29186153411865,
-16.2949638366699,19.6971359252930,
4.80670738220215,-0.569741725921631,
19.5901317596436,-41.9906959533691,
36.0944671630859,-37.8930282592773,
47.8668937683106,13.8729896545410,
32.0063514709473,49.4430809020996,
-16.2323532104492,26.8278694152832,
-53.4796142578125,-12.6533832550049,
-36.0535697937012,-19.2406902313232,
16.7614059448242,4.35225820541382,
42.1458206176758,16.9519348144531,
18.4334888458252,3.44599962234497,
-12.7967634201050,-11.6902465820313,
-9.23312568664551,-12.2660646438599,
8.68293666839600,-5.53368568420410,
-3.40480279922485,5.10091876983643,
-39.2449951171875,23.7878761291504,
-53.5886993408203,31.8903427124023,
-30.7475166320801,11.8693504333496,
-11.1587495803833,-22.0930442810059,
-22.0104885101318,-41.6320114135742,
-35.8125419616699,-45.3634414672852,
-22.4500637054443,-56.4357070922852,
2.93702483177185,-77.3997344970703,
14.7729473114014,-77.2686767578125,
23.3898258209229,-38.0643577575684,
48.7261848449707,0.661735653877258,
69.1356658935547,-6.10449171066284,
46.3814964294434,-34.1062088012695,
-4.11287498474121,-30.0008316040039,
-26.5473365783691,-0.651077985763550,
-2.38809084892273,0.157621622085571,
18.4841613769531,-39.2212753295898,
-5.19070577621460,-60.7506256103516,
-36.9528846740723,-20.3028945922852,
-25.8285408020020,35.9701194763184,
7.24746751785278,41.1199760437012,
1.68771553039551,5.02981996536255,
-45.2579460144043,-5.27393531799316,
-68.5662384033203,28.2625427246094,
-32.0283813476563,49.9866104125977,
23.8532428741455,27.1908035278320,
40.2094650268555,1.18700897693634,
10.7578830718994,22.9106140136719,
-24.8228034973145,60.1022148132324,
-40.9892921447754,42.3192634582520,
-39.2788543701172,-27.2839717864990,
-23.0188007354736,-71.4997100830078,
11.5293197631836,-37.3361701965332,
44.8997344970703,36.0833854675293,
50.5286102294922,67.8167877197266,
34.4902915954590,36.0705413818359,
22.0372085571289,-5.38251113891602,
17.5960407257080,-5.98814535140991,
4.05440473556519,22.7321548461914,
-13.7106838226318,38.4426269531250,
-7.07406330108643,21.0966815948486,
25.9256916046143,-2.47868061065674,
43.3244323730469,-1.34493362903595,
9.05511093139648,23.6417694091797,
-42.7144927978516,29.7039813995361,
-51.6413803100586,-11.3069667816162,
-17.4973945617676,-71.0574645996094,
-0.107648074626923,-90.9071273803711,
-23.0712203979492,-51.7323455810547,
-42.9476318359375,4.95927858352661,
-15.1852779388428,21.5931682586670,
37.6791152954102,-9.64016723632813,
61.9273300170898,-37.1862602233887,
47.6879158020020,-25.3340511322022,
28.1778373718262,8.56109523773193,
23.2353458404541,33.1903915405273,
16.2346115112305,46.4355545043945,
-6.27891874313355,61.8259506225586,
-29.8215198516846,70.7876815795898,
-40.5522232055664,44.7857284545898,
-46.3171386718750,-7.41571378707886,
-54.7471733093262,-40.0887145996094,
-49.5725860595703,-25.7649250030518,
-16.0926418304443,4.49157905578613,
20.0410594940186,2.85332918167114,
25.7147045135498,-23.0596885681152,
2.45058822631836,-29.2418613433838,
-16.5646553039551,5.41190528869629,
-11.0194969177246,42.1069335937500,
-0.472455441951752,39.4618415832520,
-7.85985183715820,7.57242155075073,
-23.4005317687988,-18.2104244232178,
-21.4163093566895,-16.8583679199219,
1.87367582321167,6.25240850448608,
20.1714267730713,36.7773094177246,
17.4088420867920,61.2225151062012,
-5.80640411376953,56.9782638549805,
-39.4907226562500,13.4059658050537,
-60.4719810485840,-50.3508872985840,
-47.4870986938477,-87.6329040527344,
1.48951923847198,-76.4586181640625,
45.5012359619141,-38.9933586120606,
40.4402008056641,-6.51805210113525,
-12.7808856964111,11.1918020248413,
-62.5403976440430,12.8336553573608,
-64.1136245727539,-7.01986789703369,
-29.6197681427002,-43.6897087097168,
5.15701627731323,-67.2982254028320,
34.8446960449219,-55.8582153320313,
68.7550201416016,-21.8291702270508,
85.6432876586914,-5.13683176040649,
55.6247100830078,-12.0608959197998,
-5.61078405380249,-10.9466400146484,
-45.2917213439941,17.8354225158691,
-38.0056915283203,49.5801124572754,
-14.3481512069702,52.2604598999023,
-8.90549659729004,35.0362167358398,
-5.22779083251953,27.1806297302246,
20.1091346740723,30.2496013641357,
43.1533393859863,22.3930473327637,
23.2969284057617,-6.15807008743286,
-20.9069938659668,-31.9435653686523,
-29.9544048309326,-36.3865509033203,
6.62266063690186,-33.2278938293457,
27.7591056823730,-39.3244361877441,
-0.684744119644165,-47.7230606079102,
-34.6032524108887,-42.1507759094238,
-15.7074661254883,-29.3304443359375,
27.8294429779053,-30.7869548797607,
28.7760391235352,-47.4592666625977,
-18.2882499694824,-48.5170631408691,
-43.5405464172363,-14.7176074981689,
-7.98105382919312,31.5819530487061,
35.1977500915527,54.2288208007813,
19.2634277343750,33.5877571105957,
-38.3574714660645,-10.9187316894531,
-60.5227050781250,-49.5001907348633,
-19.1129055023193,-66.4628829956055,
30.3452701568604,-64.9580230712891,
32.7694358825684,-52.3649024963379,
0.231372475624084,-33.6152992248535,
-11.6833581924438,-14.5280647277832,
17.3462142944336,-0.575486063957214,
48.1727790832520,-1.02623033523560,
40.1958961486816,-18.7584438323975,
6.23957681655884,-37.4419250488281,
-6.76809835433960,-30.8286323547363,
13.4419040679932,9.89348411560059,
37.2349510192871,53.9816932678223,
30.6965560913086,60.1417770385742,
1.78693318367004,23.9919548034668,
-13.7040576934814,-15.6150436401367,
-3.22396039962769,-17.9414348602295,
8.24454975128174,10.9823627471924,
-3.74204730987549,32.8313140869141,
-25.0971240997314,29.5789852142334,
-30.0939292907715,14.5875062942505,
-16.3993587493897,9.92150402069092,
-2.80528974533081,8.03900718688965,
-1.91475367546082,-5.76051092147827,
-0.691242456436157,-31.0210285186768,
18.1646823883057,-46.5614433288574,
48.7244377136231,-35.4858703613281,
65.6840515136719,-4.51513719558716,
59.5847167968750,26.2482128143311,
39.6445426940918,37.8869056701660,
17.1516780853272,28.0054054260254,
-8.39936256408691,2.92472600936890,
-34.4299087524414,-24.1990108489990,
-40.3875083923340,-41.1220283508301,
-14.4026823043823,-46.5799026489258,
23.7095832824707,-46.9304199218750,
31.1857757568359,-38.5058403015137,
-2.03883886337280,-13.1013221740723,
-33.2684783935547,19.4899063110352,
-23.7821254730225,32.6315612792969,
9.36555099487305,13.4912157058716,
13.6865701675415,-13.0322980880737,
-21.6065654754639,-14.2818813323975,
-52.9445838928223,5.14754915237427,
-48.1932144165039,3.39640259742737,
-28.9651317596436,-38.3619308471680,
-27.6983680725098,-79.8070983886719,
-30.6613445281982,-74.6111679077148,
2.27424550056458,-34.3240699768066,
60.9393043518066,-8.01404190063477,
85.7597427368164,-13.3804626464844,
47.2896499633789,-23.7533302307129,
-11.0447654724121,-15.6927995681763,
-32.1786842346191,2.44885849952698,
-14.4254684448242,14.8358039855957,
3.05117821693420,22.8619308471680,
4.17226934432983,28.1068744659424,
7.99478149414063,14.9104871749878,
17.7580013275147,-20.5768623352051,
14.1825189590454,-43.3996162414551,
-12.5915832519531,-24.4587688446045,
-35.7760963439941,5.43591594696045,
-26.9541816711426,-3.80168795585632,
1.06766402721405,-41.5656013488770,
17.6446800231934,-49.2652511596680,
14.7445755004883,-9.93661594390869,
17.5724086761475,31.7567958831787,
36.7279319763184,37.5405807495117,
45.5031089782715,31.5016975402832,
20.5218334197998,48.2622184753418,
-26.5591030120850,63.2610702514648,
-55.6322708129883,33.0807342529297,
-38.8584861755371,-15.5155735015869,
8.03599548339844,-16.0374450683594,
46.6617050170898,32.9975662231445,
56.9281997680664,55.1915817260742,
43.3597106933594,12.2102527618408,
20.7962226867676,-36.2272605895996,
-3.61399364471436,-20.7584590911865,
-28.3260498046875,30.0988845825195,
-47.3682556152344,42.4090385437012,
-47.2132301330566,5.75586700439453,
-22.5156955718994,-16.1243743896484,
7.64868879318237,14.5621623992920,
12.0194301605225,51.1106376647949,
-18.2328872680664,36.6894340515137,
-50.2307510375977,-15.1779270172119,
-41.4308776855469,-49.7469596862793,
11.8795900344849,-46.2042465209961,
65.1004409790039,-26.2121696472168,
69.6830520629883,-5.41454935073853,
30.8144474029541,16.4238071441650,
-6.77036714553833,35.3933906555176,
-11.0667343139648,39.1641731262207,
5.36178016662598,31.8174877166748,
8.32023143768311,29.8906383514404,
-8.32478427886963,38.0961303710938,
-26.7184123992920,40.1675720214844,
-28.1915512084961,19.3870277404785,
-16.3624572753906,-7.60055351257324,
-6.13551616668701,-20.5785331726074,
-9.00763416290283,-25.1696434020996,
-19.3443527221680,-37.7483940124512,
-26.4092063903809,-49.0872573852539,
-23.0053119659424,-41.0148162841797,
-14.6358880996704,-12.7958889007568,
-11.2289628982544,12.1656312942505,
-13.4012804031372,15.3356294631958,
-7.57680845260620,1.92978942394257,
16.0756645202637,-13.1825485229492,
31.6226959228516,-21.7964229583740,
11.4383068084717,-16.6413478851318,
-30.5059165954590,7.78138542175293,
-46.6673622131348,45.1441078186035,
-17.1117134094238,62.9984207153320,
17.2495727539063,42.2885131835938,
3.68000984191895,7.82258510589600,
-44.2405624389648,0.226439118385315,
-63.7624549865723,21.2624988555908,
-29.2546806335449,38.5699615478516,
15.1242990493774,35.9267501831055,
21.9205856323242,33.4758682250977,
4.42797279357910,45.4393539428711,
7.85496377944946,52.6713752746582,
31.5193614959717,30.2007350921631,
38.8028030395508,-8.49457740783691,
16.8018188476563,-27.3635807037354,
-1.73746275901794,-25.4743995666504,
6.99820899963379,-30.7797298431397,
21.6763439178467,-43.9430465698242,
8.57645606994629,-33.6499099731445,
-25.8388576507568,7.18430900573731,
-46.4756202697754,38.9220504760742,
-35.7347946166992,28.9455184936523,
-10.6373701095581,3.57369732856751,
12.2957801818848,4.00101184844971,
24.7229804992676,24.2198314666748,
12.6492042541504,25.8581809997559,
-21.9358501434326,3.30192947387695,
-52.4318771362305,-0.805946111679077,
-50.5046501159668,25.0479373931885,
-22.3143997192383,40.4325942993164,
-4.12776803970337,10.5644044876099,
-6.45708322525024,-31.8678264617920,
-0.500279426574707,-35.8875083923340,
30.3512878417969,-7.26500082015991,
52.4732704162598,7.24100017547607,
30.6028804779053,-9.00110530853272,
-6.06962490081787,-23.3917102813721,
0.432915806770325,-12.8930263519287,
44.6178894042969,6.61397838592529,
56.8313140869141,7.83383417129517,
6.46609354019165,0.586879611015320,
-53.7371520996094,11.7933816909790,
-56.5178985595703,38.4592132568359,
-9.09557056427002,51.8562088012695,
28.9586162567139,42.4610748291016,
25.5490989685059,21.8476696014404,
1.31414377689362,0.0932804644107819,
-16.1664180755615,-18.1192550659180,
-28.2006034851074,-26.4732227325439,
-33.9356651306152,-27.7104492187500,
-20.7180957794189,-32.6602516174316,
3.76787900924683,-44.8247184753418,
12.2237367630005,-44.0424423217773,
-3.18353056907654,-6.29719400405884,
-6.49929857254028,46.8274345397949,
21.8792114257813,59.5617294311523,
51.5282325744629,14.6694593429565,
40.0511474609375,-28.3168430328369,
3.39067220687866,-10.7660093307495,
-5.62162780761719,35.9520606994629,
23.9181404113770,36.8484153747559,
41.4897613525391,-15.0074911117554,
10.8875141143799,-48.6330375671387,
-27.9142913818359,-11.4450807571411,
-19.6798057556152,50.0356712341309,
27.0457172393799,59.1848526000977,
53.6813087463379,11.2767753601074,
30.8917446136475,-32.7294616699219,
-7.84988784790039,-30.7105121612549,
-26.5460624694824,-5.84225511550903,
-26.4565010070801,12.7366685867310,
-32.0476608276367,21.5416526794434,
-45.4247589111328,25.8418312072754,
-45.9833297729492,11.4269456863403,
-19.3187656402588,-25.2799510955811,
21.1998310089111,-49.6843719482422,
55.8707313537598,-32.9471206665039,
69.2109832763672,10.8938055038452,
53.1271705627441,41.3192405700684,
18.8686447143555,39.2769966125488,
-5.83679294586182,21.3115634918213,
-9.83985614776611,3.67268109321594,
-10.0910949707031,-20.1873817443848,
-17.8923797607422,-46.8536109924316,
-17.1561927795410,-48.8365516662598,
7.98178577423096,-15.4947338104248,
43.2600173950195,25.7828464508057,
48.2189216613770,41.1400375366211,
20.9428062438965,29.9445686340332,
10.7899074554443,13.9379472732544,
43.2121391296387,5.45085096359253,
73.6677017211914,-5.53033971786499,
45.8113861083984,-16.9672164916992,
-14.2709188461304,-14.1949014663696,
-36.6580162048340,5.36867046356201,
-3.00263786315918,19.3935050964355,
21.8507099151611,4.34885644912720,
-5.02599859237671,-22.7156028747559,
-37.8198242187500,-33.0819015502930,
-12.5049457550049,-17.0430927276611,
53.0696983337402,4.44990587234497,
80.5763854980469,11.9221506118774,
40.3626976013184,4.32513093948364,
-11.9403438568115,-11.4529209136963,
-21.0277214050293,-28.9437980651855,
-2.76662778854370,-43.2495155334473,
1.07697618007660,-51.0784912109375,
-5.85719347000122,-49.3796615600586,
8.66763496398926,-42.3687362670898,
46.8181114196777,-28.6333312988281,
66.5199661254883,0.163878440856934,
45.0566291809082,41.1988754272461,
-1.61337065696716,68.8633804321289,
-32.7761993408203,66.6711807250977,
-30.1018676757813,47.8523406982422,
-3.82520198822022,36.1751289367676,
28.1123847961426,34.6835098266602,
45.0896301269531,30.2968025207520,
32.1533012390137,27.3651065826416,
3.04501724243164,40.2574806213379,
-4.33787727355957,61.6287384033203,
20.3215408325195,56.6693267822266,
45.8110656738281,11.6006431579590,
38.3101768493652,-30.0925235748291,
4.21366834640503,-22.8321857452393,
-26.4581756591797,15.0584678649902,
-40.4508132934570,22.1543636322022,
-50.9730377197266,-17.3475131988525,
-58.9813957214356,-54.2681503295898,
-41.8209838867188,-46.1258163452148,
3.70882511138916,-11.7030458450317,
37.1965599060059,17.1333999633789,
27.4937610626221,36.7651405334473,
-4.24382734298706,60.8657836914063,
-16.7682800292969,68.7425918579102,
-6.56251525878906,30.9943237304688,
-1.92962443828583,-32.2374343872070,
-7.47034978866577,-52.8799781799316,
-3.25558352470398,-11.0606412887573,
11.8268299102783,39.1696624755859,
4.46430873870850,38.7867813110352,
-35.4067459106445,-1.47193682193756,
-64.3910827636719,-32.1092033386231,
-37.2427406311035,-36.2646980285645,
19.1955738067627,-28.5301513671875,
43.0031738281250,-11.8984565734863,
21.8315219879150,19.1126022338867,
1.07718288898468,48.4262161254883,
11.4477243423462,41.7144393920898,
22.9419021606445,2.25496387481689,
3.66580057144165,-16.8770751953125,
-23.4261245727539,14.1588153839111,
-13.9743652343750,57.0041732788086,
26.7793445587158,56.9015884399414,
47.8299484252930,19.7228794097900,
24.3291854858398,-1.65211701393127,
-10.2209281921387,13.8640270233154,
-12.9351196289063,39.4428291320801,
4.10395526885986,43.2326545715332,
-2.56639957427979,25.7126693725586,
-37.9312896728516,2.85146379470825,
-60.8103523254395,-18.2365226745605,
-38.3658638000488,-36.0326271057129,
13.0331935882568,-33.8115806579590,
41.1685523986816,-7.23121881484985,
18.4108943939209,17.7072849273682,
-21.7481155395508,9.82434654235840,
-29.5398941040039,-25.0722064971924,
3.78558826446533,-48.3673286437988,
35.2717781066895,-44.3338470458984,
19.9043235778809,-28.6236820220947,
-32.7147026062012,-19.9910163879395,
-64.5158767700195,-23.3269081115723,
-39.9358520507813,-28.6589393615723,
6.38231658935547,-29.2423553466797,
13.5302238464355,-18.7002105712891,
-25.5248603820801,5.23730325698853,
-57.0738143920898,36.3956298828125,
-35.1937065124512,48.4584693908691,
14.3654346466064,32.8267631530762,
28.3722000122070,9.80539894104004,
-12.6701278686523,0.392065554857254,
-55.3447265625000,-8.56503772735596,
-46.8254470825195,-39.5501365661621,
0.507684707641602,-72.0271911621094,
29.4536628723145,-64.6859893798828,
10.1178359985352,-17.9093551635742,
-24.8963623046875,22.7367877960205,
-31.7708663940430,22.9216880798340,
-15.5079956054688,8.34883975982666,
-14.0488872528076,18.5618495941162,
-31.9073905944824,41.6034393310547,
-38.9288558959961,30.3632144927979,
-12.0580387115479,-14.0674381256104,
22.0091571807861,-45.6537704467773,
22.6379203796387,-41.1136512756348,
-6.55670595169067,-28.3474349975586,
-18.6249408721924,-33.7877426147461,
5.27215480804443,-31.6296215057373,
33.1177940368652,-0.434577941894531,
25.3947811126709,29.2722816467285,
-8.79674625396729,12.8089799880981,
-27.3278770446777,-29.3680419921875,
-13.8347845077515,-36.8245277404785,
-0.865056514739990,6.77733039855957,
-16.4788284301758,40.2235260009766,
-48.2603225708008,10.9244689941406,
-62.6919364929199,-45.8270568847656,
-47.8037414550781,-66.1012191772461,
-23.6111278533936,-43.9721565246582,
-11.4671068191528,-26.2950248718262,
-13.7848548889160,-36.7558364868164,
-14.6121053695679,-55.6754112243652,
-2.05538845062256,-57.9154548645020,
22.0120563507080,-43.6442527770996,
45.1986351013184,-27.0056076049805,
57.3617362976074,-11.4347877502441,
53.8365440368652,-5.66290664672852,
42.6745948791504,-17.7335491180420,
34.7345008850098,-36.2455177307129,
32.5051689147949,-22.6785964965820,
31.7654895782471,28.3293476104736,
26.4885978698730,64.6570358276367,
16.9529514312744,41.6478805541992,
5.54693126678467,-9.04034900665283,
-4.40151977539063,-23.5604038238525,
-13.8866291046143,4.11327648162842,
-25.8726844787598,23.2676353454590,
-39.4786605834961,1.55662655830383,
-39.2279396057129,-25.6170806884766,
-13.6504678726196,-16.7906112670898,
27.0903263092041,14.0630874633789,
52.1050338745117,23.3120956420898,
44.1797370910645,18.6571941375732,
21.4557266235352,33.5040473937988,
13.7988576889038,64.8021926879883,
19.4776954650879,70.9262771606445,
9.89313793182373,40.8488311767578,
-19.8070049285889,14.8140716552734,
-31.3998031616211,13.5683441162109,
1.94984555244446,10.3059730529785,
49.3899116516113,-15.0279455184937,
53.4898338317871,-32.3148269653320,
5.16553974151611,-9.74498081207275,
-43.8593101501465,27.3807163238525,
-45.5536041259766,22.0248508453369,
-14.5512504577637,-25.0403327941895,
1.53493237495422,-47.1051216125488,
-3.58716034889221,-12.0822029113770,
-1.44928455352783,33.8129768371582,
23.5987071990967,39.9441032409668,
45.8615570068359,15.4474868774414,
35.9652252197266,-5.55952310562134,
7.51215171813965,-16.5045108795166,
-5.53267860412598,-30.2243022918701,
-2.58753347396851,-42.7807426452637,
-7.93779468536377,-38.9670028686523,
-23.0293254852295,-34.2323341369629,
-17.1239452362061,-48.7544441223145,
22.6513328552246,-63.9357986450195,
57.0074806213379,-35.4764976501465,
35.9926795959473,30.2539272308350,
-23.4114952087402,63.4302291870117,
-50.3001747131348,27.8024921417236,
-14.4958095550537,-23.2519569396973,
38.0446128845215,-27.6919918060303,
44.0525741577148,-0.626497149467468,
6.59972810745239,4.48744630813599,
-13.6728363037109,-16.7429809570313,
14.5076007843018,-16.4122848510742,
58.3414802551270,28.4950866699219,
63.7857208251953,74.0907058715820,
29.0757865905762,79.6438903808594,
-3.48068046569824,62.1711120605469,
-4.51665210723877,50.3118476867676,
11.0783290863037,33.9713249206543,
16.2009773254395,-0.442966938018799,
0.411440610885620,-24.5566539764404,
-22.9426116943359,-5.84946393966675,
-33.8915557861328,25.7668094635010,
-35.4720497131348,18.0841140747070,
-34.0058898925781,-19.7675762176514,
-28.1949501037598,-29.7639293670654,
-19.6314277648926,5.05899190902710,
-18.5049285888672,27.3946208953857,
-33.5227394104004,-7.73626279830933,
-53.1525421142578,-53.7374420166016,
-46.8694610595703,-39.0172042846680,
-8.67298030853272,22.5805053710938,
24.1343917846680,55.7570419311523,
5.76872491836548,37.7171096801758,
-45.9566268920898,19.8611202239990,
-65.6910171508789,28.6084671020508,
-15.7504415512085,28.9308223724365,
60.0452766418457,-3.00721216201782,
88.6814346313477,-33.3444023132324,
54.3685188293457,-20.8454055786133,
4.50125360488892,13.6250839233398,
-20.7046413421631,21.8495483398438,
-18.1852817535400,4.55307340621948,
-5.94419527053833,4.94694805145264,
5.47794246673584,24.6805763244629,
9.79445171356201,19.2471733093262,
-4.37943458557129,-16.8233585357666,
-33.7070198059082,-32.8652839660645,
-51.7392234802246,-10.3324537277222,
-44.3751068115234,4.08906698226929,
-28.9376506805420,-24.3944778442383,
-25.8891162872314,-50.7968864440918,
-22.4705562591553,-20.9337120056152,
-4.81578779220581,40.6991233825684,
6.32599973678589,59.8500823974609,
-15.0159854888916,23.2162303924561,
-47.1336860656738,-2.65125250816345,
-43.6499671936035,23.5144710540772,
-0.777389049530029,55.7091255187988,
18.9400177001953,44.5226860046387,
-22.2514934539795,15.4007196426392,
-77.1675415039063,13.4198150634766,
-74.8265075683594,27.0145626068115,
-23.3813152313232,11.0758876800537,
7.01499509811401,-35.2372436523438,
-12.3996257781982,-67.0529403686523,
-29.7311382293701,-65.9461059570313,
5.63574314117432,-54.9044151306152,
62.8437423706055,-50.3325691223145,
74.1372528076172,-34.8549728393555,
28.6584205627441,-1.61760354042053,
-18.3845329284668,14.5511941909790,
-20.1691875457764,-9.43072605133057,
10.8529710769653,-32.0917778015137,
34.9923286437988,-11.5462455749512,
41.7828140258789,30.5541343688965,
47.0096054077148,41.4956512451172,
52.3925399780273,19.2912464141846,
39.8505287170410,6.93319368362427,
6.39967536926270,25.4371833801270,
-18.3612766265869,45.1945343017578,
-13.9795722961426,41.1890144348145,
6.40037631988525,29.2362518310547,
9.62436771392822,28.0447559356689,
-14.4277315139771,18.8641681671143,
-38.2240829467773,-17.4932689666748,
-34.9659652709961,-45.6442337036133,
-11.1738281250000,-22.8616752624512,
8.60114002227783,31.6939735412598,
20.3194274902344,53.9165725708008,
33.7267112731934,20.4891242980957,
45.6342010498047,-17.8988151550293,
36.4678878784180,-15.5511741638184,
-0.130316078662872,7.96950626373291,
-29.8817386627197,4.52726745605469,
-21.1499977111816,-29.8227424621582,
16.3475608825684,-50.9610214233398,
33.2350311279297,-36.0474967956543,
5.12685489654541,-11.8938570022583,
-35.7230682373047,-11.7246913909912,
-44.6419944763184,-23.2224903106689,
-22.6915893554688,-15.3535614013672,
-10.2741470336914,12.7391881942749,
-30.6764354705811,25.7237205505371,
-59.1767616271973,0.845971584320068,
-53.8291320800781,-40.6475105285645,
-15.0719318389893,-58.0887298583984,
22.2360820770264,-33.9083061218262,
35.5487785339356,-0.724304437637329,
37.9243392944336,7.06042385101318,
38.0787353515625,-6.67158269882202,
25.1943721771240,-14.5874567031860,
-5.18689632415772,-2.93089866638184,
-29.1575756072998,8.45556640625000,
-16.0430850982666,-3.00000190734863,
18.0237083435059,-30.3310527801514,
21.2844333648682,-37.6061859130859,
-15.0923919677734,-12.5046606063843,
-39.1590385437012,18.1598358154297,
-9.31536674499512,19.3467540740967,
42.6386146545410,-0.989759802818298,
48.0780868530273,-7.59639310836792,
4.32852888107300,18.0909004211426,
-22.4555339813232,46.8366546630859,
7.18712997436523,36.9853057861328,
44.6276855468750,-6.77507352828980,
24.1895599365234,-41.0350303649902,
-40.8160095214844,-38.4444351196289,
-71.5218429565430,-20.1820793151855,
-33.7947540283203,-18.0286178588867,
21.4573001861572,-29.0057926177979,
26.1957702636719,-27.4854564666748,
-17.6203975677490,-8.45411109924316,
-51.5597915649414,7.59638786315918,
-41.1040344238281,11.7937135696411,
-8.30883598327637,22.0237598419189,
14.3150596618652,46.8577957153320,
20.0886936187744,65.9605712890625,
23.4603519439697,56.2561607360840,
31.0805644989014,28.6203231811523,
30.5970516204834,8.96274375915527,
13.1457386016846,2.94683933258057,
-10.0109939575195,-6.14551544189453,
-17.7904434204102,-17.5865688323975,
-2.71038007736206,-12.2381248474121,
21.4662761688232,7.56175422668457,
34.3477287292481,18.9894695281982,
24.1700630187988,8.47185039520264,
7.37035083770752,-4.58249664306641,
1.18102288246155,2.34270071983337,
2.31517720222473,20.8448963165283,
-6.98727798461914,26.1979904174805,
-31.8824558258057,17.3660240173340,
-51.4873962402344,16.2242050170898,
-37.6061820983887,27.3938751220703,
7.18006420135498,34.8510551452637,
46.9471855163574,28.3891754150391,
50.5359649658203,19.6275863647461,
20.2708263397217,11.3623971939087,
-11.2045392990112,-6.16536283493042,
-23.9269123077393,-33.3449401855469,
-25.9988040924072,-44.9888381958008,
-33.9395866394043,-23.3114967346191,
-45.1732215881348,14.1929807662964,
-41.7512588500977,32.8536224365234,
-16.8655662536621,22.9440155029297,
10.4925212860107,9.68505382537842,
16.4670028686523,9.60531711578369,
1.24145674705505,8.27474975585938,
-14.8648223876953,-4.88404273986816,
-14.3428754806519,-16.4400539398193,
-1.53213667869568,-13.2480325698853,
1.30388987064362,-1.38870692253113,
-11.4140958786011,1.07031726837158,
-31.1114234924316,-5.45830869674683,
-35.9478836059570,-8.96879196166992,
-17.0073471069336,-9.91090202331543,
10.3615875244141,-15.6035518646240,
17.7086467742920,-17.4731483459473,
-7.20518493652344,1.99658322334290,
-41.7249145507813,33.8804206848145,
-50.3891868591309,37.5749740600586,
-18.3065490722656,-5.72488927841187,
23.8234100341797,-58.2162246704102,
35.7924842834473,-66.6844940185547,
11.2722253799438,-31.3567848205566,
-14.2086629867554,-3.00894737243652,
-3.24986505508423,-16.7628002166748,
40.5595169067383,-45.7330093383789,
77.1322555541992,-44.0786514282227,
77.0926895141602,-4.64506101608276,
52.0356674194336,32.7553558349609,
31.8648052215576,37.4517860412598,
29.4923458099365,20.0620594024658,
31.2852153778076,12.1602287292480,
17.3513278961182,18.5780372619629,
-9.50166797637940,19.4742813110352,
-30.5522632598877,0.743518471717835,
-32.0790596008301,-23.4385795593262,
-16.9989318847656,-37.1450920104981,
-1.51627564430237,-40.3623008728027,
1.65163218975067,-45.1894836425781,
-7.47099685668945,-51.4257583618164,
-17.8434543609619,-36.5459823608398,
-17.5793228149414,0.0503435134887695,
-10.7891016006470,32.3195953369141,
-12.2180957794189,33.2802124023438,
-25.0797634124756,15.4003181457520,
-30.4042758941650,10.2302904129028,
-16.2082862854004,27.8152236938477,
7.64560651779175,46.1777954101563,
14.6353378295898,43.0116691589356,
1.44364380836487,32.0105743408203,
-6.26274013519287,36.6309700012207,
6.45724105834961,49.5266761779785,
23.6183452606201,40.9781761169434,
22.2251491546631,4.06560707092285,
3.88333845138550,-35.6536483764648,
-9.11639308929443,-53.1158638000488,
-6.90064859390259,-52.9704513549805,
-4.48378849029541,-53.2350769042969,
-14.0119628906250,-53.3800582885742,
-23.8142433166504,-30.6891403198242,
-19.5811252593994,10.0569076538086,
-6.30215978622437,27.4040298461914,
-1.10669672489166,-3.74717283248901,
-6.11189365386963,-53.9944877624512,
-5.55312871932983,-62.3625679016113,
12.2133903503418,-16.8428058624268,
32.9663314819336,25.7887630462647,
32.8409767150879,12.9743347167969,
12.6835613250732,-32.4791069030762,
0.992800712585449,-38.5080299377441,
14.3568143844605,14.2482976913452,
33.6963539123535,64.2746887207031,
25.9087009429932,49.4919013977051,
-5.76851320266724,-12.9529314041138,
-23.8956470489502,-46.0685272216797,
-4.80508708953857,-17.6760597229004,
29.1955509185791,34.8375091552734,
41.2413063049316,51.0299339294434,
28.5100498199463,23.9453716278076,
16.2471218109131,-12.7795066833496,
10.3555784225464,-29.7640991210938,
-2.07437920570374,-20.0542736053467,
-19.1716136932373,8.41076660156250,
-16.1005420684814,40.0563964843750,
12.7104883193970,55.4173812866211,
34.6972236633301,36.3066520690918,
25.4768619537354,-5.02766704559326,
5.90867948532105,-32.8490486145020,
10.8635931015015,-33.6194038391113,
31.7183780670166,-28.0776062011719,
31.2402305603027,-39.2487869262695,
6.56231594085693,-60.7296028137207,
-2.80842018127441,-59.4619483947754,
21.6208572387695,-18.2998466491699,
39.2657356262207,33.4958229064941,
10.0012207031250,52.4545707702637,
-40.7952995300293,27.4643135070801,
-61.4327583312988,-13.4084997177124,
-37.5085258483887,-29.9911308288574,
-5.54930400848389,-7.71170902252197,
4.37868595123291,26.9053249359131,
3.92845845222473,35.1259193420410,
9.84430313110352,6.12040805816650,
16.5476570129395,-30.5846252441406,
8.62344837188721,-34.9824333190918,
-7.74552297592163,-11.4734001159668,
-18.9178504943848,5.89418888092041,
-25.8658866882324,-4.92206764221191,
-31.3086051940918,-24.9178466796875,
-20.0044364929199,-26.2983169555664,
18.2037601470947,-9.51138210296631,
59.5721817016602,-5.61678504943848,
61.6428756713867,-20.2480010986328,
24.7310619354248,-29.0244331359863,
-9.14964580535889,-19.0361442565918,
-3.94737696647644,-0.766021966934204,
27.6615161895752,8.60854339599609,
44.1404991149902,8.61527442932129,
36.8482589721680,5.07260990142822,
27.8047409057617,-10.2849264144897,
26.3037128448486,-40.6870918273926,
18.9486713409424,-55.9412117004395,
-0.801955580711365,-29.4143714904785,
-20.6554889678955,16.3595409393311,
-24.1623802185059,24.7960796356201,
-6.51047277450562,-19.1923732757568,
27.3792648315430,-60.9523010253906,
61.2082252502441,-43.3050460815430,
68.7754669189453,12.7011423110962,
32.2910270690918,37.7397270202637,
-22.3178787231445,6.10949230194092,
-44.5475654602051,-31.5092887878418,
-11.4111700057983,-23.0641994476318,
30.5917854309082,17.1348361968994,
25.3249511718750,31.2772388458252,
-16.6825447082520,-0.958197355270386,
-34.8920249938965,-36.2262191772461,
-8.21282958984375,-29.8473167419434,
21.9311504364014,8.48420333862305,
21.1393203735352,29.8776130676270,
9.18999481201172,14.1702604293823,
22.1876220703125,-15.3336992263794,
51.4089279174805,-27.4382572174072,
58.0584869384766,-15.8736066818237,
38.2717285156250,-0.301290333271027,
27.4823398590088,-1.04050707817078,
37.0617752075195,-12.3931169509888,
38.2038230895996,-24.9279747009277,
9.81697654724121,-36.5765151977539,
-22.8060054779053,-47.4737815856934,
-26.4043045043945,-50.5720558166504,
-11.4165058135986,-39.4199180603027,
-2.02321219444275,-16.3101272583008,
1.93235135078430,0.150493264198303,
17.3803424835205,-6.26731491088867,
37.2051963806152,-25.7584114074707,
34.9038734436035,-23.2966976165772,
8.40686702728272,8.78790855407715,
-8.73587894439697,37.1201477050781,
0.724299550056458,21.0818157196045,
12.4628162384033,-28.9429626464844,
-1.12902796268463,-62.4848518371582,
-24.6674365997314,-49.8107833862305,
-29.6537609100342,-20.6367340087891,
-18.9863452911377,-18.3255348205566,
-16.4144935607910,-36.5566024780273,
-19.7677783966064,-40.2290573120117,
-3.35780310630798,-17.6381473541260,
35.6959991455078,1.83611273765564,
60.2421531677246,7.29260063171387,
41.0492553710938,18.1967544555664,
-0.136657238006592,47.8704490661621,
-18.1866397857666,67.9872360229492,
-2.86127424240112,48.7730789184570,
16.2237358093262,13.1778907775879,
14.7106504440308,9.24495506286621,
0.770533859729767,46.2472496032715,
-11.2377538681030,73.6360549926758,
-20.4823894500732,49.0396003723145,
-28.3246517181397,-12.8227024078369,
-31.7377395629883,-58.4127807617188,
-29.6874599456787,-59.6965408325195,
-22.8508968353272,-28.3440971374512,
-18.3888645172119,11.2441768646240,
-17.8661289215088,41.8795433044434,
-19.9209842681885,49.6827278137207,
-23.4390525817871,35.5090141296387,
-25.0530872344971,12.0981445312500,
-14.6105651855469,-5.24563884735107,
2.21139049530029,-14.8168783187866,
1.28891348838806,-29.8210926055908,
-25.8225097656250,-53.4353637695313,
-42.4242782592773,-70.8812789916992,
-14.4671764373779,-67.7379608154297,
35.3955268859863,-46.1124343872070,
40.7810134887695,-16.6697311401367,
-16.4029064178467,17.5979843139648,
-69.9901733398438,43.0095367431641,
-54.8253364562988,36.0073585510254,
6.29648494720459,-3.35054445266724,
30.6708850860596,-40.8085975646973,
-6.75406789779663,-33.6882476806641,
-40.7789192199707,10.3163824081421,
-13.3134756088257,35.3529891967773,
48.1557846069336,11.6185626983643,
77.5176239013672,-26.3977279663086,
59.6809310913086,-24.5649375915527,
37.1205024719238,16.6205749511719,
39.4882621765137,48.3900909423828,
50.5278015136719,41.1157989501953,
46.6289634704590,17.7634925842285,
26.1406021118164,8.82380485534668,
4.62872695922852,8.74864292144775,
-11.9416341781616,-7.21244955062866,
-17.4541378021240,-34.4810600280762,
-1.33067536354065,-42.2226943969727,
32.3784561157227,-15.6869239807129,
47.5196609497070,24.2559757232666,
22.9858779907227,45.7568016052246,
-17.6621398925781,43.4813880920410,
-34.4844284057617,36.4464187622070,
-24.3419952392578,32.5627861022949,
-12.3315277099609,25.1463680267334,
-13.0742874145508,7.62074756622314,
-16.1198348999023,-15.0771045684814,
-11.0318708419800,-25.3523597717285,
-15.7879772186279,-12.2683134078980,
-40.3365631103516,16.4753265380859,
-61.7854652404785,30.5980491638184,
-55.0662193298340,10.9095115661621,
-29.5310001373291,-25.9240322113037,
-15.6455554962158,-42.2011070251465,
-19.5188159942627,-18.2157688140869,
-25.4647884368897,19.0158939361572,
-28.2169609069824,20.3910446166992,
-36.1774482727051,-19.3028888702393,
-44.3525962829590,-57.8954277038574,
-33.6830978393555,-60.2372474670410,
-3.29075336456299,-34.2666740417481,
16.2461910247803,-16.7060394287109,
0.490114212036133,-21.3625946044922,
-24.9913730621338,-38.4679794311523,
-18.4533443450928,-54.0228500366211,
18.8980827331543,-57.9728736877441,
45.2722358703613,-41.1260871887207,
42.8546485900879,2.15659928321838,
35.3842658996582,50.0491828918457,
39.6228485107422,61.6970787048340,
39.1609725952148,22.0326633453369,
11.5185661315918,-32.2017517089844,
-24.6978473663330,-49.9314460754395,
-35.3302497863770,-28.5760002136230,
-16.5351047515869,1.45897781848907,
1.02726721763611,14.8419780731201,
1.47400641441345,6.39014959335327,
-0.254448711872101,-19.1248531341553,
7.74525547027588,-44.7762298583984,
9.71667385101318,-45.5458183288574,
-1.13890480995178,-3.61829900741577,
-4.78129529953003,49.2676887512207,
11.1833715438843,58.3370208740234,
25.0001621246338,12.0186548233032,
13.2872085571289,-26.0995693206787,
-12.5320873260498,-9.12909412384033,
-27.4631309509277,25.9214286804199,
-27.6975383758545,5.56533670425415,
-29.7013549804688,-62.9939460754395,
-29.4173316955566,-96.4056091308594,
-4.52804565429688,-47.9853668212891,
34.4135742187500,26.2566871643066,
37.6306610107422,40.6296424865723,
-2.22914195060730,-6.42261266708374,
-30.2710838317871,-44.0661430358887,
-3.23988842964172,-30.3197708129883,
41.7923049926758,6.67577981948853,
45.9443244934082,30.2893962860107,
10.8071517944336,40.3037490844727,
-8.58207130432129,51.6556930541992,
2.86097383499146,51.8488273620606,
2.87284541130066,28.4109039306641,
-28.2467155456543,2.28092527389526,
-47.2991142272949,2.41862487792969,
-18.5287036895752,25.6049365997314,
15.2821340560913,39.9035072326660,
0.240380167961121,24.4496135711670,
-48.5245704650879,-6.46821975708008,
-66.9768295288086,-20.0895195007324,
-42.7108078002930,-15.4146842956543,
-28.0240345001221,-8.75091743469238,
-43.0703544616699,-14.8714265823364,
-46.6391754150391,-39.9987525939941,
-1.27107143402100,-69.8827743530273,
57.6161460876465,-71.5267257690430,
69.1477050781250,-23.1278228759766,
31.0553436279297,44.5792541503906,
0.816772460937500,71.3052978515625,
4.57671451568604,30.4876384735107,
10.6617355346680,-23.5641098022461,
-12.0515556335449,-27.8375453948975,
-46.5178451538086,13.4024343490601,
-58.2287445068359,28.8436203002930,
-38.9621849060059,-18.7576694488525,
-4.37062168121338,-79.4812850952148,
32.0688095092773,-82.8989715576172,
59.4924125671387,-24.7900543212891,
71.3248672485352,35.5709915161133,
59.3390846252441,57.1224441528320,
31.8707256317139,52.0130538940430,
5.48206233978272,49.3482398986816,
-14.0882759094238,50.7639732360840,
-33.4975776672363,36.6612701416016,
-50.1380043029785,4.40032863616943,
-45.8538665771484,-30.0537929534912,
-23.9899597167969,-51.4555206298828,
-3.11736869812012,-57.1084938049316,
7.48657369613648,-51.9375152587891,
12.6564445495605,-39.8159942626953,
12.3049087524414,-23.8517894744873,
-4.87567329406738,-8.25578689575195,
-37.7632789611816,10.4044532775879,
-55.1888313293457,33.6162948608398,
-32.9572029113770,49.2328872680664,
10.1615562438965,46.1076202392578,
32.8141250610352,28.4672775268555,
23.5791873931885,15.9365520477295,
13.3890380859375,20.5956878662109,
12.1804943084717,27.8947486877441,
-2.40287971496582,17.3947048187256,
-36.1151390075684,-7.85482597351074,
-53.7822456359863,-18.4836254119873,
-22.2571086883545,0.621108770370483,
27.5467720031738,31.1792907714844,
41.1063270568848,44.3977012634277,
12.8081455230713,29.8746604919434,
-11.1561679840088,8.33562088012695,
-6.05425691604614,-0.445536792278290,
-2.19177842140198,9.11081695556641,
-26.4648513793945,23.6282424926758,
-48.0320014953613,26.0061473846436,
-25.1021347045898,7.80186939239502,
23.2349395751953,-23.4012527465820,
38.7210159301758,-47.8457794189453,
12.3314666748047,-46.7223815917969,
-10.3448266983032,-25.3159465789795,
4.71739816665649,-4.24211263656616,
38.0926551818848,1.59834313392639,
51.0035629272461,-0.418034881353378,
36.3329696655273,2.43386578559876,
12.0172729492188,11.1467514038086,
-9.98747920989990,17.7107563018799,
-24.3958511352539,20.9905281066895,
-18.0187377929688,26.8026103973389,
12.3532886505127,32.4006805419922,
41.3945693969727,20.4668159484863,
40.8910865783691,-11.9267454147339,
26.7482109069824,-38.3937988281250,
32.4397087097168,-34.4071884155273,
50.7358932495117,-2.27395915985107,
39.4813880920410,24.7487220764160,
-11.4318675994873,22.6768379211426,
-53.4446372985840,5.13333511352539,
-38.2279243469238,-5.52309417724609,
15.3233270645142,-9.23849964141846,
42.3889999389648,-20.4419231414795,
17.6192607879639,-34.8629074096680,
-18.7768707275391,-30.2750530242920,
-24.0165252685547,-0.782006502151489,
2.90017676353455,21.5902671813965,
33.3141593933106,8.94479084014893,
48.3989715576172,-17.4382190704346,
48.9895172119141,-9.57993412017822,
38.8800277709961,39.1138877868652,
23.3915157318115,76.8797225952148,
9.86297225952148,56.1526908874512,
2.78749728202820,-2.76536059379578,
-3.39124584197998,-30.0905475616455,
-15.9760389328003,3.33976030349731,
-32.9456253051758,46.5986938476563,
-39.4294738769531,32.2046089172363,
-30.5084018707275,-35.4303894042969,
-20.6252689361572,-84.7573623657227,
-19.1040401458740,-63.9408226013184,
-18.0813980102539,0.0188597440719605,
-7.74155521392822,39.1817474365234,
6.25074434280396,26.5608177185059,
11.8366537094116,3.16134834289551,
3.20024991035461,10.4369020462036,
-8.32641410827637,32.4205818176270,
-16.9277935028076,31.2912845611572,
-25.4025764465332,7.93504953384399,
-32.0112762451172,-6.30435657501221,
-24.8527412414551,-0.325120627880096,
1.24185776710510,-5.39094161987305,
27.4032707214355,-34.9664726257324,
30.2331752777100,-51.0162811279297,
9.15121841430664,-17.1200218200684,
-14.8008975982666,34.4150276184082,
-28.1404170989990,43.1023674011231,
-31.5369911193848,4.55740404129028,
-28.5731372833252,-26.8737964630127,
-11.4849796295166,-13.1674385070801,
20.8913230895996,10.1691465377808,
54.1016731262207,-1.40648031234741,
67.2260742187500,-29.9380683898926,
60.7971496582031,-26.4704246520996,
45.7770919799805,10.9814777374268,
27.0773906707764,33.6432876586914,
2.26094722747803,16.5107898712158,
-20.1177864074707,-7.67803812026978,
-21.7806282043457,4.32547473907471,
-3.93094754219055,38.2342643737793,
12.4447307586670,48.3321495056152,
10.0593442916870,15.9161930084229,
-4.39544248580933,-25.1684703826904,
-14.6020565032959,-39.7215538024902,
-16.5843944549561,-30.1639938354492,
-16.7414360046387,-15.6664676666260,
-10.0324764251709,-10.4923801422119,
11.3133563995361,-9.76943492889404,
41.5037727355957,-1.28420066833496,
58.3418502807617,13.1665353775024,
50.5330047607422,21.8842067718506,
32.8397979736328,16.4102897644043,
16.5833950042725,-3.80843496322632,
1.21285116672516,-29.2218227386475,
-16.8214225769043,-47.6674118041992,
-30.2661666870117,-55.2840003967285,
-33.9450111389160,-53.7597427368164,
-29.2725028991699,-37.7188415527344,
-23.1826190948486,-0.340378463268280,
-16.9773349761963,46.0431175231934,
-8.00919246673584,68.2169265747070,
-6.82529449462891,43.2454299926758,
-22.7945289611816,-9.77576637268066,
-41.5109825134277,-39.7636489868164,
-39.5148124694824,-21.9227466583252,
-22.2644901275635,11.0835075378418,
-16.0475063323975,11.3321132659912,
-25.5070896148682,-25.0629425048828,
-17.9035186767578,-50.9990081787109,
15.8212633132935,-30.8807468414307,
39.1800765991211,13.7678527832031,
13.6351661682129,33.0321044921875,
-34.9542617797852,9.21339035034180,
-42.6769218444824,-25.7942790985107,
4.22804927825928,-34.2306442260742,
46.9338111877441,-20.5896472930908,
38.3442306518555,-8.99856758117676,
6.53825283050537,-4.84911155700684,
5.17254877090454,6.21905565261841,
33.5698852539063,33.4619941711426,
46.9981803894043,54.6569252014160,
26.3939228057861,45.6756477355957,
-3.77441835403442,12.3117532730103,
-21.1723155975342,-19.7940082550049,
-31.2720260620117,-28.2858047485352,
-40.5087623596191,-10.8274478912354,
-33.8340911865234,18.9510269165039,
-4.59469079971314,39.4588546752930,
21.8313350677490,39.3526840209961,
20.9156436920166,15.4703960418701,
9.56412506103516,-14.0440835952759,
18.0715274810791,-21.8221282958984,
35.4496803283691,-1.67031359672546,
27.7528953552246,28.7789726257324,
1.14215040206909,38.6331787109375,
-4.12514495849609,16.8695640563965,
28.1052589416504,-18.4522247314453,
61.5406112670898,-33.4191589355469,
58.5634498596191,-9.91603279113770,
28.0234031677246,26.6105613708496,
7.44507503509522,41.4215202331543,
1.70407116413116,28.4708728790283,
-10.4012498855591,20.6984844207764,
-22.8663520812988,42.4579391479492,
-12.4025039672852,68.0327911376953,
17.3667240142822,52.2420196533203,
27.8442726135254,-3.34520626068115,
10.0611782073975,-48.5827560424805,
-0.933389663696289,-47.9422912597656,
13.9673032760620,-28.8705406188965,
27.8318881988525,-28.6731986999512,
11.0042896270752,-33.2692909240723,
-17.3614234924316,-8.55817031860352,
-13.0720729827881,39.9775886535645,
20.5031013488770,62.5427513122559,
36.6811637878418,39.9686470031738,
21.0762710571289,7.43271493911743,
10.4752130508423,-0.293356001377106,
25.8336944580078,6.52853965759277,
39.5976943969727,0.0480237007141113,
29.9665203094482,-16.3014640808105,
16.8741416931152,-18.1880779266357,
27.3399600982666,-10.6915683746338,
35.9576873779297,-12.4569578170776,
2.63809728622437,-20.9263248443604,
-51.6481666564941,-7.44185256958008,
-59.4734344482422,26.1464309692383,
-5.17165184020996,47.2962799072266,
44.5451812744141,40.2025947570801,
27.1844234466553,31.9359989166260,
-33.9641532897949,41.4437103271484,
-68.2128372192383,45.3684272766113,
-54.9666671752930,13.8124885559082,
-37.5121078491211,-39.5787925720215,
-39.7937316894531,-62.7246932983398,
-29.9943332672119,-40.5272445678711,
21.2557659149170,-11.4942979812622,
78.7245483398438,-14.3369703292847,
82.3864669799805,-37.8824577331543,
25.7762718200684,-48.1144638061523,
-24.6564216613770,-32.5129508972168,
-14.4036302566528,-6.08218097686768,
28.3639736175537,10.2761011123657,
35.6815376281738,9.08640575408936,
-5.46484947204590,-6.84578609466553,
-40.7478103637695,-20.1507663726807,
-21.7778244018555,-16.0206165313721,
27.8709163665772,6.61111545562744,
45.2230873107910,27.7293930053711,
10.7332000732422,30.6286563873291,
-26.2037715911865,21.1483993530273,
-25.2068519592285,20.5324783325195,
-3.59225273132324,30.6374244689941,
-5.90117454528809,26.7539443969727,
-32.6337394714356,3.61695575714111,
-42.1276588439941,-18.3074207305908,
-8.51496696472168,-19.3726215362549,
39.3894119262695,-3.98664426803589,
52.4158592224121,11.1071472167969,
22.9251251220703,20.1636676788330,
-10.7871198654175,28.3506450653076,
-18.6874561309814,29.3004665374756,
-11.2651195526123,12.0750646591187,
-14.6596946716309,-10.8385782241821,
-31.3224258422852,-14.7376585006714,
-37.3165245056152,2.40691614151001,
-15.0686197280884,9.45102119445801,
13.1521835327148,-16.5320377349854,
17.7266273498535,-49.9059906005859,
-1.80292773246765,-52.4044494628906,
-15.7260475158691,-26.6514282226563,
-1.05115032196045,-12.4105882644653,
32.3393783569336,-26.6848373413086,
56.7911300659180,-46.7760658264160,
58.5444793701172,-39.8234634399414,
43.1875534057617,-11.1121425628662,
18.5084857940674,5.76465129852295,
-9.93045234680176,-3.75522637367249,
-26.2137088775635,-23.0977916717529,
-13.8123416900635,-34.3059997558594,
24.8054008483887,-26.9530506134033,
56.1457595825195,-0.630964994430542,
55.7013282775879,27.3419170379639,
31.9021263122559,26.6712856292725,
15.4230928421021,-5.30381298065186,
16.8742580413818,-28.0187091827393,
23.6964988708496,-3.12904882431030,
22.0462646484375,43.0871734619141,
9.78448009490967,43.6517524719238,
-7.99916505813599,-19.3445339202881,
-26.8442382812500,-70.4031829833984,
-34.8993949890137,-44.4499511718750,
-19.4241733551025,18.2175292968750,
12.1168212890625,25.2000236511230,
22.8125381469727,-30.0954971313477,
-8.16590499877930,-58.5195808410645,
-52.8485870361328,-15.0317935943604,
-65.8018035888672,35.3612442016602,
-38.9369201660156,16.2977008819580,
-12.2297677993774,-42.4445381164551,
-15.1335744857788,-52.1121864318848,
-29.8925590515137,0.858051657676697,
-20.6695728302002,38.7011756896973,
14.9136810302734,8.38681983947754,
47.0090446472168,-44.3719329833984,
55.5769157409668,-49.2633857727051,
50.1111335754395,-7.84874343872070,
44.6597480773926,23.5590877532959,
35.8775215148926,16.8512744903564,
16.8186511993408,-11.7494859695435,
0.0498152077198029,-39.7848930358887,
4.94429588317871,-56.4816017150879,
28.1521854400635,-50.7112007141113,
44.5872116088867,-21.8496665954590,
33.1723442077637,7.15978622436523,
-2.28032445907593,7.85859966278076,
-35.0298843383789,-13.0221138000488,
-39.6571426391602,-16.9597129821777,
-21.0779571533203,13.6808013916016,
-6.34887123107910,37.6575736999512,
-13.0888872146606,18.3599777221680,
-28.5791110992432,-20.0170593261719,
-23.6331596374512,-22.2285804748535,
4.94079065322876,19.6027221679688,
21.6355304718018,61.7429924011231,
0.926434993743897,60.0115661621094,
-33.3338584899902,17.8363857269287,
-33.4809570312500,-24.7077350616455,
0.137058734893799,-42.5538597106934,
21.8289051055908,-37.4185867309570,
6.27988958358765,-22.7796440124512,
-15.1798458099365,-15.2910623550415,
-2.27505850791931,-25.0276908874512,
32.2949600219727,-46.1289901733398,
40.7471771240234,-53.1620025634766,
15.2974672317505,-35.3792953491211,
-8.17600917816162,-19.8600215911865,
-10.4902296066284,-32.1803321838379,
-13.6600685119629,-54.0612258911133,
-34.1860771179199,-43.3450851440430,
-41.7013893127441,4.28523969650269,
-4.88159561157227,42.1728515625000,
44.9459571838379,31.4142208099365,
50.6006584167481,-7.58410453796387,
8.73529815673828,-23.9245128631592,
-25.3753890991211,-14.3531513214111,
-11.7255725860596,-11.5078010559082,
25.9087066650391,-21.5128707885742,
37.7592010498047,-17.9495868682861,
15.6777572631836,8.74792671203613,
-8.88826656341553,20.7735519409180,
-10.1458377838135,-6.06815338134766,
10.2790546417236,-39.9344329833984,
40.4363594055176,-40.1516036987305,
58.5505409240723,-12.7345256805420,
42.0570945739746,-0.482488334178925,
-8.73919486999512,-12.1578769683838,
-50.6254081726074,-12.5440607070923,
-38.9386177062988,16.8341884613037,
12.8939180374146,44.9654922485352,
47.2285041809082,36.7652854919434,
31.2012481689453,9.20602512359619,
-3.07567858695984,-2.90338921546936,
-5.10675811767578,6.81636238098145,
23.9954586029053,22.9506874084473,
39.2880821228027,32.4177818298340,
23.1922492980957,33.6091308593750,
3.75617551803589,18.9944229125977,
3.51023507118225,-15.2725114822388,
18.0635757446289,-44.0032997131348,
31.6786537170410,-38.1625976562500,
40.3474044799805,1.86772251129150,
46.1236877441406,35.0877761840820,
36.6875648498535,39.9720611572266,
5.98718643188477,38.5487632751465,
-27.0351142883301,49.9570312500000,
-41.3966598510742,52.1247673034668,
-34.6471519470215,22.9931354522705,
-23.8079586029053,-11.2510643005371,
-12.7277803421021,-10.2221717834473,
10.5232982635498,26.2145538330078,
35.3987045288086,50.5627250671387,
29.5283756256104,33.4475250244141,
-14.1990299224854,-6.31130456924439,
-53.4882202148438,-36.6332855224609,
-47.2735061645508,-56.0564765930176,
-2.77478408813477,-69.4800262451172,
30.5839748382568,-61.6813316345215,
22.0963516235352,-21.2475624084473,
-12.0566539764404,15.2647647857666,
-41.0318298339844,9.67672729492188,
-51.8055458068848,-19.4859237670898,
-45.6544151306152,-21.3723678588867,
-23.7831192016602,15.7572040557861,
-1.75053322315216,48.9670906066895,
-6.88713264465332,47.7723922729492,
-41.3875579833984,27.5836544036865,
-70.4250183105469,16.5931415557861,
-59.6748237609863,4.00591087341309,
-26.0978374481201,-24.5375785827637,
-13.5674943923950,-40.1223678588867,
-30.0405445098877,-11.2858028411865,
-40.9323272705078,26.9780635833740,
-22.9195652008057,11.8937263488770,
-2.31270670890808,-46.0125122070313,
-12.0491170883179,-68.0102233886719,
-35.0706672668457,-25.8211765289307,
-28.1859493255615,15.3076601028442,
9.01795959472656,-4.60728263854981,
37.4968223571777,-46.2053260803223,
31.4901256561279,-28.4284629821777,
6.04273700714111,46.5816192626953,
-13.1343250274658,90.9327239990234,
-18.1244697570801,59.0662040710449,
-13.1306991577148,9.01537322998047,
1.90001857280731,1.09723627567291,
17.3015003204346,22.8814315795898,
15.6590967178345,29.5372524261475,
-9.45149993896484,16.7723560333252,
-32.1828384399414,8.85542106628418,
-31.0725784301758,2.29284787178040,
-24.3067741394043,-21.4738616943359,
-40.5798568725586,-42.0175743103027,
-60.7788200378418,-26.0547046661377,
-39.2419319152832,13.5125379562378,
20.0816402435303,22.1133804321289,
60.6049270629883,-13.9550447463989,
42.8284988403320,-35.4451942443848,
-5.31598806381226,-1.35102653503418,
-26.0088253021240,38.8431510925293,
-9.08430290222168,13.8734989166260,
12.9256067276001,-55.2294692993164,
18.0991954803467,-84.3426666259766,
13.7933368682861,-35.5684356689453,
7.40962409973145,29.3004608154297,
-7.10930633544922,34.4546394348145,
-20.6728935241699,-17.7739276885986,
-13.0846242904663,-55.8803291320801,
8.00645637512207,-42.6279830932617,
7.12667179107666,0.0320479869842529,
-23.3238525390625,32.1701889038086,
-45.1895141601563,40.6788520812988,
-27.5190620422363,35.4311370849609,
11.9496879577637,24.0574417114258,
34.0258979797363,13.4000921249390,
30.4561786651611,14.2195167541504,
29.2155399322510,27.4702033996582,
30.4584140777588,31.6607341766357,
9.94342041015625,7.69042158126831,
-27.0716419219971,-33.5387573242188,
-39.6579551696777,-59.3429870605469,
-10.2658920288086,-54.7234001159668,
21.6095695495605,-48.3421821594238,
17.0307235717773,-66.4478836059570,
-6.74138689041138,-89.1941146850586,
-10.7133407592773,-71.9739379882813,
6.54172182083130,-12.7833328247070,
9.59073638916016,35.7259635925293,
-11.0738668441772,27.6072216033936,
-19.0871028900147,-10.8313159942627,
13.1522617340088,-18.2177066802979,
59.0961151123047,22.6244201660156,
71.3583602905273,55.0447311401367,
40.3956260681152,33.2096099853516,
-4.31248903274536,-16.0871658325195,
-27.3377189636230,-29.6834812164307,
-17.8982219696045,3.92464542388916,
15.1445426940918,36.5510482788086,
47.6552581787109,29.5579452514648,
48.2204093933106,3.38900828361511,
6.40236949920654,3.86802673339844,
-47.5972862243652,29.5285358428955,
-67.7985458374023,40.2756881713867,
-34.9066886901856,13.1119804382324,
18.3194541931152,-19.4686622619629,
42.0366973876953,-16.1911849975586,
24.7526626586914,23.6488437652588,
-2.46734213829041,58.5079154968262,
-6.21149826049805,54.3989067077637,
10.2803144454956,21.5807075500488,
23.5908451080322,-3.04898953437805,
15.6750001907349,-1.82758998870850,
-1.00431656837463,11.7422981262207,
-8.30980014801025,17.7288322448730,
-5.48044204711914,11.8712415695190,
-9.39488124847412,5.82102537155151,
-28.8994712829590,7.78515768051148,
-53.1598587036133,10.7643384933472,
-58.8742599487305,7.68751859664917,
-42.3047561645508,-1.03173482418060,
-14.9753026962280,-9.89824485778809,
8.91843032836914,-14.1451568603516,
24.6954574584961,-7.63028335571289,
34.9147186279297,9.41428661346436,
40.1426200866699,25.0850658416748,
36.0874061584473,23.7368202209473,
25.7911281585693,-1.87842965126038,
17.5931053161621,-31.2918300628662,
19.5531616210938,-37.5227432250977,
30.4893112182617,-17.9064350128174,
38.6167068481445,7.20424079895020,
31.7739353179932,16.4581336975098,
9.49162769317627,7.36916875839233,
-17.3247985839844,-6.32010650634766,
-35.6811828613281,-10.5069665908813,
-42.0690841674805,-4.20181274414063,
-41.7025299072266,5.28261804580689,
-41.7838897705078,7.68913269042969,
-40.3197059631348,-0.435179769992828,
-36.4907684326172,-7.42076826095581,
-31.2575950622559,0.410746276378632,
-28.5222377777100,19.5832939147949,
-26.8020687103272,22.8106746673584,
-22.3498744964600,-4.54003334045410,
-13.1502590179443,-39.4031715393066,
-8.76265525817871,-44.1469688415527,
-9.85632324218750,-17.4588527679443,
-10.3871965408325,3.57942819595337,
-2.73534345626831,-12.6114130020142,
8.24470901489258,-47.0161361694336,
10.4463872909546,-56.2669296264648,
-5.41236686706543,-26.5254173278809,
-30.9609355926514,9.68486976623535,
-41.5873603820801,22.3451690673828,
-25.9538345336914,9.08341026306152,
5.74049949645996,-12.8266506195068,
25.0691623687744,-35.0005035400391,
22.3159580230713,-50.9421310424805,
15.4091567993164,-48.8926811218262,
34.7945327758789,-26.5111732482910,
71.6114349365234,-3.47027301788330,
82.6348648071289,-0.504463195800781,
48.3008880615234,-13.5757503509521,
1.71756553649902,-22.3682880401611,
-11.6495895385742,-21.5946712493897,
4.15705299377441,-30.8546752929688,
6.83401584625244,-55.4151268005371,
-18.8377227783203,-64.3515090942383,
-36.3777809143066,-32.0057716369629,
-14.7352972030640,21.1567516326904,
19.5102958679199,58.7019805908203,
23.3269081115723,66.3923645019531,
4.85175037384033,53.6340713500977,
11.2181921005249,30.5274848937988,
47.6436462402344,2.69943928718567,
65.8027267456055,-14.2227602005005,
32.3844642639160,-3.59997415542603,
-18.4840240478516,19.7445793151855,
-32.9704055786133,18.5033264160156,
-12.3018760681152,-7.96320438385010,
3.47374057769775,-14.7364635467529,
-4.28678226470947,18.7318134307861,
-12.7922668457031,47.9715270996094,
-4.01890182495117,28.2993125915527,
9.88625335693359,-15.8301334381104,
18.6475963592529,-23.0787220001221,
30.6148834228516,6.12328624725342,
46.9019355773926,20.7745666503906,
39.4059410095215,-2.21242523193359,
-7.80938720703125,-19.1070632934570,
-57.7342491149902,4.19428539276123,
-61.1779251098633,27.6667289733887,
-19.4004344940186,1.72600698471069,
15.9335269927979,-50.9697227478027,
10.4783210754395,-61.1408996582031,
-14.6757450103760,-16.9356861114502,
-20.1318073272705,22.9618568420410,
-2.20725727081299,19.3982563018799,
10.3660764694214,-2.54444408416748,
-0.783291935920715,-6.24755144119263,
-21.9510898590088,-5.58559226989746,
-33.4713249206543,-29.6142635345459,
-20.6572132110596,-66.7762680053711,
16.0382690429688,-72.4759674072266,
57.4635276794434,-30.5612659454346,
77.3539123535156,21.9949607849121,
59.4157333374023,45.6334190368652,
20.3977642059326,38.3533096313477,
-6.04178190231323,20.3455410003662,
-3.67062854766846,-0.135277926921844,
18.8588027954102,-18.7750892639160,
38.6013793945313,-24.4190731048584,
47.0950736999512,-9.36904335021973,
40.8429298400879,16.5115470886230,
10.4140567779541,35.7670249938965,
-37.7136688232422,37.5151214599609,
-73.6961975097656,22.7377834320068,
-67.6343154907227,1.22514367103577,
-23.1139755249023,-16.9686508178711,
22.1121387481689,-25.6020240783691,
39.0666427612305,-20.3512020111084,
34.4841079711914,-7.32359790802002,
31.0219383239746,1.32976257801056,
32.3151245117188,9.24275016784668,
32.4722862243652,23.6620998382568,
27.3823394775391,36.5396347045898,
29.4516696929932,34.3373107910156,
36.8878784179688,15.4742221832275,
31.1353797912598,0.553290307521820,
3.64530086517334,-2.03751349449158,
-26.9089298248291,-9.73085689544678,
-35.3957939147949,-32.4154510498047,
-14.5038690567017,-47.5074157714844,
15.8062515258789,-19.0352554321289,
33.5294952392578,42.4115142822266,
32.0007743835449,80.1508941650391,
23.0274829864502,58.5633850097656,
21.3846111297607,9.96499824523926,
31.7282848358154,-14.2892904281616,
42.4608230590820,-6.97683620452881,
33.1654281616211,1.16061341762543,
1.21761488914490,-9.13475990295410,
-31.3324127197266,-25.1992683410645,
-31.5069274902344,-29.6259899139404,
-3.93533229827881,-29.8337688446045,
15.8333225250244,-26.5931911468506,
5.80408382415772,-6.53838109970093,
-16.8276023864746,27.9625911712647,
-22.4296493530273,43.4602851867676,
-1.78519296646118,16.4368019104004,
26.1955814361572,-22.6248264312744,
39.5278930664063,-16.1982154846191,
32.6858863830566,36.5314407348633,
7.13051605224609,66.3901672363281,
-24.1237716674805,32.2408866882324,
-29.8689136505127,-25.5025234222412,
6.42989540100098,-30.9292030334473,
50.3685684204102,19.6301517486572,
48.7985649108887,52.5240821838379,
-1.61370968818665,16.3391799926758,
-36.1376838684082,-47.9402313232422,
-7.18429899215698,-58.8808441162109,
45.2646980285645,-5.40436983108521,
44.5754470825195,48.8418884277344,
-9.17274093627930,43.3864173889160,
-39.6606178283691,-4.98212718963623,
0.0876245498657227,-33.1579742431641,
56.6599617004395,-12.5461044311523,
45.9928703308106,29.6268501281738,
-25.5062961578369,47.9311637878418,
-76.3175125122070,37.6793327331543,
-54.2924270629883,28.4911079406738,
0.508056402206421,30.8338165283203,
21.0155906677246,29.4499149322510,
3.44822883605957,8.67201614379883,
-4.87883949279785,-21.8813037872314,
18.2284431457520,-28.3293018341064,
40.7599372863770,2.44142532348633,
21.1811332702637,42.5604324340820,
-32.8175659179688,56.1590843200684,
-70.6364746093750,39.5411415100098,
-60.9408454895020,11.3110218048096,
-20.8892631530762,-11.9800262451172,
16.0286560058594,-30.0288486480713,
33.4143562316895,-43.6895561218262,
35.9248657226563,-34.4604110717773,
32.6826438903809,4.73698186874390,
21.4149398803711,44.1577415466309,
-0.700560808181763,42.8847579956055,
-17.7550849914551,-6.72160148620606,
-18.4768791198730,-58.6647682189941,
-8.30236721038818,-67.8512878417969,
0.0636719912290573,-36.5347023010254,
1.85095024108887,-4.63529586791992,
5.74724483489990,1.40565013885498,
16.7738475799561,-3.43339896202087,
25.6857395172119,4.05131673812866,
19.6631946563721,23.0603275299072,
2.84697175025940,30.9206905364990,
-7.94540977478027,10.7757797241211,
-7.76995468139648,-24.9090747833252,
-6.25927209854126,-47.2023086547852,
-16.9344062805176,-39.2774353027344,
-36.1432418823242,-5.28990888595581,
-43.5360832214356,29.4792366027832,
-25.2915897369385,39.9549674987793,
7.79427337646484,20.5464401245117,
30.2063255310059,-9.19185352325440,
26.5835475921631,-27.6122035980225,
6.41029071807861,-30.1282863616943,
-11.1857357025146,-28.1180210113525,
-17.3083839416504,-31.1160087585449,
-15.7949686050415,-34.5337677001953,
-13.3459920883179,-28.7301025390625,
-10.0922861099243,-14.6476469039917,
-8.18218994140625,-0.0598560571670532,
-8.83671188354492,14.2009105682373,
-9.93832492828369,31.7631206512451,
-8.11648464202881,41.5955543518066,
-3.05302548408508,28.2068424224854,
-1.87503004074097,-6.37334108352661,
-3.12170147895813,-34.9992713928223,
1.04881632328033,-28.5181846618652,
16.6819152832031,7.89111900329590,
30.8534927368164,44.4875602722168,
28.8928127288818,58.8056793212891,
12.5544137954712,52.7732505798340,
-11.6976833343506,40.2843093872070,
-40.2465133666992,23.8112411499023,
-61.5538978576660,9.22252845764160,
-52.7457199096680,3.64532184600830,
-7.65729427337647,10.6251087188721,
39.0686340332031,13.1869592666626,
41.4805297851563,-0.938912868499756,
-4.03986024856567,-25.1345539093018,
-46.1498870849609,-32.8671417236328,
-48.5410003662109,-16.5623455047607,
-32.6933708190918,4.00302267074585,
-32.5630722045898,8.99935150146484,
-37.0874023437500,1.85035431385040,
-17.1284770965576,-2.71353578567505,
15.1060037612915,-6.97993469238281,
17.9199256896973,-22.8953399658203,
-9.91808795928955,-47.3177032470703,
-22.0153293609619,-59.2939910888672,
6.96024274826050,-51.3089981079102,
36.4670906066895,-44.4890060424805,
23.8870429992676,-53.0855941772461,
-5.95674562454224,-61.7978782653809,
-0.113114833831787,-41.1139907836914,
39.1321411132813,9.06209850311279,
52.8619689941406,51.9467544555664,
16.0719718933105,57.5517272949219,
-22.7549552917480,36.4868927001953,
-17.3912792205811,21.2569427490234,
12.6916732788086,23.8253593444824,
19.2298393249512,25.2419052124023,
-4.77616596221924,1.89900040626526,
-20.4815006256104,-40.7309112548828,
-3.78305506706238,-71.2167510986328,
23.5526371002197,-60.9015541076660,
34.6811027526856,-14.8162317276001,
32.5569953918457,25.3112869262695,
33.8128967285156,31.3115215301514,
41.0657272338867,8.84845352172852,
44.8994483947754,-7.09572649002075,
46.7334060668945,0.230291545391083,
49.2110900878906,17.6610450744629,
42.6439170837402,18.4378604888916,
13.0405750274658,1.87951707839966,
-23.7254772186279,-14.2908220291138,
-37.6769332885742,-18.9091243743897,
-15.1436424255371,-10.0977134704590,
14.8104763031006,10.0998678207397,
13.7245788574219,33.4382247924805,
-19.6708049774170,39.1223335266113,
-41.7248115539551,12.0604963302612,
-22.6127052307129,-35.6922111511231,
17.7381649017334,-59.6624832153320,
37.8640022277832,-42.7633361816406,
22.1105022430420,-11.3362913131714,
1.24451673030853,-4.44119167327881,
8.56913757324219,-23.9114074707031,
40.5591087341309,-35.0903015136719,
52.3381576538086,-18.5013732910156,
22.3956813812256,6.26076650619507,
-27.2845973968506,14.7037525177002,
-49.5527801513672,12.1012077331543,
-35.6529884338379,16.3848724365234,
-19.0822105407715,27.9811992645264,
-32.3420066833496,26.4218864440918,
-62.0166740417481,0.974652767181397,
-60.6296157836914,-33.1840400695801,
-14.8724575042725,-56.2757301330566,
31.6927185058594,-59.0804481506348,
34.4220466613770,-45.7132720947266,
5.83921623229981,-26.2386322021484,
0.234029233455658,-7.35604333877564,
41.7952156066895,-1.43102753162384,
87.4140472412109,-5.61196327209473,
80.8956909179688,-4.07627677917481,
22.6688156127930,16.7480945587158,
-35.2161483764648,39.7167778015137,
-59.6354179382324,39.8502044677734,
-55.7991409301758,11.3790969848633,
-43.7214393615723,-23.2375507354736,
-25.8763465881348,-34.3189964294434,
6.41442680358887,-15.4845991134644,
35.1576347351074,15.7369108200073,
36.6168251037598,34.7955932617188,
13.9077253341675,26.7668685913086,
-2.37728857994080,-4.38344526290894,
3.38443636894226,-35.6737556457520,
10.6634988784790,-45.4210739135742,
-3.68982291221619,-38.1261940002441,
-24.4998855590820,-41.9624938964844,
-15.4253158569336,-62.8083496093750,
26.7219200134277,-70.1267547607422,
55.6694602966309,-41.3004646301270,
39.9574203491211,-0.201843261718750,
1.06659555435181,9.86894035339356,
-12.8061895370483,-13.8794307708740,
16.0979003906250,-30.9684505462647,
49.0565185546875,-13.7919378280640,
52.5191116333008,15.1897296905518,
30.0640068054199,23.6081256866455,
10.4955492019653,24.8414363861084,
3.50928139686584,40.9244194030762,
-2.82241821289063,55.1329803466797,
-16.5113620758057,35.3437194824219,
-25.5726490020752,-8.50593090057373,
-17.5211296081543,-24.7327880859375,
2.95733642578125,2.18636560440063,
13.6808691024780,31.5973930358887,
-2.88695859909058,19.1517105102539,
-35.6440811157227,-16.2303352355957,
-51.2881660461426,-34.1120452880859,
-28.1636562347412,-30.8709316253662,
22.6996078491211,-32.8121871948242,
61.0621337890625,-37.7272720336914,
58.5421180725098,-12.6116485595703,
29.6805648803711,42.0520706176758,
11.5356273651123,69.7384567260742,
16.5938205718994,39.8499031066895,
34.4908409118652,-9.25385093688965,
45.6448020935059,-23.1568241119385,
45.6695289611816,-4.98789215087891,
33.7742538452148,-0.196514546871185,
11.9474430084229,-28.3602504730225,
-10.2865858078003,-54.8881072998047,
-15.2319793701172,-44.2308883666992,
1.02495861053467,-7.18839359283447,
15.5540924072266,25.6442661285400,
9.07813739776611,43.7619705200195,
-6.12033605575562,49.7457427978516,
-2.99564456939697,44.6324729919434,
17.9773159027100,35.8209419250488,
23.5010986328125,39.9916114807129,
-4.30494976043701,58.2323799133301,
-41.7665824890137,61.3711967468262,
-55.2348365783691,32.2107162475586,
-43.6172981262207,-3.09721732139587,
-30.9555091857910,-3.22939395904541,
-27.0853862762451,28.2505035400391,
-19.6787986755371,42.3231506347656,
0.122499585151672,11.6689968109131,
17.0608749389648,-29.1000099182129,
20.1492290496826,-33.5568656921387,
19.4454631805420,-4.90514755249023,
31.7720661163330,23.9358634948730,
44.3515930175781,39.2747039794922,
28.9981803894043,43.8292236328125,
-13.6587677001953,32.0242996215820,
-43.8822097778320,-5.18123674392700,
-28.7031059265137,-44.5262756347656,
17.2466278076172,-42.8450126647949,
52.2767944335938,7.03551673889160,
48.9814186096191,56.4810829162598,
21.1511611938477,60.2817230224609,
-0.357814550399780,30.6006031036377,
-8.51388072967529,11.8124132156372,
-16.4598140716553,11.4235849380493,
-33.5045623779297,8.27646446228027,
-49.2684936523438,0.870152175426483,
-47.5377922058106,12.6476850509644,
-26.7726001739502,40.6592216491699,
-12.7137918472290,45.4790916442871,
-19.5743083953857,5.62829732894898,
-26.7025356292725,-44.7598114013672,
1.28153920173645,-53.1267280578613,
52.5357818603516,-18.6114349365234,
72.7571411132813,18.8528175354004,
35.0067710876465,35.9842834472656,
-21.3068275451660,44.5885620117188,
-32.0818138122559,53.5362243652344,
2.81767034530640,41.1573791503906,
21.1946716308594,-3.17095851898193,
-6.52483463287354,-48.1320152282715,
-35.6046218872070,-59.5595436096191,
-13.2686014175415,-36.4266395568848,
41.8142967224121,-8.54023170471191,
65.8191909790039,6.63571834564209,
41.2156372070313,15.6565113067627,
15.1441698074341,22.5741386413574,
19.4122428894043,18.7904415130615,
31.1982192993164,1.26402914524078,
10.6221532821655,-13.3650817871094,
-32.2415161132813,-14.2316484451294,
-53.6716651916504,-13.5817003250122,
-35.8637390136719,-21.1754550933838,
-1.83002901077271,-26.4010391235352,
17.8341751098633,-14.3212366104126,
16.9218463897705,4.44061613082886,
8.23058414459229,2.60037231445313,
0.682892799377441,-21.6792030334473,
3.96108150482178,-39.4746818542481,
22.7107715606689,-28.3322315216064,
42.6223258972168,-1.09745657444000,
33.0051422119141,7.25844621658325,
-8.21548271179199,-6.64347457885742,
-52.1960792541504,-15.7913541793823,
-61.3798294067383,0.790139555931091,
-32.2042884826660,24.7875995635986,
0.822767734527588,27.4770584106445,
4.25540494918823,3.99792242050171,
-19.1797447204590,-21.5238323211670,
-37.7570266723633,-19.0247230529785,
-30.3649616241455,11.7272291183472,
2.41032171249390,39.9740486145020,
36.2946395874023,39.3998527526856,
42.3359451293945,18.6921157836914,
21.5208797454834,7.09462833404541,
3.90167164802551,20.7407989501953,
18.3352127075195,39.9277648925781,
49.8975830078125,36.7590141296387,
54.6245727539063,15.8563776016235,
16.0269279479980,15.2666883468628,
-26.9083347320557,43.1671295166016,
-29.8872089385986,53.7164192199707,
-5.40547084808350,12.9153156280518,
-6.85049486160278,-42.6276969909668,
-41.3949012756348,-46.6530227661133,
-56.2827835083008,7.71305465698242,
-16.8471336364746,51.5978126525879,
32.0032768249512,30.6062297821045,
23.9297237396240,-19.3184051513672,
-35.9682350158691,-31.6516799926758,
-76.2118072509766,-4.88180780410767,
-55.1152458190918,12.9929256439209,
-15.3248643875122,4.34055709838867,
-10.8717813491821,4.30729675292969,
-35.2093963623047,25.5368614196777,
-39.0611572265625,28.8276977539063,
-10.0863838195801,-7.95057678222656,
15.9619350433350,-40.6234741210938,
10.2060661315918,-18.5646286010742,
-8.68390274047852,29.9708881378174,
-16.5813236236572,33.2270812988281,
-13.3062763214111,-20.2712707519531,
-9.05653381347656,-64.4937667846680,
2.44921016693115,-42.6080780029297,
30.9691333770752,12.7538585662842,
63.6568183898926,35.9692916870117,
71.4982070922852,15.9563446044922,
42.2830734252930,-9.65772342681885,
0.203851699829102,-16.7895603179932,
-24.1392822265625,-12.5351324081421,
-25.2309494018555,-5.20587396621704,
-13.7861146926880,9.47818565368652,
-3.89154505729675,31.5491981506348,
-7.42744731903076,42.8331336975098,
-26.1060733795166,32.8758811950684,
-42.4720268249512,5.39470720291138,
-35.8924026489258,-22.6108188629150,
-5.74093437194824,-45.0747528076172,
24.3416786193848,-59.1891555786133,
32.3323783874512,-52.5763778686523,
27.4224033355713,-27.6534957885742,
34.6139373779297,-10.0994863510132,
54.1877937316895,-13.9949207305908,
61.6797714233398,-23.2665729522705,
41.3072776794434,-20.9545974731445,
10.1942911148071,-12.2792387008667,
-11.3182353973389,-10.5084733963013,
-21.3834514617920,-16.4738388061523,
-28.3717918395996,-18.9331512451172,
-28.3703498840332,-23.7885990142822,
-12.9038562774658,-49.1760978698731,
6.87739181518555,-76.2880020141602,
8.41059017181397,-60.6889877319336,
-11.6402101516724,0.950942039489746,
-24.0497817993164,46.6802330017090,
-5.73750257492065,30.4769802093506,
26.2531147003174,-5.58109235763550,
36.3660774230957,6.75686120986939,
16.3455314636230,50.8292884826660,
-14.8407859802246,48.6504249572754,
-34.4464187622070,-21.3948192596436,
-40.0786743164063,-79.6797485351563,
-34.0457382202148,-56.2041664123535,
-22.1352138519287,8.63295173645020,
-12.4754524230957,20.0874080657959,
-15.3617792129517,-31.0428619384766,
-25.1871089935303,-70.2620697021484,
-15.7425403594971,-51.2880592346191,
21.1480026245117,-8.03004550933838,
54.7042350769043,16.0493431091309,
48.6760139465332,29.0575771331787,
9.98929405212402,50.0875740051270,
-15.5980157852173,56.1838531494141,
-3.13477373123169,22.3773231506348,
24.2767295837402,-24.5015563964844,
30.1537780761719,-31.0881633758545,
13.4974298477173,2.37747788429260,
1.82535517215729,24.4116859436035,
5.41586303710938,7.72596359252930,
7.30746507644653,-9.67759704589844,
0.314741551876068,14.1632671356201,
-1.14195013046265,52.7957344055176,
14.4853763580322,52.8807678222656,
28.2545661926270,9.47175121307373,
14.1290826797485,-31.7234611511230,
-20.2901573181152,-34.4472465515137,
-37.1855278015137,-6.31771278381348,
-21.2587833404541,15.0080528259277,
-0.568964004516602,11.2358980178833,
-6.09318351745606,-0.0109558701515198,
-29.1822738647461,3.80085730552673,
-35.9538726806641,20.0785198211670,
-14.5688982009888,26.3750667572022,
7.16525983810425,6.87235307693481,
7.99842691421509,-24.7372608184814,
-3.86662697792053,-33.3044700622559,
-9.29728698730469,-8.16072750091553,
-10.3263053894043,18.9387264251709,
-21.1484088897705,13.4441280364990,
-34.1713256835938,-13.9797782897949,
-29.0247097015381,-20.7424678802490,
-3.77481365203857,5.21898221969605,
13.0746698379517,28.1178188323975,
5.06056308746338,9.08468151092529,
-7.33499288558960,-38.7203140258789,
3.21195507049561,-63.8217506408691,
32.1703376770020,-41.0182647705078,
50.2069396972656,1.86903643608093,
45.2685356140137,19.7357463836670,
31.7083911895752,1.58497405052185,
23.1730098724365,-23.9497814178467,
10.6080055236816,-28.7062053680420,
-12.3864631652832,-14.4012851715088,
-33.0266418457031,-2.12315011024475,
-28.5995635986328,-3.51499509811401,
3.39489054679871,-9.73015213012695,
39.1184120178223,-5.53763294219971,
56.3342514038086,7.57386112213135,
54.8107032775879,11.1715803146362,
41.9180603027344,-2.30727934837341,
19.3355083465576,-20.2054500579834,
-13.3762731552124,-20.6939582824707,
-40.6727142333984,0.136398553848267,
-39.5006828308106,18.7014598846436,
-8.88876724243164,10.8425350189209,
16.2661685943604,-20.6822185516357,
-1.36070954799652,-40.4837036132813,
-47.6645278930664,-22.4942073822022,
-66.2987136840820,15.5820074081421,
-30.6919002532959,30.9698638916016,
22.1936416625977,8.43822765350342,
37.2488517761231,-18.6785812377930,
10.1378421783447,-11.1055040359497,
-15.9705381393433,17.4067478179932,
-18.0660152435303,16.3896312713623,
-13.1639041900635,-22.7487964630127,
-14.8178148269653,-53.0193862915039,
-6.70285320281982,-32.8059043884277,
23.0220870971680,17.2235717773438,
38.8393478393555,44.0289764404297,
4.60118198394775,29.8230037689209,
-54.0614395141602,4.52084779739380,
-75.2254486083984,-10.0565176010132,
-39.0457305908203,-16.7966194152832,
10.8814630508423,-16.7443695068359,
28.3479003906250,7.22274017333984,
19.5051784515381,48.9430770874023,
5.00408935546875,62.6075210571289,
-5.71302461624146,15.5931377410889,
-12.8119916915894,-54.6766738891602,
-4.33045101165772,-81.4394149780273,
28.5946884155273,-48.2158393859863,
56.8834114074707,-3.51387858390808,
42.2638130187988,8.29998397827148,
-0.194899082183838,-1.64615511894226,
-20.3825454711914,-2.53165292739868,
0.720487117767334,11.9867897033691,
24.9318027496338,23.7766132354736,
16.0085372924805,31.1822948455811,
-10.2770357131958,47.5989952087402,
-30.3818740844727,64.7527618408203,
-42.1562957763672,57.0919876098633,
-60.4311218261719,22.2956008911133,
-71.8863449096680,-2.38367390632629,
-43.8987770080566,10.1713752746582,
9.98494911193848,37.6132049560547,
36.9202690124512,36.9550170898438,
8.11969947814941,-1.04124665260315,
-40.8628082275391,-38.9369850158691,
-55.8112449645996,-36.5433692932129,
-27.9710102081299,-2.66736507415772,
6.42706394195557,24.3829383850098,
21.3573722839355,23.5699310302734,
16.6933956146240,8.57696342468262,
-0.467560291290283,2.31462860107422,
-30.8716144561768,9.48755073547363,
-63.2085227966309,14.6389122009277,
-68.0310287475586,2.89171218872070,
-26.9786586761475,-17.1627712249756,
37.2743682861328,-26.6053256988525,
74.2730331420898,-23.9894962310791,
59.6604347229004,-19.8162269592285,
21.3235263824463,-20.0072746276855,
-0.341583997011185,-12.6782999038696,
5.59521818161011,7.06045913696289,
17.0827503204346,22.4575786590576,
15.3287973403931,8.83827686309815,
6.36318016052246,-29.1952629089355,
7.61097431182861,-47.7204704284668,
10.6692972183228,-20.6888294219971,
-1.75667953491211,23.2173309326172,
-27.5367527008057,33.7147521972656,
-35.8861007690430,-1.70886468887329,
-6.22434520721436,-40.0622367858887,
43.3075561523438,-38.1707763671875,
70.5543746948242,-1.88248431682587,
57.4951667785645,29.5929012298584,
23.9743576049805,36.7732887268066,
0.936432123184204,31.0248394012451,
-8.73698329925537,26.2553501129150,
-17.7730636596680,15.6160984039307,
-30.6870517730713,-12.5980262756348,
-33.1183547973633,-45.7204933166504,
-14.2048091888428,-58.9323883056641,
17.6035594940186,-46.8651275634766,
41.0336112976074,-27.7699871063232,
45.0511093139648,-19.8391819000244,
38.6543655395508,-21.8561496734619,
36.5298080444336,-23.1306228637695,
37.8446197509766,-15.3711147308350,
35.5267791748047,-0.756095767021179,
30.9804000854492,6.09465312957764,
28.5828304290772,-1.31780362129211,
26.2720222473145,-14.0263319015503,
13.6808109283447,-12.6180715560913,
-6.69387340545654,18.3257408142090,
-14.1529216766357,55.3836555480957,
2.98021316528320,54.7731132507324,
24.0104675292969,10.8833732604980,
14.9336986541748,-28.7788963317871,
-18.3526515960693,-26.8414268493652,
-36.1975975036621,-4.81128978729248,
-21.2003803253174,-1.55304884910584,
-3.42488193511963,-15.5240478515625,
-15.3129940032959,-13.2794456481934,
-38.5271644592285,5.08455562591553,
-33.6771011352539,-5.38340568542481,
-0.489101052284241,-51.4069824218750,
22.9998931884766,-68.2634277343750,
15.6912527084351,-13.5039463043213,
1.40662384033203,52.4211387634277,
4.93513441085815,42.2515411376953,
7.76132726669312,-27.7293491363525,
-13.4882946014404,-61.1226692199707,
-39.5823898315430,-20.0368423461914,
-32.4265441894531,27.0204582214355,
6.66334438323975,20.8932437896729,
36.3063659667969,-6.62485361099243,
29.5235900878906,2.37317347526550,
3.85711693763733,25.4518833160400,
-13.2782468795776,0.373789310455322,
-12.8510599136353,-60.7183799743652,
2.94955110549927,-81.8178100585938,
36.4888687133789,-40.0759811401367,
74.9373626708984,-0.331415057182312,
81.7608413696289,-8.35769367218018,
34.8056564331055,-20.8443355560303,
-29.4382972717285,10.1097965240479,
-49.0498352050781,49.5581207275391,
-11.2937278747559,35.5769691467285,
26.0631885528564,-17.6740245819092,
16.0191383361816,-35.4609146118164,
-22.3442344665527,13.7015991210938,
-42.6187362670898,70.1578216552734,
-26.8719444274902,66.8966751098633,
-2.45454597473145,17.1795139312744,
4.35412597656250,-20.4367885589600,
4.29413747787476,-21.6914234161377,
16.8016242980957,-5.75269508361816,
36.8322448730469,7.16726398468018,
39.8521881103516,6.10276556015015,
17.9889163970947,-13.4475126266480,
-11.8868322372437,-41.9661064147949,
-14.9222660064697,-54.1786651611328,
23.1184883117676,-34.9552688598633,
74.5379486083984,-0.979023456573486,
84.0158386230469,14.5583515167236,
27.6215934753418,6.42939472198486,
-46.6887321472168,6.58112430572510,
-70.0394973754883,23.5911407470703,
-29.9419345855713,26.0064868927002,
17.7056617736816,-5.60196304321289,
21.3633785247803,-32.4570426940918,
0.0783522054553032,-8.30051422119141,
-2.40043401718140,54.6115798950195,
12.0597124099731,91.6534881591797,
-2.18119192123413,67.8390426635742,
-51.2517318725586,15.4046840667725,
-80.0755538940430,-19.3606853485107,
-49.0468673706055,-33.6539421081543,
14.5340709686279,-47.9421691894531,
50.3780021667481,-54.2175559997559,
42.0435142517090,-24.2122859954834,
21.4578094482422,38.5040168762207,
12.6045417785645,84.3278579711914,
7.33789587020874,75.0753479003906,
-1.09607875347137,28.7996177673340,
-8.03245639801025,-9.37629699707031,
-12.9117794036865,-17.2579059600830,
-30.9307842254639,-1.39003467559814,
-59.6985130310059,17.0663757324219,
-68.4516296386719,24.8224258422852,
-39.3161582946777,21.7871398925781,
-7.77069282531738,14.6922788619995,
-18.0397739410400,10.9448041915894,
-61.2306709289551,14.5875120162964,
-82.6668777465820,14.0899400711060,
-53.4285774230957,-0.499007225036621,
-5.12691307067871,-16.4803161621094,
15.9568128585815,-19.4727210998535,
8.32653999328613,-15.3318099975586,
6.10245418548584,-19.6939811706543,
23.2823925018311,-24.5681190490723,
37.7540626525879,-4.21299457550049,
26.9779663085938,40.0429115295410,
-2.61555814743042,64.0970153808594,
-32.1531715393066,35.3228950500488,
-51.5944824218750,-17.8750076293945,
-55.6680374145508,-41.0630760192871,
-41.3594322204590,-27.7992401123047,
-19.9985637664795,-20.6241016387939,
-7.51530122756958,-42.4077186584473,
-18.5706577301025,-57.8563613891602,
-46.9411888122559,-30.5949230194092,
-68.0726928710938,15.1088275909424,
-59.3143005371094,23.7833709716797,
-23.1411247253418,-13.0608186721802,
22.1170902252197,-47.7011032104492,
45.9042816162109,-38.8852272033691,
25.6637153625488,-2.89619421958923,
-17.9894351959229,18.0920810699463,
-30.8244209289551,11.0490074157715,
10.9883308410645,-1.57508301734924,
61.3130073547363,-1.76896357536316,
53.4060821533203,5.72668695449829,
-12.3675136566162,9.52068138122559,
-56.6134529113770,4.77617597579956,
-26.2830848693848,-9.81748771667481,
36.2960624694824,-23.9556007385254,
50.4729270935059,-22.8286399841309,
7.23973941802979,1.71643805503845,
-28.3809623718262,27.3299770355225,
-15.8982362747192,22.5097427368164,
6.13350391387939,-14.8541841506958,
-4.42261028289795,-46.8616905212402,
-32.8647270202637,-41.4529266357422,
-35.1175613403320,-11.4094953536987,
-8.85944175720215,-2.30590605735779,
5.53913021087647,-24.7490329742432,
-9.67795467376709,-46.5169219970703,
-25.2221260070801,-40.2686309814453,
-13.9887075424194,-17.3099956512451,
13.3568792343140,-7.81950712203980,
26.4124660491943,-22.3905429840088,
19.9410610198975,-38.0784416198731,
11.1342906951904,-29.3962707519531,
9.01659393310547,5.22381877899170,
12.3132619857788,40.6524200439453,
20.7455215454102,52.0616378784180,
31.3837337493897,36.0340614318848,
30.7344875335693,19.9882850646973,
9.38299655914307,29.3438529968262,
-18.5927429199219,59.1222267150879,
-21.2133731842041,68.9032287597656,
9.71702289581299,32.3369560241699,
43.9394187927246,-19.8124179840088,
44.3194694519043,-32.6352233886719,
14.8447360992432,1.02681350708008,
-6.16774320602417,38.0057754516602,
2.67432689666748,35.3793106079102,
21.1988773345947,12.7332725524902,
17.2118911743164,15.5423574447632,
-13.1161565780640,49.8046226501465,
-43.9058189392090,71.8490829467773,
-53.2667579650879,48.1537322998047,
-46.4539070129395,-5.03791618347168,
-36.2640953063965,-47.5495567321777,
-23.8911819458008,-58.0278511047363,
-4.13685083389282,-47.6198806762695,
20.1066303253174,-30.8503952026367,
28.7221736907959,-14.9422140121460,
16.2157688140869,-7.04137229919434,
-3.35099148750305,-19.5421905517578,
-10.7795648574829,-48.3251075744629,
-3.53931975364685,-72.5681915283203,
6.50308227539063,-68.7422332763672,
4.94418191909790,-37.4465408325195,
-5.92974185943604,-2.53948783874512,
-17.5905513763428,15.6228218078613,
-31.8868656158447,15.8163728713989,
-48.9588317871094,11.9671916961670,
-54.3259849548340,8.98508644104004,
-30.6071472167969,8.33668041229248,
16.4206504821777,6.61250448226929,
43.3626251220703,7.75674343109131,
18.2765369415283,13.2273674011230,
-42.1639823913574,15.4509248733521,
-74.4594039916992,10.3188304901123,
-49.1029357910156,1.59732210636139,
-8.98282623291016,-3.68165516853333,
-7.38134574890137,-9.27023887634277,
-39.1791000366211,-19.9272117614746,
-47.1647644042969,-30.7049789428711,
-8.28887176513672,-29.2519969940186,
33.1637191772461,-7.61829757690430,
29.5057430267334,21.6393795013428,
-2.46991896629334,40.9212760925293,
-12.4670867919922,42.2257575988770,
0.919122457504273,28.9664573669434,
-7.28969955444336,11.6801595687866,
-43.4213104248047,-5.80341672897339,
-55.3162727355957,-20.5585823059082,
-6.75109291076660,-32.7083435058594,
56.6161499023438,-38.4056243896484,
58.9336280822754,-32.1976318359375,
-0.0754851102828980,-10.0574731826782,
-50.0213699340820,15.8153762817383,
-45.8855476379395,27.1061668395996,
-18.4901905059814,18.0086746215820,
-14.5821485519409,0.0784158706665039,
-24.8881320953369,-15.9776992797852,
-11.0149812698364,-25.2567806243897,
30.1470794677734,-22.4395809173584,
52.9749488830566,0.798259735107422,
35.5126228332520,38.3953704833984,
2.28388428688049,60.2882423400879,
-13.2618513107300,50.6370887756348,
-8.21629810333252,29.7139606475830,
-4.10407733917236,32.8749694824219,
-8.77896785736084,56.5264167785645,
-21.0388202667236,59.9696769714356,
-36.5799446105957,30.1763362884522,
-57.3062095642090,-1.52102077007294,
-70.0710525512695,-5.60595273971558,
-57.0537414550781,0.851958453655243,
-21.1427574157715,-10.5672588348389,
12.7335662841797,-31.2472667694092,
32.7332878112793,-32.5498046875000,
44.0110969543457,-9.82561779022217,
52.6281623840332,9.58710670471191,
46.5989952087402,11.9178962707520,
16.9643573760986,13.5346708297730,
-22.6493301391602,23.8493595123291,
-46.2141532897949,22.0205249786377,
-50.6934280395508,-7.57964611053467,
-49.3573036193848,-42.7541198730469,
-42.8867454528809,-58.8974418640137,
-11.9111509323120,-54.0399322509766,
44.2672996520996,-44.3098793029785,
86.9883422851563,-27.2159938812256,
78.9058609008789,-1.94622492790222,
30.5835151672363,13.0555772781372,
0.0802739262580872,-2.99095153808594,
14.5985193252563,-31.9983024597168,
48.3568496704102,-28.9254112243652,
50.7521247863770,11.5331764221191,
15.3548078536987,39.7929420471191,
-17.2113609313965,13.4274425506592,
-12.9908008575439,-39.1823387145996,
17.3944511413574,-53.4523200988770,
39.7658958435059,-11.3472757339478,
40.6558036804199,43.1499061584473,
28.0234832763672,63.5090751647949,
15.8385477066040,48.1601600646973,
1.97645008563995,21.6434669494629,
-11.7635641098022,3.54080533981323,
-15.2310075759888,-10.1123142242432,
2.76443600654602,-17.7821941375732,
36.4859008789063,-14.9058732986450,
61.7679214477539,0.0136826634407043,
65.5033721923828,16.8178882598877,
47.6084632873535,24.1057071685791,
21.8171195983887,16.5405216217041,
-0.872409701347351,-0.384727716445923,
-17.4651203155518,-19.0581340789795,
-29.1845760345459,-28.5674896240234,
-35.4367828369141,-25.3857765197754,
-36.0841598510742,-18.9269981384277,
-32.9850387573242,-19.4260101318359,
-27.5053634643555,-30.9526023864746,
-23.7651977539063,-48.7272338867188,
-15.0589103698730,-60.5072708129883,
6.33319187164307,-61.2964897155762,
38.4764900207520,-51.5251884460449,
58.9983749389648,-35.8558387756348,
44.6462593078613,-17.8482170104980,
-2.56792855262756,1.65134727954865,
-44.8240547180176,20.5318546295166,
-45.7088737487793,31.5467700958252,
-5.98960971832275,28.2736148834229,
30.5455837249756,10.6778335571289,
30.6870822906494,-6.93146371841431,
2.02624130249023,-12.5984210968018,
-13.4925403594971,-4.69454717636108,
5.66872882843018,5.40976619720459,
36.0284767150879,9.76282501220703,
39.8981742858887,3.25913548469543,
20.8770198822022,-7.86743783950806,
16.2889652252197,-16.0448951721191,
39.6293678283691,-13.7030582427979,
54.4498634338379,-0.633009433746338,
22.6351699829102,14.4016656875610,
-35.3734283447266,16.8121528625488,
-60.7718429565430,5.97810745239258,
-29.0651836395264,-11.5328397750855,
8.95661354064941,-27.4465827941895,
0.224314212799072,-37.4950218200684,
-33.1684951782227,-35.9427299499512,
-37.2830886840820,-19.6498126983643,
-5.80495595932007,-6.84988117218018,
13.1744670867920,-18.7687702178955,
-1.91443920135498,-51.3389244079590,
-14.0349254608154,-66.1343917846680,
10.9315538406372,-34.5972061157227,
43.3835639953613,24.1007804870605,
35.4040718078613,58.6546440124512,
-3.77437758445740,43.6184043884277,
-21.7395229339600,-0.622612953186035,
-11.3078880310059,-35.1010208129883,
-15.3015537261963,-39.8521652221680,
-43.1089591979981,-20.4130764007568,
-45.3423080444336,6.95023202896118,
4.63257503509522,22.5300140380859,
54.0979461669922,10.7426185607910,
45.5990600585938,-17.0070590972900,
7.04439496994019,-35.1612777709961,
7.75023126602173,-30.9390106201172,
47.9335823059082,-19.5881195068359,
55.8207740783691,-16.1926727294922,
4.32724189758301,-20.5003261566162,
-40.3368682861328,-24.2566757202148,
-19.4693031311035,-25.0416107177734,
25.4939270019531,-21.8343372344971,
12.9398937225342,-7.07035970687866,
-48.7920150756836,16.4460849761963,
-76.9007339477539,21.2524662017822,
-32.3042335510254,-9.42142391204834,
27.6331939697266,-43.6616058349609,
35.4205398559570,-35.3238410949707,
-0.0850667953491211,12.6648139953613,
-24.6467952728272,41.3068161010742,
-18.4313163757324,22.6291198730469,
-12.9957656860352,-4.73614549636841,
-26.0275478363037,2.31051731109619,
-34.9598350524902,32.9745368957520,
-22.0311813354492,50.5108680725098,
-0.0656547546386719,42.8628234863281,
13.0241184234619,26.9348278045654,
20.6823329925537,10.2136211395264,
30.8089485168457,-17.2759876251221,
40.1987342834473,-40.0634651184082,
40.3121910095215,-32.9652709960938,
33.7118568420410,-5.46587133407593,
32.5514450073242,0.422599077224731,
35.4166374206543,-20.4942188262939,
28.2888622283936,-18.2932281494141,
16.9093399047852,23.5193080902100,
23.5593070983887,50.7673110961914,
45.6225318908691,22.7512989044189,
49.6561355590820,-19.8516407012939,
20.8991088867188,-11.4014797210693,
-14.3895759582520,34.6924285888672,
-25.6843643188477,41.9973030090332,
-18.3410415649414,-12.1421813964844,
-17.8279247283936,-57.9810523986816,
-25.0580120086670,-49.1461944580078,
-13.4401912689209,-27.5371837615967,
22.2643146514893,-34.7717361450195,
51.0376243591309,-34.9444007873535,
45.2943000793457,18.6193046569824,
18.5987167358398,75.9782180786133,
-5.93029737472534,54.3903923034668,
-19.5436496734619,-29.0059299468994,
-22.5922298431397,-66.4096984863281,
-3.86629676818848,-11.8881244659424,
27.6095027923584,53.6038970947266,
37.0555267333984,45.4157981872559,
2.72869586944580,-0.678912043571472,
-38.7792015075684,1.26965618133545,
-38.7262458801270,45.3838539123535,
0.362493276596069,49.4008140563965,
22.7802066802979,-7.68578577041626,
4.27382373809814,-52.3302803039551,
-18.0347061157227,-42.3255386352539,
-6.48820114135742,-18.3537044525147,
19.8313503265381,-26.1550979614258,
26.8760967254639,-38.9135169982910,
25.5324821472168,-11.1830005645752,
37.9365119934082,34.6159744262695,
46.2230491638184,43.1297645568848,
17.9939613342285,10.9231433868408,
-32.7956619262695,-2.24817800521851,
-54.8977737426758,29.8475284576416,
-31.8183498382568,57.2608985900879,
-8.30291461944580,39.6603813171387,
-19.9799919128418,4.11000299453735,
-45.8344993591309,-11.7213125228882,
-49.4750213623047,-9.71574974060059,
-35.1207313537598,-14.0674343109131,
-29.1360321044922,-19.7499294281006,
-22.8796234130859,-7.66944932937622,
0.00900799036026001,19.4557437896729,
20.3776149749756,35.7561683654785,
2.61468362808228,36.5118484497070,
-37.9453468322754,37.3179588317871,
-47.8151359558106,40.2139968872070,
-8.63885402679443,22.4734859466553,
25.9952259063721,-14.0733795166016,
7.40857267379761,-29.2265205383301,
-38.5223426818848,-6.92275428771973,
-49.1031188964844,14.5395488739014,
-14.1040840148926,-2.58178019523621,
15.0788106918335,-40.9511260986328,
9.91787052154541,-53.4929656982422,
-1.64326572418213,-28.6397209167480,
13.6524801254272,2.21402740478516,
41.6839828491211,11.2841148376465,
47.6770935058594,7.43741607666016,
33.7641754150391,1.70238614082336,
28.9532947540283,-11.6472768783569,
39.6253051757813,-30.4720249176025,
38.0004081726074,-32.5562477111816,
7.29778575897217,-7.95675516128540,
-28.0387496948242,15.0187788009644,
-28.6531105041504,2.54131174087524,
3.77932119369507,-31.2042865753174,
29.1556930541992,-40.5663833618164,
25.6147975921631,-10.8141059875488,
12.8657207489014,26.9642925262451,
13.1566896438599,40.3646087646484,
21.1090354919434,34.2994613647461,
7.27652502059937,35.5507659912109,
-35.1487083435059,50.2042007446289,
-68.3419876098633,52.0908508300781,
-57.7006340026856,25.0004959106445,
-17.3782730102539,-17.5563068389893,
8.36391544342041,-48.5528526306152,
-5.72332763671875,-48.3904762268066,
-28.5041007995605,-25.5822219848633,
-18.7475872039795,-5.83908319473267,
22.0059013366699,-7.81675243377686,
46.8796844482422,-20.4021129608154,
20.5397663116455,-12.6177139282227,
-28.5129566192627,22.8896064758301,
-43.8812370300293,51.7632026672363,
-8.71946144104004,42.0801849365234,
32.5187988281250,1.64377975463867,
27.4497318267822,-22.7983646392822,
-20.5619106292725,-2.05095243453980,
-55.3675460815430,28.8903903961182,
-33.9014205932617,22.0171680450439,
23.7710571289063,-21.3878459930420,
64.8848266601563,-53.3516693115234,
64.6293258666992,-48.3526344299316,
35.8363113403320,-18.0917739868164,
2.30657482147217,10.0069379806519,
-24.1839103698730,30.3555889129639,
-38.3449249267578,36.8696556091309,
-37.6437911987305,10.8789787292480,
-27.2222061157227,-46.5601806640625,
-23.8804759979248,-81.4677734375000,
-23.6949481964111,-45.5530014038086,
-7.58480739593506,27.5919132232666,
25.5720634460449,52.9048995971680,
47.3012084960938,5.63218688964844,
28.0949611663818,-39.0980682373047,
-12.4137239456177,-18.8527202606201,
-29.6116142272949,24.3737354278564,
-12.2462806701660,10.4341573715210,
3.17780923843384,-55.8353576660156,
-5.64166021347046,-86.9907531738281,
-16.8870754241943,-42.6128120422363,
-3.32847094535828,11.6271200180054,
30.2558097839355,5.67506837844849,
55.2834548950195,-35.7599105834961,
61.2514419555664,-43.8544692993164,
54.0117721557617,-7.06994915008545,
34.0673217773438,19.1198558807373,
-3.51620149612427,2.33993482589722,
-35.6723213195801,-24.1483440399170,
-28.1531047821045,-30.1849498748779,
16.5788917541504,-25.0644893646240,
55.5943145751953,-24.4876194000244,
56.5833587646484,-19.9605140686035,
36.1974716186523,5.38452053070068,
21.3296127319336,38.5119285583496,
5.33986330032349,41.9238014221191,
-28.4334487915039,11.8898248672485,
-65.2891159057617,-14.5097169876099,
-65.5817337036133,-11.5470228195190,
-23.2975788116455,13.7401905059814,
14.1809368133545,34.1115646362305,
6.27976560592651,29.3988018035889,
-24.7174549102783,-3.17637395858765,
-29.1372661590576,-34.9802436828613,
4.85632896423340,-32.1530952453613,
36.5976219177246,8.30616950988770,
30.6962318420410,48.3470382690430,
-1.29012560844421,46.8782958984375,
-25.6152381896973,13.3120737075806,
-21.9911651611328,2.32490563392639,
0.756912112236023,36.7683372497559,
22.3563613891602,69.4166030883789,
31.2484779357910,49.1120681762695,
23.6053199768066,-4.72807455062866,
4.23949527740479,-30.6287803649902,
-12.0644149780273,-15.7815656661987,
-15.8568134307861,-9.47955894470215,
-11.9229192733765,-39.0341758728027,
-12.0602884292603,-63.8535041809082,
-15.6155376434326,-35.5348968505859,
-15.8084697723389,19.5803546905518,
-15.9594001770020,37.6136703491211,
-23.3477191925049,7.53950691223145,
-34.1350326538086,-16.5003395080566,
-35.8064308166504,3.17668938636780,
-20.5189971923828,33.3598136901856,
-0.803450822830200,18.9075565338135,
8.89043235778809,-26.3523502349854,
13.3645668029785,-47.6402740478516,
24.1938705444336,-18.3627204895020,
35.6517906188965,26.8916549682617,
38.3164100646973,45.2765083312988,
34.7574348449707,28.3113746643066,
35.1427955627441,5.87856817245483,
32.9974403381348,6.85438203811646,
14.0941419601440,28.1558609008789,
-14.1673851013184,44.7163276672363,
-16.8204288482666,34.4525299072266,
16.7683849334717,2.39194512367249,
47.8014984130859,-13.1890106201172,
31.7138080596924,15.7402362823486,
-20.5098495483398,58.0690727233887,
-55.5003890991211,51.5480041503906,
-44.3934669494629,-11.7385540008545,
-21.4217166900635,-67.2092056274414,
-26.2221221923828,-60.8800086975098,
-47.7892341613770,-15.4245929718018,
-46.2643966674805,2.34760975837708,
-12.3025255203247,-18.8082523345947,
21.2182750701904,-23.2376537322998,
20.7357940673828,21.4487571716309,
-11.6561002731323,65.8312225341797,
-40.3483238220215,55.1382484436035,
-38.0522308349609,7.87336492538452,
-8.11812686920166,-17.5132274627686,
20.6280879974365,-5.97164201736450,
21.0333175659180,-2.16391515731812,
-6.36519861221314,-26.2860260009766,
-33.3259811401367,-40.4880180358887,
-32.4949760437012,-12.9682779312134,
-14.2530918121338,21.2756366729736,
-11.9692420959473,11.1999263763428,
-25.1193103790283,-36.7656593322754,
-19.5555458068848,-66.2906494140625,
16.0773410797119,-47.8591003417969,
45.6812286376953,-19.7893009185791,
29.9454879760742,-23.4399223327637,
-15.8887338638306,-41.5716476440430,
-39.3690910339356,-30.2011528015137,
-22.0281314849854,10.5775156021118,
0.171730697154999,43.1401138305664,
1.67774605751038,38.7011184692383,
-3.18709778785706,13.2699785232544,
1.99474108219147,3.28049397468567,
3.83228921890259,13.4981632232666,
-12.8890905380249,21.1925735473633,
-24.5526084899902,14.8217592239380,
-2.52121424674988,9.91743469238281,
31.0193023681641,22.6567592620850,
22.6784057617188,42.0302429199219,
-36.2289695739746,41.2344474792481,
-84.3629074096680,6.84132099151611,
-72.1777267456055,-36.5098228454590,
-22.7682285308838,-43.6399688720703,
1.00065732002258,-2.87356472015381,
-16.4814014434814,44.8073997497559,
-31.3031749725342,45.7414855957031,
-10.7271757125855,-2.54912137985230,
21.6377105712891,-51.0961189270020,
28.9944076538086,-51.7382087707520,
12.6249284744263,-13.3147258758545,
7.97836875915527,20.6599121093750,
26.6075096130371,28.0970516204834,
37.8596992492676,28.6272811889648,
14.8450946807861,37.8138198852539,
-31.6519813537598,44.2250251770020,
-62.1155090332031,31.8612117767334,
-55.4229049682617,7.92435550689697,
-26.0061893463135,-10.4499406814575,
4.25854110717773,-19.1175594329834,
29.1190338134766,-25.8091220855713,
39.6983222961426,-25.5653438568115,
31.7232456207275,-6.35662078857422,
8.47556972503662,19.5322704315186,
-5.83640861511231,23.4614601135254,
8.70903587341309,3.32774400711060,
38.8065147399902,-10.0662279129028,
41.0541534423828,8.84999561309815,
-1.63939499855042,40.2404479980469,
-53.3803749084473,42.0013122558594,
-65.9564971923828,9.97815322875977,
-31.0300064086914,-22.0568542480469,
10.6476888656616,-27.7104396820068,
20.8472328186035,-17.0272312164307,
4.88471412658691,-9.66404819488525,
2.35275745391846,-10.0592088699341,
26.6199226379395,-6.05564546585083,
53.5464057922363,6.91215276718140,
51.6064529418945,13.4735822677612,
23.2322349548340,2.67334032058716,
3.42845344543457,-18.9499416351318,
15.1624460220337,-29.7738418579102,
38.7188415527344,-13.2580585479736,
34.0866546630859,29.9699726104736,
-9.34260177612305,68.8821640014648,
-54.2449836730957,62.6528358459473,
-66.5008010864258,11.8629341125488,
-52.0419082641602,-30.5315723419189,
-40.0208511352539,-23.1816768646240,
-46.1802062988281,12.7075862884521,
-47.3929748535156,16.9621162414551,
-29.1733169555664,-30.2747097015381,
-8.87097454071045,-73.9661941528320,
-9.64412117004395,-62.8970031738281,
-23.1151924133301,-19.4706954956055,
-18.1965293884277,-0.400780916213989,
8.22122955322266,-10.0148696899414,
28.5758266448975,0.177302837371826,
24.6465110778809,38.2292518615723,
15.4349613189697,52.5871810913086,
23.6652545928955,15.5810832977295,
38.0127601623535,-27.4340877532959,
27.4127750396729,-15.9885063171387,
-12.1452093124390,30.5531806945801,
-51.6704597473145,40.8950271606445,
-66.1322250366211,-5.58483314514160,
-58.7218437194824,-49.2013702392578,
-37.0494613647461,-40.9619178771973,
-3.51059556007385,-0.878544092178345,
34.8318824768066,22.6529598236084,
52.8038711547852,19.5877342224121,
34.6568679809570,7.18280506134033,
2.73241949081421,-14.4883289337158,
-4.08858823776245,-45.6624221801758,
16.5243377685547,-58.4541358947754,
28.5418682098389,-22.6954803466797,
8.67517089843750,36.3177947998047,
-22.2754192352295,51.2659721374512,
-22.4116554260254,3.13057065010071,
15.8044099807739,-46.2284545898438,
49.7685699462891,-30.0382347106934,
40.7160835266113,36.6081962585449,
0.813079357147217,77.9158096313477,
-22.1618061065674,58.3882713317871,
2.08929157257080,18.4336433410645,
43.0976867675781,10.0401086807251,
48.0924034118652,33.2168960571289,
1.57447171211243,51.1390075683594,
-53.6038208007813,44.4834175109863,
-67.4318618774414,31.3487510681152,
-45.3563957214356,26.8669052124023,
-28.0369987487793,19.0475940704346,
-31.2943191528320,-3.99284601211548,
-29.9468250274658,-26.1251678466797,
-5.09656429290772,-18.6926631927490,
24.1923103332520,15.2122764587402,
25.5340785980225,37.3453445434570,
4.85120820999146,23.7090816497803,
-4.98792123794556,-11.0374984741211,
2.49147105216980,-24.2471446990967,
3.66666913032532,2.30733466148376,
-11.8138628005981,41.8241386413574,
-21.3569011688232,56.9580764770508,
-8.75457859039307,39.0775070190430,
3.22746562957764,9.60446071624756,
-15.4061203002930,-3.72430396080017,
-45.9521026611328,4.51716566085815,
-47.2981567382813,15.0336856842041,
-14.3616161346436,8.95787429809570,
13.1325273513794,-11.0069103240967,
2.48143291473389,-24.1266403198242,
-27.1025257110596,-24.1255741119385,
-39.6072311401367,-21.4520454406738,
-29.3394565582275,-22.2113018035889,
-16.1734104156494,-23.7286586761475,
-9.61049747467041,-19.9358081817627,
-1.93582856655121,-20.1571617126465,
2.82258319854736,-36.1809349060059,
-3.85846424102783,-55.7635803222656,
-9.69270610809326,-60.6522750854492,
8.76811981201172,-52.3727226257324,
46.9972839355469,-47.3630828857422,
66.1161651611328,-44.7647819519043,
41.6902694702148,-23.8963775634766,
-1.58751428127289,9.84375095367432,
-20.3663768768311,16.6174945831299,
-6.96145629882813,-16.9081821441650,
3.98671054840088,-46.8156509399414,
-3.50319457054138,-23.2884330749512,
-16.4381942749023,33.4673080444336,
-23.8485469818115,58.7037582397461,
-33.5362586975098,26.8839759826660,
-43.4903221130371,-17.8743190765381,
-35.3266296386719,-32.8704032897949,
-4.20184850692749,-33.8785591125488,
23.5328884124756,-46.1605987548828,
22.7104358673096,-53.7314910888672,
10.3569192886353,-28.2066116333008,
16.4703044891357,4.76168537139893,
35.1261520385742,1.76647818088532,
31.8993053436279,-36.9088859558106,
1.37783908843994,-54.5254859924316,
-9.78088760375977,-25.0168304443359,
20.2476863861084,16.6660594940186,
55.7694778442383,29.1797351837158,
52.5340347290039,22.4212303161621,
18.8250446319580,24.3588180541992,
-1.12553215026855,26.4064178466797,
4.40468311309814,0.587287187576294,
7.45201349258423,-39.5432510375977,
-9.42906284332275,-45.6017913818359,
-29.2520370483398,-11.9832172393799,
-33.5763015747070,11.9723901748657,
-31.3493938446045,-9.02562046051025,
-33.1895332336426,-51.7395439147949,
-20.7878055572510,-72.8252563476563,
20.0497322082520,-58.5727539062500,
62.0017471313477,-31.9224624633789,
62.2909507751465,-5.42817974090576,
21.7897834777832,21.7308959960938,
-15.4008235931396,41.6893730163574,
-18.1999797821045,34.7161750793457,
5.00448513031006,6.70681810379028,
25.2956333160400,-12.3297128677368,
25.9264221191406,-11.9764699935913,
12.8422307968140,-6.63434123992920,
-3.25211787223816,-5.00504446029663,
-10.5968189239502,11.3553771972656,
-2.21621656417847,49.0582771301270,
14.6828565597534,69.9015045166016,
15.5095281600952,35.7376289367676,
-3.76112413406372,-35.7162628173828,
-18.0436401367188,-78.4298171997070,
-11.3563385009766,-59.5140647888184,
-9.82480430603027,-18.6183929443359,
-35.1702537536621,-2.33653783798218,
-65.2769088745117,-7.46876811981201,
-63.5531768798828,0.559966802597046,
-30.7035999298096,23.2377662658691,
-5.81401109695435,24.3308963775635,
-7.36219215393066,-8.31547164916992,
-7.75847959518433,-39.7138137817383,
10.4179162979126,-33.0442352294922,
12.1629333496094,1.02653527259827,
-23.7454147338867,24.5219554901123,
-54.8564224243164,23.6443405151367,
-29.8763980865479,20.9215660095215,
23.9755401611328,30.3326797485352,
26.9028949737549,37.6657333374023,
-35.7280082702637,26.2090969085693,
-86.0289382934570,6.86896324157715,
-59.9709930419922,-4.69512939453125,
-1.52161347866058,-1.70119321346283,
5.24259662628174,6.32960605621338,
-40.4362907409668,12.5854616165161,
-66.9017028808594,16.4658241271973,
-38.4785156250000,19.2087497711182,
-7.93557262420654,19.2761878967285,
-27.2773189544678,13.0768280029297,
-64.8210220336914,-0.551153004169464,
-57.8047714233398,-20.2305259704590,
-6.56045007705689,-43.1019439697266,
28.1117286682129,-58.0735092163086,
13.9985485076904,-59.5333557128906,
-9.11822319030762,-55.9192886352539,
4.64355611801148,-53.4530296325684,
46.6031532287598,-42.2322082519531,
61.6903800964356,-20.8760147094727,
26.6903038024902,-5.93698692321777,
-16.2583961486816,-10.8063926696777,
-24.3888969421387,-20.6720695495605,
7.21967697143555,-12.8663721084595,
43.9873542785645,5.30890941619873,
50.0037612915039,5.65740489959717,
19.8784980773926,-12.5595741271973,
-17.8627872467041,-12.9297838211060,
-32.7479591369629,20.6730308532715,
-18.4597682952881,42.3980751037598,
6.08104562759399,14.5738945007324,
20.7664375305176,-29.6042156219482,
24.9071121215820,-23.9994049072266,
32.7238807678223,28.0493354797363,
40.4839439392090,54.3282356262207,
21.5089378356934,19.5352687835693,
-30.4833393096924,-20.5955638885498,
-72.5775527954102,-11.9697427749634,
-61.3741531372070,21.0054168701172,
-5.66429758071899,13.2255392074585,
37.6362838745117,-32.5586318969727,
30.2546081542969,-48.3312149047852,
-6.07437849044800,-4.05786132812500,
-28.1710529327393,40.9099693298340,
-30.5401020050049,27.7140045166016,
-33.0751266479492,-26.7412319183350,
-41.4902763366699,-62.5927467346191,
-38.3997879028320,-58.9656333923340,
-17.4254379272461,-41.9945297241211,
0.297145187854767,-31.5020637512207,
1.81721127033234,-25.4355468750000,
0.553377091884613,-27.3935737609863,
9.46328639984131,-42.2143936157227,
19.6250991821289,-59.9333076477051,
14.6445865631104,-51.1731109619141,
1.69505167007446,-14.9208860397339,
-4.12532377243042,4.05599164962769,
2.30449819564819,-25.3045749664307,
8.43254852294922,-70.2342147827148,
8.62231159210205,-74.7656326293945,
12.8951826095581,-35.7597427368164,
20.3140392303467,4.51287698745728,
18.4342079162598,16.6141262054443,
7.66068983078003,6.99853849411011,
6.33040952682495,0.843547165393829,
18.7795047760010,5.18975830078125,
22.8561477661133,15.5628986358643,
1.48662090301514,31.7810325622559,
-31.3597049713135,44.0749740600586,
-46.2155532836914,36.1337585449219,
-36.4781150817871,6.66940116882324,
-24.2817726135254,-15.9575309753418,
-20.8989734649658,-7.95726442337036,
-13.2305803298950,5.21509075164795,
5.46431207656860,-7.29009628295898,
21.7532138824463,-28.3350257873535,
23.0087108612061,-15.0969295501709,
16.9519672393799,38.4764785766602,
14.6115932464600,84.9383239746094,
4.37704753875732,76.7572555541992,
-26.5749320983887,27.1012496948242,
-58.5065498352051,-18.4855270385742,
-55.4902076721191,-36.1116561889648,
-16.4429950714111,-31.2244663238525,
16.4150524139404,-8.38300228118897,
4.77911472320557,23.0151252746582,
-35.7943954467773,33.5786285400391,
-52.2558517456055,-1.28641772270203,
-24.2210941314697,-52.0582351684570,
20.4723243713379,-55.7537345886231,
39.1520652770996,8.16790962219238,
18.9511871337891,78.8579864501953,
-20.2687683105469,86.3468399047852,
-45.9133033752441,35.4952697753906,
-41.3457450866699,-13.2616748809814,
-17.8970012664795,-27.2167606353760,
0.00783510506153107,-31.6321468353272,
1.05725264549255,-54.0755577087402,
3.56214308738709,-69.3729934692383,
26.8656654357910,-43.0574684143066,
56.3877143859863,9.34035015106201,
54.2340812683106,41.5310783386231,
7.44357776641846,33.4432678222656,
-44.2269706726074,15.8711719512939,
-51.0344848632813,24.2237033843994,
-17.8292865753174,46.9883155822754,
9.22510147094727,50.4008789062500,
1.13802123069763,21.0914039611816,
-22.7876873016357,-11.3134031295776,
-29.6786098480225,-15.7171020507813,
-14.4805660247803,3.65531134605408,
3.39388132095337,16.6608772277832,
15.3052158355713,2.57670998573303,
25.6675243377686,-26.9695510864258,
35.3724327087402,-37.7403602600098,
32.3818511962891,-11.4785919189453,
15.1460599899292,34.3883972167969,
-5.61295604705811,57.4676551818848,
-17.4187602996826,36.2373428344727,
-22.8333911895752,-13.1035270690918,
-32.6985473632813,-53.0408973693848,
-43.0739288330078,-57.5752906799316,
-42.6536560058594,-32.8769035339356,
-34.5647315979004,-6.32860517501831,
-31.5197219848633,-1.66447627544403,
-35.3248596191406,-24.1992568969727,
-28.8125762939453,-56.0803909301758,
-2.99480772018433,-66.7126083374023,
17.7161064147949,-42.5176925659180,
4.51289463043213,-6.43388509750366,
-32.6230812072754,4.10728502273560,
-44.1135406494141,-20.1108837127686,
-3.29436826705933,-47.6750564575195,
50.7623786926270,-50.1467628479004,
61.5898551940918,-35.0988235473633,
25.8707199096680,-25.1655178070068,
-5.31623077392578,-20.6105079650879,
4.71373271942139,-4.36166000366211,
29.1700210571289,21.9693660736084,
25.9819068908691,26.2226428985596,
-0.840948462486267,-4.83963775634766,
-14.1414585113525,-33.0349693298340,
-1.74769341945648,-24.3434467315674,
9.50913333892822,3.16164398193359,
-4.39516925811768,10.4316272735596,
-30.0123310089111,-2.86347627639771,
-34.0228424072266,5.62220954895020,
-12.2321386337280,44.1112823486328,
6.39996433258057,64.1962127685547,
-2.60243415832520,33.4443130493164,
-26.1741580963135,-11.1336536407471,
-32.1564636230469,-14.1180381774902,
-2.96463894844055,17.8270301818848,
38.2861137390137,24.3085632324219,
44.3944587707520,-11.3621044158936,
0.580600261688232,-35.2464599609375,
-48.4574737548828,-9.26966667175293,
-49.5365982055664,29.7049007415772,
-2.90711307525635,26.1275997161865,
33.7244415283203,-16.1868457794189,
17.7424545288086,-40.7953872680664,
-25.4195346832275,-19.0176277160645,
-39.5726394653320,21.0309867858887,
-14.6004247665405,41.5409393310547,
3.48011350631714,37.6811065673828,
-13.5673961639404,22.9388542175293,
-41.0766639709473,1.18313741683960,
-39.9234619140625,-25.0212726593018,
-11.9350290298462,-38.6912727355957,
10.6037206649780,-37.5980491638184,
14.9564704895020,-40.1575202941895,
19.9399356842041,-54.8391876220703,
39.4852027893066,-55.5254402160645,
57.3306121826172,-14.8583641052246,
56.0297660827637,46.0576667785645,
38.6274261474609,76.9607238769531,
21.2889995574951,57.9670562744141,
9.00158500671387,20.8448066711426,
-4.12891054153442,3.51409816741943,
-18.4520492553711,-1.73721706867218,
-25.0076828002930,-17.4836921691895,
-19.7669086456299,-33.8656044006348,
-9.03477096557617,-23.8932628631592,
1.84384965896606,14.6352195739746,
14.1424398422241,46.2628059387207,
20.7426624298096,46.0847511291504,
15.7944879531860,26.1939296722412,
-1.41017723083496,13.1872158050537,
-17.9826927185059,19.0532627105713,
-21.6263732910156,28.9887161254883,
-13.6278429031372,31.7482910156250,
-9.85660171508789,22.6640663146973,
-22.1106700897217,4.06186628341675,
-41.0024108886719,-16.8605651855469,
-43.2226867675781,-26.3987407684326,
-14.1603097915649,-11.8529109954834,
31.4378299713135,11.7533798217773,
51.5751075744629,21.3071613311768,
20.9662532806397,15.5503072738647,
-36.7314033508301,14.9562044143677,
-68.3960647583008,25.2539997100830,
-52.7399406433106,21.8587093353272,
-20.2203235626221,-19.6317138671875,
-7.00431108474731,-77.8580703735352,
-6.16340923309326,-99.9176788330078,
7.61099624633789,-67.1661453247070,
34.6952743530273,-13.9823493957520,
45.6983833312988,10.8646011352539,
30.2334117889404,1.07702994346619,
16.3068542480469,-19.2022132873535,
27.6008663177490,-29.6362915039063,
49.2563056945801,-29.8083000183105,
52.0597305297852,-21.8518333435059,
39.6790466308594,-5.55206060409546,
35.6211357116699,13.7171707153320,
39.5904655456543,18.4088497161865,
29.8345317840576,0.401751518249512,
6.78718948364258,-25.8690319061279,
2.07355594635010,-36.4980621337891,
26.3713893890381,-23.4552021026611,
52.2779464721680,5.79641151428223,
41.6577453613281,37.1605186462402,
0.202260017395020,53.0068626403809,
-34.6702346801758,37.1537933349609,
-43.1099853515625,3.84403038024902,
-31.7464752197266,-17.1240425109863,
-13.5913276672363,-7.38265800476074,
11.6244182586670,13.5248546600342,
32.6112442016602,9.01459407806397,
25.6976566314697,-21.5543289184570,
-8.51901531219482,-40.3396377563477,
-36.8817291259766,-29.6902160644531,
-36.0026588439941,-16.7322444915772,
-19.0668334960938,-31.6558418273926,
-14.7124681472778,-53.6104927062988,
-30.9472942352295,-39.6355247497559,
-43.2671394348145,6.25730895996094,
-27.6045742034912,31.9176692962647,
10.2630729675293,3.74181842803955,
41.3475227355957,-41.5458869934082,
44.0642509460449,-47.5012474060059,
8.89633941650391,-17.6837768554688,
-39.2568244934082,1.25187659263611,
-48.1284294128418,-16.7896499633789,
0.727260351181030,-39.2972831726074,
59.7442932128906,-28.2508182525635,
58.2243041992188,5.15381050109863,
-6.42410135269165,24.5703582763672,
-53.7179679870606,18.9521007537842,
-26.2447586059570,7.29267454147339,
32.1135368347168,5.65342569351196,
32.7694740295410,4.78987026214600,
-24.5938873291016,-8.07321453094482,
-50.9169883728027,-27.3086719512939,
8.54994392395020,-28.0667381286621,
86.6952743530273,2.89674258232117,
87.6276321411133,46.8439216613770,
11.0442905426025,67.3836212158203,
-52.9148750305176,48.1240043640137,
-43.6537666320801,5.33320808410645,
0.266660332679749,-18.8777065277100,
11.9362268447876,-2.50428295135498,
-10.3466091156006,26.7192115783691,
-22.8641490936279,31.9746513366699,
-7.33751344680786,14.9037466049194,
7.43901634216309,1.77395200729370,
-5.04552698135376,1.87590444087982,
-28.2973098754883,1.29927909374237,
-34.7154960632324,-5.76734018325806,
-30.4692916870117,-0.805100381374359,
-30.5898532867432,18.6624832153320,
-34.2402572631836,15.1021366119385,
-25.3849124908447,-33.6154975891113,
-5.89429569244385,-83.6421737670898,
0.921897828578949,-70.2232589721680,
-19.6841926574707,-7.44652986526489,
-42.1393051147461,23.9474315643311,
-34.1073493957520,-17.5919628143311,
-0.553272962570190,-71.8332748413086,
27.5165786743164,-60.3696479797363,
28.4419918060303,1.04970455169678,
10.1572093963623,31.9756793975830,
-3.44223022460938,0.236305117607117,
4.51842355728149,-42.2117919921875,
33.2919044494629,-38.9746932983398,
64.8162307739258,0.696115732192993,
76.5182723999023,29.5952663421631,
58.5349693298340,34.1677398681641,
23.4906654357910,38.0060043334961,
-4.21184825897217,48.8123474121094,
-10.6534729003906,46.2552986145020,
-5.02529239654541,23.6090583801270,
1.24106907844543,4.79284906387329,
7.00441884994507,7.86409950256348,
12.7780714035034,31.6987724304199,
11.0158348083496,55.0059051513672,
4.10728883743286,55.7738380432129,
-2.16280198097229,33.5248718261719,
-5.24280405044556,7.25576210021973,
-11.4410266876221,-0.841269850730896,
-19.8435344696045,21.2068557739258,
-12.1928787231445,44.5760383605957,
19.7216148376465,29.2542076110840,
48.0296401977539,-17.5587329864502,
39.5446777343750,-36.6149864196777,
0.403678894042969,-0.0616161823272705,
-21.3452224731445,43.3744659423828,
-4.10370349884033,27.7338199615479,
14.3953151702881,-32.3230476379395,
-6.62401390075684,-55.8323554992676,
-51.5302619934082,-13.0215721130371,
-68.4861984252930,24.1910400390625,
-40.3283500671387,-12.5171298980713,
0.603736817836762,-81.0225677490234,
18.9375000000000,-77.4388275146484,
15.0258493423462,15.3126802444458,
7.87870550155640,96.5192871093750,
4.05414867401123,82.4496459960938,
1.13328599929810,10.5403556823730,
2.59418010711670,-24.0226764678955,
6.16395044326782,5.41498661041260,
1.96397960186005,33.4217567443848,
-15.2014045715332,6.09264945983887,
-25.6825542449951,-49.9669837951660,
-15.5822448730469,-71.3946380615234,
-5.56614828109741,-37.8089523315430,
-14.8108987808228,10.4372901916504,
-25.4629230499268,27.8143596649170,
-2.60002088546753,11.8667736053467,
47.1909790039063,-11.0733919143677,
74.2271347045898,-5.87399816513062,
46.3823966979981,35.8967819213867,
-3.31638646125793,80.9979019165039,
-21.1567535400391,78.6809692382813,
-3.27676916122437,23.0296401977539,
14.7806196212769,-38.0445861816406,
21.2312297821045,-53.9308547973633,
27.1830673217773,-22.8823699951172,
30.5189609527588,10.9605550765991,
9.62324523925781,18.2777976989746,
-34.1459121704102,12.3631467819214,
-58.2938919067383,7.05680370330811,
-38.0560913085938,-8.97752380371094,
1.09778523445129,-40.8865737915039,
16.5014400482178,-63.4943122863770,
11.5266323089600,-49.8835487365723,
15.0130805969238,-17.5449695587158,
27.9447040557861,-5.26827621459961,
21.3709716796875,-19.4459991455078,
-10.8588705062866,-26.7416419982910,
-19.4277782440186,-4.47569751739502,
23.2170314788818,23.2571926116943,
78.7103271484375,28.9813728332520,
85.7932891845703,12.6144227981567,
33.3186416625977,-0.355303347110748,
-26.5128326416016,0.511325716972351,
-47.4530067443848,8.16593360900879,
-36.1932334899902,19.8059463500977,
-28.3343753814697,33.9801559448242,
-39.7119636535645,32.7941017150879,
-53.5040931701660,-0.00750690698623657,
-47.5870552062988,-45.4515304565430,
-14.5370855331421,-60.4136581420898,
34.4099044799805,-30.8929824829102,
69.3175277709961,11.1915779113770,
61.2680282592773,20.1426239013672,
12.7508516311646,-4.11873626708984,
-33.1618957519531,-28.6111564636230,
-33.6242828369141,-31.1621303558350,
7.20937061309814,-23.9116458892822,
44.0754127502441,-20.8854064941406,
42.8486480712891,-24.3719196319580,
12.7246770858765,-30.8359127044678,
-6.84861612319946,-39.6710472106934,
1.05466032028198,-42.3672485351563,
20.0868587493897,-26.5754146575928,
28.4215373992920,9.08666133880615,
23.3270950317383,35.6540031433106,
11.2633857727051,23.3776550292969,
2.74161434173584,-18.9787406921387,
-1.48473346233368,-55.2184677124023,
-5.00886726379395,-52.3070755004883,
-9.13204002380371,-20.0346546173096,
-13.9338493347168,14.5333509445190,
-11.4994831085205,39.7588920593262,
-3.60448074340820,58.8630790710449,
0.570452630519867,68.8321304321289,
-4.23782444000244,61.2709655761719,
-9.34057617187500,36.7095451354981,
-0.203566938638687,20.7369689941406,
20.3893642425537,30.4562377929688,
24.8674640655518,52.6931228637695,
-1.02836501598358,51.5528450012207,
-34.8892211914063,10.0154113769531,
-41.8228607177734,-47.8477783203125,
-14.3823480606079,-79.5209808349609,
20.1106700897217,-69.5436096191406,
34.6865615844727,-34.5251655578613,
29.4923915863037,-2.95800852775574,
16.8301906585693,5.30361175537109,
3.57130837440491,-0.662567138671875,
-11.8445968627930,-4.79968833923340,
-22.4874687194824,1.80827224254608,
-18.0186824798584,18.5219726562500,
-5.71600198745728,36.7316856384277,
-0.837527394294739,50.0014953613281,
-8.82645034790039,47.4731369018555,
-15.0139617919922,26.4767360687256,
-7.63441801071167,-1.57991003990173,
2.87864398956299,-11.4620351791382,
2.94874095916748,12.0700626373291,
-6.62364578247070,42.1614646911621,
-14.4694833755493,35.3589439392090,
-18.9930572509766,-12.0690212249756,
-33.0996589660645,-56.8962020874023,
-49.4827384948731,-53.5203170776367,
-39.1987228393555,-14.6535968780518,
5.98569250106812,18.0740871429443,
50.4625129699707,31.2214412689209,
47.6833839416504,42.3767051696777,
-2.04143285751343,57.5479202270508,
-48.3342437744141,54.8903617858887,
-52.4488983154297,23.8576717376709,
-24.8295631408691,-4.95689487457275,
1.44967663288116,2.18828368186951,
18.9927310943604,26.5480384826660,
35.8897171020508,32.2354965209961,
42.7783508300781,14.3724069595337,
17.6538467407227,-0.344295203685761,
-32.0853424072266,-2.16229128837585,
-59.8914718627930,-10.9916057586670,
-38.6306915283203,-29.1540660858154,
2.10834527015686,-24.3380527496338,
11.6187534332275,12.1128387451172,
-9.12110614776611,41.1459999084473,
-20.1050949096680,19.7438468933105,
3.42498779296875,-31.1932640075684,
35.8372688293457,-48.1339149475098,
37.4977378845215,-16.2752246856689,
14.2631788253784,13.6094932556152,
4.68288755416870,-6.06528997421265,
19.7914676666260,-49.6931343078613,
31.8112850189209,-58.1871070861816,
12.3991289138794,-19.1915283203125,
-26.2648468017578,20.7105636596680,
-43.0359268188477,19.2103042602539,
-19.7342948913574,-15.6459894180298,
8.28163719177246,-45.1255035400391,
-3.41691207885742,-45.7527236938477,
-45.5722274780273,-26.3981723785400,
-67.5539703369141,-5.11540365219116,
-40.0197944641113,9.92541599273682,
4.62260818481445,10.9238958358765,
13.1594524383545,-6.47897768020630,
-13.1572017669678,-32.2134780883789,
-24.6278991699219,-44.7795677185059,
4.49210548400879,-29.5393657684326,
34.0030937194824,2.47638440132141,
17.3683605194092,23.1119556427002,
-27.6861972808838,17.9479942321777,
-41.5196266174316,-1.26227211952209,
-5.08030176162720,-7.24178171157837,
37.4633216857910,5.41916751861572,
39.2687454223633,26.4927406311035,
7.17947196960449,36.2757034301758,
-18.5671253204346,23.1020088195801,
-15.3601036071777,-9.07473468780518,
5.95968198776245,-41.6351966857910,
31.4453773498535,-47.1648979187012,
50.0982894897461,-15.8068161010742,
50.7527313232422,32.0165557861328,
25.9567260742188,60.6387176513672,
-5.55395555496216,50.4041366577148,
-13.4237995147705,18.9679431915283,
8.70766162872315,1.44179773330688,
30.2007427215576,11.7754945755005,
22.8461227416992,37.8062438964844,
2.10992646217346,56.8193054199219,
-2.42001914978027,58.2979202270508,
8.91879558563232,50.6891250610352,
7.90417385101318,43.2637252807617,
-20.2634220123291,37.2910614013672,
-45.4265022277832,23.9678745269775,
-33.3695144653320,0.460813701152802,
5.98875522613525,-18.7419586181641,
24.3093109130859,-13.4589109420776,
-3.25367784500122,14.3147048950195,
-46.1121253967285,39.2381477355957,
-54.5207252502441,34.9507217407227,
-20.7441463470459,3.52755188941956,
17.2460842132568,-21.6956729888916,
17.5042209625244,-19.6992549896240,
-18.5889205932617,1.85813653469086,
-48.5314445495606,17.3071308135986,
-42.3726348876953,11.7883987426758,
-8.82049751281738,-13.6624526977539,
19.5452747344971,-41.1758613586426,
24.8344860076904,-53.1673889160156,
21.3681335449219,-40.5651321411133,
27.9983196258545,-17.5120792388916,
40.9282150268555,-6.22143745422363,
30.6314468383789,-12.8667621612549,
-6.39168405532837,-13.0593118667603,
-33.8360252380371,10.9832696914673,
-21.1078567504883,41.6948966979981,
10.6863708496094,41.3928031921387,
13.0684480667114,9.91504478454590,
-27.1309013366699,-8.99863243103027,
-63.2914123535156,9.18366241455078,
-48.2586631774902,30.5209655761719,
1.91757130622864,15.2714900970459,
33.5151214599609,-24.4057502746582,
28.7117824554443,-39.6518402099609,
6.21809625625610,-14.0000629425049,
-14.9348821640015,13.9588537216187,
-36.8957481384277,7.87682390213013,
-56.6015739440918,-16.6737232208252,
-49.1316337585449,-29.5906085968018,
-10.6754102706909,-30.3790168762207,
15.8018474578857,-35.9543380737305,
0.146682977676392,-44.5610923767090,
-26.2481708526611,-39.8401184082031,
-11.6047687530518,-27.2120075225830,
39.0897178649902,-28.6224174499512,
59.9864349365234,-41.1031570434570,
17.4398193359375,-39.3281745910645,
-33.6306838989258,-15.0669822692871,
-20.3830471038818,2.34838652610779,
42.3306045532227,-7.09368133544922,
76.7434005737305,-22.1060123443604,
37.8862113952637,-8.26288795471191,
-33.8496398925781,24.1661491394043,
-64.1224441528320,31.9040603637695,
-28.4468231201172,4.31263732910156,
29.1029930114746,-24.0822620391846,
51.3746452331543,-23.1441898345947,
23.1752758026123,-8.18179798126221,
-21.2420520782471,-7.65520381927490,
-35.5519447326660,-17.4800872802734,
-8.76188087463379,-13.1710147857666,
26.8786487579346,13.1643695831299,
24.4834938049316,36.4766883850098,
-20.3131561279297,39.7730369567871,
-63.7796401977539,29.6726512908936,
-73.6055068969727,21.1457405090332,
-57.4700469970703,10.1947259902954,
-36.6764411926270,-10.3494844436646,
-16.5289001464844,-26.4763278961182,
6.46349954605103,-19.2968826293945,
22.9977855682373,8.65141582489014,
13.9115619659424,34.4714279174805,
-14.7821187973022,38.4836769104004,
-29.9336929321289,25.6762351989746,
-23.6916103363037,9.24692058563232,
-24.9807872772217,-3.74392247200012,
-48.0171775817871,-15.5978279113770,
-63.8047523498535,-25.3587455749512,
-37.2472801208496,-28.7571697235107,
10.8628177642822,-26.3509788513184,
29.7722702026367,-14.9280853271484,
9.79355335235596,6.40769481658936,
-9.67352676391602,27.6120643615723,
-0.792338848114014,27.8775539398193,
16.4868297576904,-0.747028827667236,
11.6793451309204,-31.6126117706299,
-1.82407331466675,-29.8916110992432,
5.74009323120117,7.78619050979614,
26.5382843017578,48.8251762390137,
21.1702175140381,63.3713150024414,
-18.7438087463379,53.1030960083008,
-52.6468391418457,40.7540321350098,
-51.9402732849121,30.3308792114258,
-31.3476200103760,10.4174327850342,
-23.9550952911377,-21.5849914550781,
-23.9964523315430,-51.9201202392578,
-8.71966552734375,-68.1494674682617,
22.8447875976563,-62.2169227600098,
44.3269653320313,-34.7897949218750,
44.4592666625977,3.57010865211487,
44.6538810729981,26.3548488616943,
59.1466598510742,20.6468296051025,
68.0276947021484,2.98795413970947,
50.5927963256836,-3.63957524299622,
23.1882266998291,-1.00188553333282,
10.3866891860962,-12.4888124465942,
10.4851007461548,-41.8502693176270,
-2.67009210586548,-53.7675743103027,
-36.2957687377930,-27.0717506408691,
-63.2582511901856,5.80871391296387,
-59.8995933532715,6.21384334564209,
-35.5267295837402,-14.4202022552490,
-11.5247364044189,-19.5065040588379,
1.49081254005432,-10.4994125366211,
5.38476181030273,-23.9183349609375,
-1.87063765525818,-65.7144927978516,
-16.0267066955566,-77.3405609130859,
-15.2264804840088,-24.7190322875977,
5.86282920837402,49.0366401672363,
22.3395748138428,72.8507614135742,
-0.0616267882287502,38.1204643249512,
-45.0931472778320,9.36424732208252,
-62.8287010192871,21.3434848785400,
-25.6797180175781,42.6356086730957,
30.6211853027344,34.6152534484863,
50.3092193603516,7.69220972061157,
24.3277244567871,1.79583668708801,
-10.0099792480469,21.4462985992432,
-25.9528694152832,39.9816284179688,
-24.7208271026611,29.1091823577881,
-16.1386623382568,-9.09158992767334,
1.89268100261688,-52.2350311279297,
24.6387329101563,-72.4885940551758,
40.4005928039551,-48.0009193420410,
37.1226921081543,8.79227638244629,
14.8839807510376,49.3012466430664,
-17.5376796722412,22.5643711090088,
-47.1591606140137,-50.1665420532227,
-53.5124549865723,-89.9946746826172,
-24.0261230468750,-56.6866798400879,
23.6754798889160,7.63292980194092,
46.4005622863770,36.7901344299316,
21.7150611877441,28.4492168426514,
-12.9258890151978,26.1742687225342,
-13.0083208084106,48.6417388916016,
5.94127893447876,63.5724754333496,
-6.47048950195313,42.5013275146484,
-56.1386871337891,10.3600540161133,
-84.7866134643555,-1.54079198837280,
-52.8045158386231,-6.82701253890991,
5.74050521850586,-29.2978916168213,
30.8621749877930,-59.3750648498535,
20.2560844421387,-64.8739318847656,
23.9807567596436,-43.0066680908203,
56.2850761413574,-25.5802898406982,
74.5699462890625,-25.8030357360840,
52.1974601745606,-28.1998901367188,
17.6023902893066,-25.5169696807861,
11.0327262878418,-29.0177669525147,
22.8426742553711,-36.1979064941406,
20.8015003204346,-19.0102882385254,
5.27447652816773,33.3515090942383,
-0.542521476745606,69.2026290893555,
4.83760261535645,36.9248733520508,
-1.97451198101044,-32.7316474914551,
-25.2038688659668,-59.2439880371094,
-35.3063812255859,-14.9878711700439,
-14.5077896118164,45.8599357604981,
9.02755928039551,61.1949958801270,
3.82856655120850,34.2416687011719,
-20.9106826782227,3.92827844619751,
-35.3527374267578,-9.85547542572022,
-33.9207382202148,-21.0266323089600,
-28.6465167999268,-33.9284629821777,
-16.4066543579102,-42.5875549316406,
6.84621953964233,-49.0745735168457,
28.9400749206543,-62.8294410705566,
23.5531749725342,-65.6303710937500,
-6.55241680145264,-34.9170227050781,
-22.7322673797607,12.9891433715820,
-1.42224717140198,28.7754383087158,
33.2697868347168,-3.88123464584351,
43.4885139465332,-38.8860054016113,
28.3181037902832,-37.1231613159180,
9.71497154235840,-8.06321048736572,
-9.41718578338623,4.85354375839233,
-38.8331451416016,-10.0559482574463,
-60.6425285339356,-21.7508411407471,
-44.1308364868164,-16.2075099945068,
9.26461315155029,-7.44550323486328,
55.7555084228516,-3.61355209350586,
56.8888893127441,10.4765968322754,
28.8320655822754,37.3448982238770,
12.1268367767334,47.3595504760742,
17.2489948272705,23.4637451171875,
24.7878017425537,-10.1898908615112,
23.0415458679199,-18.1627120971680,
22.0734214782715,-9.59362792968750,
23.8392925262451,-18.4099788665772,
17.6340732574463,-46.2576828002930,
11.2045726776123,-56.2984695434570,
22.5522785186768,-26.9654445648193,
51.4474105834961,13.7997331619263,
64.6626052856445,30.5337028503418,
38.5711784362793,26.7981109619141,
-4.27236080169678,26.2575263977051,
-25.6101131439209,23.3689994812012,
-19.0603103637695,0.980816841125488,
-14.9445304870605,-31.6465129852295,
-26.7737655639648,-43.8932800292969,
-31.3856372833252,-27.8592815399170,
-19.1479358673096,-7.15910911560059,
-7.69893789291382,-4.22653055191040,
-11.9610919952393,-13.4274730682373,
-15.7516679763794,-17.1787452697754,
2.62096166610718,-10.8903923034668,
29.7244701385498,1.33244681358337,
32.4582252502441,19.1188125610352,
12.9639625549316,31.4353504180908,
3.52654552459717,12.9250946044922,
14.9410552978516,-30.7428588867188,
18.7710304260254,-53.8874816894531,
-7.16899204254150,-28.4891586303711,
-31.8105831146240,10.8659124374390,
-14.2904958724976,10.5057201385498,
29.9136543273926,-22.0230541229248,
49.1385993957520,-24.9058570861816,
24.6216945648193,21.9792251586914,
-3.43726634979248,66.6117248535156,
5.58642673492432,54.2618446350098,
36.4681053161621,10.8544187545776,
44.8394355773926,-2.27449703216553,
15.4342870712280,15.8467359542847,
-21.5179119110107,14.4888086318970,
-33.4208984375000,-18.8911056518555,
-22.0453281402588,-41.5078430175781,
-5.46940422058106,-24.4585876464844,
3.24456453323364,3.75792598724365,
-1.78901863098145,3.36948633193970,
-17.7453861236572,-22.4794349670410,
-30.4525413513184,-42.3333930969238,
-26.5089130401611,-46.5897521972656,
-10.7810068130493,-43.7135925292969,
2.17316794395447,-25.9926471710205,
2.34905552864075,16.0562019348145,
-13.1884899139404,51.8427200317383,
-36.5549621582031,33.4872474670410,
-59.3617897033691,-26.4161224365234,
-62.7421607971191,-53.1288528442383,
-30.1581821441650,-11.7672348022461,
21.2822265625000,39.6434860229492,
42.4658241271973,27.8786315917969,
12.0112342834473,-28.1969089508057,
-28.3969573974609,-41.7893714904785,
-26.5958957672119,16.6796627044678,
2.60887956619263,75.8216094970703,
4.99997854232788,65.1810913085938,
-25.2647533416748,9.17235374450684,
-34.2339897155762,-18.3428840637207,
11.7370681762695,-1.29936170578003,
68.2285919189453,10.7835655212402,
70.1070632934570,-11.4950389862061,
20.1127490997314,-32.8267707824707,
-23.4878940582275,-16.6351203918457,
-28.4120292663574,14.5037975311279,
-11.7143459320068,18.4737606048584,
7.67842245101929,-3.80611586570740,
27.6941089630127,-9.63928604125977,
39.9076805114746,20.0945167541504,
18.6257553100586,47.1787681579590,
-29.6009559631348,33.2314453125000,
-50.1807823181152,-4.17571735382080,
-12.0329799652100,-19.0210514068604,
51.2686195373535,3.14695620536804,
72.7094116210938,33.4815826416016,
36.2375488281250,39.7379417419434,
-8.17308044433594,24.1461601257324,
-15.4559383392334,10.8905696868896,
3.76846623420715,9.20635604858398,
12.1431350708008,2.45399522781372,
-0.755950808525085,-19.0515975952148,
-18.4446678161621,-37.1590270996094,
-24.2377796173096,-32.3283729553223,
-15.4915075302124,-6.00938606262207,
1.35773050785065,16.6677188873291,
13.0689449310303,16.7275581359863,
6.27205324172974,5.11520338058472,
-22.9420433044434,3.76047897338867,
-53.3346366882324,10.8269720077515,
-55.1486129760742,-0.175188064575195,
-19.9735851287842,-32.1219596862793,
25.5088882446289,-49.3720970153809,
39.1414794921875,-20.7929801940918,
13.1914720535278,34.8883132934570,
-25.1185245513916,54.2133255004883,
-44.1225051879883,9.78859519958496,
-33.2127761840820,-53.1259994506836,
-11.5629014968872,-70.7483596801758,
-3.12985682487488,-34.9189071655273,
-16.2958965301514,4.94578075408936,
-37.2872352600098,13.0179443359375,
-46.9389801025391,0.543001174926758,
-36.3150215148926,-3.60552549362183,
-14.4049339294434,-2.17533659934998,
7.32256841659546,-17.3948230743408,
24.9304523468018,-40.0349807739258,
40.1436576843262,-35.2856941223145,
48.1445770263672,8.99812889099121,
34.5413818359375,54.0545921325684,
-0.772273659706116,56.3534317016602,
-36.4914665222168,15.8221635818481,
-51.2654533386231,-23.6681995391846,
-45.8206062316895,-31.8836097717285,
-35.4423103332520,-21.9176845550537,
-30.9843463897705,-15.7886819839478,
-26.7852611541748,-12.4357261657715,
-18.6430034637451,1.32275307178497,
-11.4729261398315,22.4148464202881,
-6.58150243759155,26.6200122833252,
4.75096368789673,2.60303330421448,
21.8446521759033,-27.6110267639160,
29.8447360992432,-37.5734977722168,
12.7891798019409,-25.8518104553223,
-16.7507324218750,-14.6085567474365,
-31.9927825927734,-16.7728614807129,
-23.7676277160645,-26.1831321716309,
-13.4629783630371,-28.9748458862305,
-17.5436840057373,-21.7964057922363,
-25.3409118652344,-9.47179031372070,
-19.3559169769287,7.04282760620117,
4.39094352722168,25.0092449188232,
24.1744174957275,36.5512847900391,
24.7746810913086,34.2876510620117,
10.1817684173584,22.7209091186523,
-2.09056782722473,9.77470874786377,
-1.45383894443512,-2.64695572853088,
8.88820362091065,-17.7726783752441,
17.5262565612793,-29.2615432739258,
16.6504058837891,-30.1246643066406,
9.99406909942627,-22.2568435668945,
9.15954399108887,-20.6712493896484,
16.6776561737061,-35.5602073669434,
17.6689186096191,-49.8052101135254,
-0.124305009841919,-43.1905403137207,
-31.3764610290527,-14.2047252655029,
-50.3171310424805,19.8799953460693,
-42.7161026000977,43.8790702819824,
-16.6010189056397,54.3049964904785,
7.61449575424194,53.7220001220703,
18.2995510101318,42.7155952453613,
15.7303485870361,29.9052391052246,
3.30816602706909,21.6548881530762,
-13.4750308990479,14.6014642715454,
-24.7102584838867,-3.61718964576721,
-15.7689609527588,-31.7340488433838,
8.67728424072266,-44.4627914428711,
28.4399375915527,-20.2733955383301,
24.3602180480957,24.6989288330078,
-4.40693473815918,50.4429855346680,
-40.6211547851563,43.7057571411133,
-60.8152427673340,24.1038532257080,
-51.6635513305664,14.5287990570068,
-18.9008045196533,16.5647754669189,
11.0814304351807,21.0608139038086,
11.4870901107788,25.1671657562256,
-16.2704696655273,28.8431091308594,
-34.3041534423828,19.3210773468018,
-9.17287158966065,-5.05002307891846,
34.3949508666992,-26.2362232208252,
39.1906738281250,-22.9162120819092,
-10.4042835235596,-6.39187526702881,
-60.0718040466309,-6.71410131454468,
-51.5711898803711,-26.3233184814453,
1.88028788566589,-33.3153724670410,
31.8886470794678,-4.95376777648926,
7.80677700042725,32.3653678894043,
-26.8172302246094,42.6995086669922,
-21.6154136657715,25.1967144012451,
9.40102767944336,4.39471054077148,
23.4069442749023,0.827125787734985,
16.2923030853272,8.27277565002441,
22.1627845764160,14.7009668350220,
45.5265312194824,17.4888420104980,
48.7880439758301,11.4360008239746,
12.8021945953369,-4.20072507858276,
-18.5391101837158,-18.3115005493164,
-3.25066661834717,-13.5956058502197,
33.5895347595215,15.0654602050781,
34.3906669616699,45.2097587585449,
-5.32344388961792,57.1405982971191,
-28.6717548370361,53.6021499633789,
-3.69144701957703,41.9423141479492,
26.0855331420898,19.3427886962891,
10.3449611663818,-12.5860376358032,
-32.2117919921875,-40.9524612426758,
-46.3334007263184,-47.9413261413574,
-22.1557235717773,-26.7823352813721,
-5.15534877777100,7.27663707733154,
-25.6423435211182,35.4445724487305,
-53.7578163146973,38.9189262390137,
-52.0872268676758,6.26904487609863,
-23.5038089752197,-46.8521728515625,
-4.59956216812134,-75.4360504150391,
-7.54377317428589,-46.2471733093262,
-12.5743751525879,14.5048198699951,
-11.5680437088013,40.7325897216797,
-13.6428747177124,9.75805473327637,
-19.6418228149414,-28.0699443817139,
-21.3517990112305,-19.4800529479980,
-11.5909070968628,26.4558773040772,
-1.98434090614319,46.4639358520508,
-5.44510555267334,13.8997001647949,
-17.3184432983398,-32.5678901672363,
-19.2519645690918,-46.9404106140137,
-0.377580642700195,-28.7346439361572,
32.5709342956543,-10.6694374084473,
57.1537857055664,-5.47488069534302,
49.3441734313965,-4.03987598419189,
-1.12282454967499,-0.550701916217804,
-59.4372406005859,-5.69640302658081,
-70.6627655029297,-20.4119739532471,
-18.5761432647705,-21.3939094543457,
46.4271888732910,-2.99976873397827,
58.1496925354004,12.6147766113281,
8.64320564270020,0.701940774917603,
-46.2312583923340,-29.6823825836182,
-53.9023857116699,-42.0130615234375,
-21.8371086120605,-13.4922199249268,
5.87696313858032,28.3236827850342,
5.94221830368042,38.7624893188477,
-11.0642156600952,12.3877143859863,
-31.5872726440430,-15.2621126174927,
-48.5835380554199,-9.92749881744385,
-52.1692924499512,19.2413692474365,
-30.5405387878418,32.3593444824219,
8.48472023010254,4.54449844360352,
30.0307407379150,-35.5000381469727,
16.5333919525147,-45.8366889953613,
-3.40720605850220,-23.3253383636475,
8.89410495758057,-6.86300325393677,
50.9149894714356,-12.1386651992798,
74.8327713012695,-10.6329660415649,
49.1010360717773,22.1392288208008,
2.31546115875244,60.5398635864258,
-19.9320659637451,53.6093864440918,
-15.0359401702881,2.23644137382507,
-13.7041397094727,-32.4360580444336,
-31.4946689605713,-16.1493759155273,
-46.8925476074219,9.04705524444580,
-38.6105041503906,-10.0629224777222,
-14.7543811798096,-59.0376091003418,
5.27578067779541,-77.0368576049805,
13.2802753448486,-50.0286331176758,
15.7053432464600,-27.5748214721680,
12.8872365951538,-42.2545166015625,
1.43572449684143,-52.8838653564453,
-8.91621971130371,-16.5342254638672,
-11.2796220779419,45.6332283020020,
-15.0590772628784,67.0620498657227,
-33.4717292785645,27.6702060699463,
-53.6767578125000,-22.0998878479004,
-55.7864570617676,-33.6485939025879,
-32.5689735412598,-14.2183399200439,
-1.07915735244751,1.35022163391113,
20.4794063568115,3.22500896453857,
27.2603588104248,4.08217763900757,
20.2507133483887,5.67772102355957,
-0.993671178817749,-2.09979414939880,
-24.3460350036621,-21.0603027343750,
-21.9401168823242,-43.5563468933106,
7.72812843322754,-59.2545852661133,
32.6989479064941,-66.4054260253906,
25.6400604248047,-58.9864921569824,
6.15242576599121,-28.2543125152588,
10.9866437911987,15.0550603866577,
37.8734092712402,39.0373840332031,
51.9556121826172,31.2441768646240,
37.2522926330566,17.4148311614990,
15.5949096679688,22.3525753021240,
5.69095516204834,39.6047477722168,
-3.52940368652344,42.8443145751953,
-28.5643711090088,23.5651245117188,
-47.7718505859375,5.84045743942261,
-31.8336830139160,2.07958650588989,
10.8419618606567,-0.245860248804092,
42.3845634460449,-8.52237701416016,
44.8526039123535,-4.80338907241821,
31.8554668426514,25.6679801940918,
13.9826879501343,56.3713912963867,
-7.83766269683838,48.8296318054199,
-23.4671173095703,3.09610319137573,
-17.8845634460449,-31.0281486511230,
6.48580789566040,-25.4797706604004,
15.1169643402100,-8.74182033538818,
-10.2072000503540,-15.2092618942261,
-38.5756111145020,-36.3524322509766,
-27.4388885498047,-28.7956008911133,
11.6289024353027,18.9997558593750,
32.3725090026856,64.2457199096680,
20.1611347198486,60.3396682739258,
11.5100135803223,17.7424621582031,
26.6085243225098,-16.5667610168457,
34.0930252075195,-12.4314527511597,
1.88467049598694,11.1593513488770,
-41.5981712341309,16.8359966278076,
-34.4500808715820,-7.89956665039063,
25.7420215606689,-30.9412841796875,
72.0742568969727,-13.7836942672730,
50.7077484130859,33.7039031982422,
-10.4905357360840,62.2064933776856,
-39.2605056762695,40.9856567382813,
-10.8584260940552,-2.99464702606201,
32.5240516662598,-18.8600883483887,
43.4140167236328,3.23197460174561,
22.2820587158203,22.9983043670654,
-8.07899665832520,7.35840034484863,
-32.2394180297852,-20.0075740814209,
-50.3534622192383,-23.0866012573242,
-57.9515914916992,-10.9540452957153,
-38.5250549316406,-16.4870414733887,
4.69177770614624,-44.2807197570801,
41.5625228881836,-55.5125923156738,
43.3685035705566,-29.6732788085938,
15.6787090301514,6.20448589324951,
-11.0868730545044,15.4051694869995,
-16.2857685089111,7.67606067657471,
-3.35564947128296,12.9038677215576,
-1.11393857002258,31.4991817474365,
-22.4243488311768,32.7630119323731,
-42.6115379333496,2.99613952636719,
-28.2518901824951,-22.6464366912842,
16.6779136657715,-10.0171165466309,
49.3846397399902,26.2613716125488,
32.0309066772461,44.4018135070801,
-17.3469963073730,26.8323764801025,
-40.2770423889160,-9.21292114257813,
-16.8344535827637,-39.7513427734375,
16.7205066680908,-52.8448944091797,
18.3751964569092,-51.4753608703613,
5.32667922973633,-42.6042861938477,
16.9152526855469,-36.9993705749512,
45.8013496398926,-41.9452781677246,
45.7939987182617,-45.4870071411133,
7.81643676757813,-24.8132839202881,
-17.4812564849854,16.0739536285400,
7.46629905700684,39.0600929260254,
43.9846763610840,19.2743206024170,
30.1286983489990,-20.4823722839355,
-26.7084751129150,-42.5007629394531,
-59.6395530700684,-41.2298240661621,
-30.2248649597168,-34.2797470092773,
24.8766746520996,-27.0598087310791,
50.1081809997559,-3.99286055564880,
41.0266151428223,29.6393547058105,
24.2527751922607,35.9158630371094,
8.95869445800781,1.04565644264221,
-9.23060417175293,-34.2612152099609,
-23.7536659240723,-27.3512020111084,
-15.7061052322388,4.11893510818481,
13.4157781600952,10.7984189987183,
37.4630279541016,-20.4428329467773,
35.3419952392578,-44.3827056884766,
14.9182567596436,-30.1273727416992,
-5.31834602355957,-5.09230375289917,
-19.0890598297119,-5.36413669586182,
-26.2910690307617,-19.9372978210449,
-21.2067527770996,-9.27865123748779,
-8.95867919921875,32.2814178466797,
-6.94901609420776,59.6423645019531,
-19.3808555603027,38.1504402160645,
-27.8523616790772,-8.87663173675537,
-9.19222640991211,-32.3242607116699,
27.6344356536865,-20.4579944610596,
44.7059097290039,-7.93856668472290,
25.6551017761230,-23.0270500183105,
-6.42368841171265,-50.4567222595215,
-17.0772438049316,-49.1478576660156,
-6.25766181945801,-7.20895576477051,
-0.311697781085968,34.7634696960449,
-8.60460758209229,28.3992328643799,
-11.2167787551880,-13.4681797027588,
9.39165210723877,-38.1176719665527,
33.3023910522461,-12.3321399688721,
27.3275775909424,30.8516941070557,
-5.39652538299561,34.1709671020508,
-25.9500923156738,-9.29092693328857,
-5.11260032653809,-48.0607948303223,
33.1588706970215,-39.2042160034180,
42.8310317993164,-3.67871189117432,
12.3978166580200,12.0521907806396,
-22.6388835906982,-3.27863407135010,
-30.6346359252930,-17.2893562316895,
-19.4561729431152,-9.62022590637207,
-14.9272127151489,-2.65002322196960,
-21.7692680358887,-27.1939888000488,
-18.0487422943115,-70.7963638305664,
6.65779399871826,-86.7726593017578,
27.9508323669434,-57.7339744567871,
17.5807838439941,-8.27651691436768,
-15.4884262084961,20.4765911102295,
-36.5951843261719,20.2283477783203,
-21.8218498229980,16.4674358367920,
12.7186450958252,25.7311820983887,
30.3713226318359,35.0680313110352,
18.4522895812988,24.4813098907471,
-1.17822825908661,-3.79708075523376,
-2.71181464195251,-29.6541061401367,
10.0109910964966,-36.1204948425293,
16.1048355102539,-26.0568981170654,
7.57834959030151,-12.3336534500122,
1.26852941513062,3.08715796470642,
13.9464874267578,30.3251571655273,
32.6407279968262,64.4223785400391,
23.4287414550781,85.2103347778320,
-21.3213481903076,75.9964599609375,
-68.9912338256836,36.1852416992188,
-76.5771255493164,-5.23091554641724,
-38.0111694335938,-26.5331764221191,
9.55338668823242,-26.2516269683838,
23.9323043823242,-18.8024787902832,
-0.531655192375183,-12.1754817962646,
-36.4415054321289,-5.74139499664307,
-50.3798217773438,-2.43343305587769,
-33.1484870910645,-9.09031105041504,
-2.90901207923889,-23.7504119873047,
15.8884773254395,-25.8418617248535,
12.9270410537720,6.28783988952637,
-0.910936713218689,57.4747657775879,
-12.5012063980103,80.7261962890625,
-20.1280651092529,45.4020500183106,
-29.1038627624512,-19.0047378540039,
-36.4409942626953,-61.0280799865723,
-28.1811275482178,-59.8615264892578,
-4.57267761230469,-47.1285972595215,
7.31921958923340,-49.8941535949707,
-8.80440139770508,-52.7644309997559,
-34.1601104736328,-29.2652206420898,
-35.1669197082520,16.4372844696045,
-5.93948745727539,49.5047035217285,
21.6465644836426,51.2223701477051,
16.6274776458740,38.1774635314941,
-7.86395120620728,25.9377231597900,
-23.8366336822510,11.0282211303711,
-23.2954158782959,-6.59605407714844,
-16.4188156127930,-10.8108243942261,
-7.85451698303223,6.39232254028320,
5.41882228851318,27.2833633422852,
12.2504138946533,30.1037197113037,
1.87737202644348,14.3595418930054,
-11.4228887557983,-7.12059926986694,
2.82882332801819,-25.3087482452393,
42.0811042785645,-39.5189094543457,
59.5677757263184,-33.6055145263672,
23.2469272613525,4.65862035751343,
-26.4046936035156,47.7355499267578,
-29.0846920013428,47.0980262756348,
17.6853828430176,4.22281265258789,
49.1456718444824,-26.5488033294678,
23.4921913146973,-13.5295734405518,
-22.6519241333008,9.54519939422607,
-33.9085884094238,-3.61069703102112,
-13.1892738342285,-38.8164176940918,
-3.23767948150635,-42.9201354980469,
-17.0538444519043,-12.1431255340576,
-21.5687484741211,3.23991799354553,
6.31704092025757,-20.0033397674561,
36.8923492431641,-35.5252990722656,
24.9048709869385,1.48128342628479,
-29.1749534606934,57.4028816223145,
-77.8523788452148,61.4335212707520,
-79.5057678222656,4.79160547256470,
-40.2164268493652,-50.1335487365723,
4.19445943832398,-51.0987205505371,
23.4133262634277,-18.0970859527588,
15.4376125335693,5.82769393920898,
3.81093144416809,10.7472333908081,
9.52586460113525,21.1177406311035,
22.7725429534912,44.2429161071777,
17.7063140869141,56.8791656494141,
-9.83946228027344,43.1468963623047,
-36.5181808471680,14.0849208831787,
-36.6789093017578,-6.67491102218628,
-13.4812355041504,-14.8253593444824,
3.61884498596191,-12.3412122726440,
3.07239580154419,4.18614435195923,
-3.81426906585693,33.7232093811035,
-5.08935832977295,60.9351119995117,
-3.95648908615112,67.9837570190430,
-2.13777518272400,51.7247886657715,
2.52614593505859,33.1098861694336,
12.9372901916504,26.7784881591797,
16.3527221679688,20.4780750274658,
7.20072841644287,1.78377127647400,
2.47150087356567,-19.3922176361084,
14.9097690582275,-18.6121654510498,
34.2923622131348,10.9474830627441,
31.6992321014404,42.5206146240234,
-0.510511875152588,49.9271736145020,
-42.5131187438965,29.9067440032959,
-68.6257781982422,5.29290485382080,
-69.1389160156250,-7.08071231842041,
-46.8033256530762,-7.92840528488159,
-12.3972835540771,-0.564985573291779,
12.5362272262573,12.6337566375732,
5.20355558395386,25.6849689483643,
-27.1975421905518,20.5000133514404,
-44.1898765563965,-0.155163526535034,
-15.8711395263672,-15.8853931427002,
32.1992225646973,-2.69483923912048,
47.7468528747559,34.1006317138672,
13.6053218841553,58.8541374206543,
-33.6444740295410,46.1783370971680,
-48.0274353027344,4.45230579376221,
-27.2220630645752,-31.7657794952393,
-5.16333055496216,-35.8253250122070,
-6.62332677841187,-11.3923978805542,
-23.6403598785400,18.7069473266602,
-38.1599235534668,31.0586891174316,
-37.9723739624023,24.4289054870605,
-22.5442352294922,21.4175739288330,
-2.89379668235779,39.0286178588867,
1.71903276443481,61.5781974792481,
-16.5248699188232,54.5547561645508,
-38.9097785949707,8.85122489929199,
-38.5067367553711,-49.8376770019531,
-16.8604316711426,-79.4154663085938,
-4.47816705703735,-62.5698928833008,
-18.5556793212891,-17.8279094696045,
-34.7840690612793,17.8955421447754,
-16.6995201110840,20.2280845642090,
20.1765861511230,-10.4157085418701,
25.0572280883789,-38.4272613525391,
-9.71717453002930,-26.7552928924561,
-38.1284065246582,20.7511291503906,
-22.4191322326660,54.4530410766602,
11.0688438415527,34.4106063842773,
15.2460660934448,-9.54253768920898,
-6.75525665283203,-16.0176048278809,
-10.7496633529663,24.7348861694336,
12.8505487442017,59.2503433227539,
23.8235893249512,49.9370536804199,
7.80615949630737,16.8485660552979,
-0.763953506946564,4.31796264648438,
26.6626300811768,17.9399394989014,
49.7251739501953,23.1170024871826,
21.9795475006104,11.6839761734009,
-30.2620391845703,-3.18460941314697,
-37.7542495727539,-16.8818073272705,
10.2916755676270,-35.0881195068359,
49.4626960754395,-42.3948478698731,
31.2837352752686,-12.4383678436279,
-8.77354907989502,38.9021949768066,
-13.9533233642578,54.8330116271973,
12.0720186233521,16.7365283966064,
14.9354486465454,-21.0971717834473,
-19.5583248138428,-7.34988021850586,
-56.2632446289063,32.7929344177246,
-65.7108688354492,33.6229896545410,
-59.5085296630859,-18.9828224182129,
-50.9253883361816,-63.4252395629883,
-29.1305122375488,-59.1132011413574,
10.2200260162354,-32.6899375915527,
42.6266822814941,-26.5820159912109,
42.9982261657715,-35.7537460327148,
21.8750820159912,-31.6339073181152,
14.1505517959595,-16.1998138427734,
31.9723281860352,-11.0023775100708,
46.8525657653809,-16.3373088836670,
42.6951866149902,-10.7191877365112,
34.0107688903809,6.54917430877686,
36.6189231872559,16.7820816040039,
46.8439178466797,9.90956687927246,
52.0060043334961,6.52614927291870,
44.6483345031738,21.2058029174805,
19.1965122222900,40.1294174194336,
-15.8137865066528,41.1863937377930,
-45.3858528137207,26.6019191741943,
-42.5865097045898,9.78282070159912,
-10.8042421340942,-11.7663316726685,
8.53113842010498,-34.7111740112305,
-16.4708843231201,-42.0842933654785,
-56.2981033325195,-23.6804485321045,
-48.3281822204590,-3.03810143470764,
11.1627521514893,-3.03303956985474,
58.4793434143066,-13.8734226226807,
44.1823577880859,2.42246580123901,
-1.03659534454346,48.7500915527344,
-17.9922847747803,85.5452804565430,
-4.12859678268433,81.3183593750000,
-14.1671009063721,50.6908607482910,
-64.4900207519531,24.6604213714600,
-98.1537933349609,4.17338848114014,
-66.8325042724609,-21.5670719146729,
-2.42382812500000,-34.5929107666016,
27.3103237152100,-16.3536396026611,
6.27826309204102,12.9263544082642,
-9.42088508605957,11.4028053283691,
15.2405452728271,-22.8247756958008,
49.7474327087402,-44.3455276489258,
50.2242965698242,-21.0412559509277,
24.3316287994385,25.5603637695313,
11.7598390579224,52.4005470275879,
20.6056747436523,48.2074279785156,
21.6995449066162,28.7976722717285,
-3.86420154571533,3.17649936676025,
-24.4562950134277,-23.3660163879395,
-10.5953149795532,-33.2308959960938,
18.8140201568604,-10.4054031372070,
19.9335746765137,24.4309196472168,
-15.6197071075439,30.1612434387207,
-57.0958442687988,1.34728169441223,
-66.6540451049805,-18.4432086944580,
-43.8341674804688,0.0331690311431885,
-11.7835674285889,35.4092063903809,
16.4611072540283,46.8182411193848,
37.9443168640137,25.2872714996338,
44.3745193481445,1.34642803668976,
24.4734134674072,0.0205167233943939,
-14.0826282501221,6.60711860656738,
-51.4024734497070,-2.03857135772705,
-65.2956237792969,-21.8189163208008,
-52.0475082397461,-30.7966060638428,
-22.8428211212158,-11.2408208847046,
5.06290912628174,24.8229789733887,
11.9231815338135,43.6803398132324,
-5.03915786743164,23.1060867309570,
-28.7180652618408,-23.5485630035400,
-33.4988250732422,-48.0140075683594,
-11.6916952133179,-24.4387321472168,
11.4554347991943,24.1711616516113,
12.3924140930176,46.0738258361816,
-3.89540386199951,18.5308570861816,
-7.39554309844971,-25.7649555206299,
15.9657173156738,-39.1428070068359,
40.4456710815430,-22.6519851684570,
35.5694656372070,-11.8666553497314,
1.28872644901276,-23.7482566833496,
-24.6493511199951,-35.6508216857910,
-7.09209823608398,-20.4939804077148,
40.1487121582031,9.09154033660889,
70.2001495361328,22.0439281463623,
50.2614669799805,15.3596200942993,
2.65454387664795,20.6844387054443,
-26.3161201477051,48.2152709960938,
-19.7768802642822,64.2501068115234,
-0.653835594654083,36.6960983276367,
4.37515926361084,-14.1409187316895,
0.0978554785251617,-31.1466865539551,
9.85796737670898,4.18315124511719,
30.2752590179443,43.3087005615234,
40.5710449218750,38.5715675354004,
37.3757400512695,4.06263446807861,
36.9088516235352,-8.92766380310059,
45.6009063720703,17.4957294464111,
44.1275939941406,42.6624488830566,
20.3229408264160,33.3347930908203,
-2.52097773551941,6.82243156433106,
0.403484821319580,2.49104118347168,
17.5434608459473,24.1432285308838,
16.4738044738770,38.6797142028809,
-5.42419052124023,27.0134601593018,
-15.0631847381592,4.85326147079468,
11.0969524383545,-7.19554424285889,
51.0042037963867,-6.06723594665527,
64.3732681274414,-0.886071681976318,
39.5153503417969,7.06734275817871,
-7.85463809967041,14.4071350097656,
-51.8342895507813,7.45337104797363,
-72.8378829956055,-20.9353637695313,
-58.9502029418945,-47.5358238220215,
-27.0925045013428,-43.7657661437988,
-11.5415315628052,-16.2413024902344,
-31.3797206878662,-0.892996609210968,
-54.1006355285645,-15.0429811477661,
-38.3864173889160,-35.8070602416992,
15.5952091217041,-30.5822525024414,
51.3857002258301,-1.32413482666016,
34.1535415649414,23.9320678710938,
-3.64419889450073,23.9599514007568,
-8.26638603210449,12.6272048950195,
21.9534969329834,13.0351982116699,
45.1005706787109,27.6767578125000,
38.9900856018066,35.3965911865234,
23.2120018005371,19.5610599517822,
24.6105842590332,-14.3981304168701,
34.7042121887207,-33.6243476867676,
33.2460365295410,-12.9531478881836,
24.8316688537598,32.5593948364258,
20.6664676666260,62.9698143005371,
8.17725658416748,63.1795234680176,
-33.5199737548828,47.1367607116699,
-86.5707321166992,27.9209022521973,
-99.0872573852539,-0.579429149627686,
-49.8678970336914,-42.0746917724609,
11.2432518005371,-65.6321868896484,
21.2518424987793,-36.6512451171875,
-15.8613777160645,18.3254127502441,
-42.0232124328613,29.5741939544678,
-23.0501785278320,-24.8026733398438,
16.5342044830322,-82.4873504638672,
33.5018043518066,-72.9102935791016,
27.4582252502441,-11.6644134521484,
27.2866554260254,25.3609752655029,
44.9322547912598,2.86429524421692,
57.7726135253906,-29.7772636413574,
47.8900756835938,-21.2207832336426,
25.2221069335938,7.60667181015015,
10.0647869110107,1.39829277992249,
4.33339977264404,-43.8253402709961,
-4.49808216094971,-71.7024612426758,
-17.0767192840576,-43.8975715637207,
-21.7726573944092,9.58846282958984,
-3.74895215034485,30.7779769897461,
22.7117385864258,9.29981231689453,
31.5077419281006,-15.9135990142822,
16.4274692535400,-22.5915813446045,
-2.13941812515259,-29.3835048675537,
-0.995589315891266,-51.1445922851563,
14.2173862457275,-66.7347793579102,
15.4795417785645,-43.7757949829102,
-6.75701951980591,1.45999586582184,
-29.1940937042236,12.8622636795044,
-26.9672660827637,-27.1788978576660,
-6.99042081832886,-63.5444793701172,
9.46778392791748,-41.1820869445801,
10.6778478622437,19.5754547119141,
9.35716342926025,46.6786842346191,
16.3328151702881,14.1342411041260,
23.9019298553467,-32.4826431274414,
22.1328105926514,-38.6178512573242,
10.5940923690796,-17.8761615753174,
-0.734993934631348,-14.9981355667114,
-3.24230504035950,-31.9394931793213,
0.509265959262848,-28.5937900543213,
2.03819966316223,9.52454280853272,
-10.1149606704712,40.3861694335938,
-32.7474441528320,29.1267299652100,
-42.8587303161621,-8.61360836029053,
-20.5607566833496,-26.9583568572998,
22.2262744903564,-16.3878211975098,
46.7598457336426,-10.8816318511963,
27.7126750946045,-27.0336208343506,
-11.3675012588501,-39.4650115966797,
-24.6960144042969,-22.5202407836914,
-0.170328378677368,10.4305553436279,
31.2204074859619,26.2264862060547,
33.0482025146484,16.2978382110596,
0.623302936553955,6.01322221755981,
-38.6235389709473,14.6063842773438,
-57.1790542602539,23.6790866851807,
-50.6389579772949,5.21549463272095,
-29.2173442840576,-31.3897418975830,
-5.20183849334717,-46.2081947326660,
9.31045722961426,-19.8167610168457,
5.85161209106445,23.2116851806641,
-9.16276073455811,46.2126998901367,
-18.5228939056397,45.6219711303711,
-4.32795715332031,42.5646743774414,
25.6827507019043,39.2862968444824,
40.3057022094727,19.5426769256592,
24.5826473236084,-16.6666908264160,
4.28517436981201,-32.5014495849609,
14.7257204055786,-6.85583019256592,
44.3715858459473,27.8998336791992,
48.4514312744141,23.1614151000977,
11.4902133941650,-18.7061138153076,
-20.9422473907471,-44.6137619018555,
-9.43184280395508,-27.3704071044922,
22.7921752929688,2.38013863563538,
20.1616420745850,6.87003898620606,
-16.6615772247314,-4.51248741149902,
-36.3817901611328,-4.67391729354858,
-17.5590934753418,5.97712135314941,
-1.77458000183105,-1.89365053176880,
-18.3599414825439,-32.2396926879883,
-33.1265296936035,-48.8711013793945,
-2.32025337219238,-30.4610939025879,
50.2249145507813,4.98685789108276,
58.3298530578613,28.7116985321045,
13.5935726165771,35.0663642883301,
-27.7997303009033,30.9094448089600,
-27.1998329162598,13.3941516876221,
-12.3950843811035,-12.7462949752808,
-24.1312999725342,-23.6369190216064,
-53.3463859558106,-4.68894100189209,
-59.0079078674316,16.3969364166260,
-37.1053123474121,3.01707530021668,
-21.7799415588379,-42.1670379638672,
-27.4157810211182,-67.4482421875000,
-34.0700683593750,-42.1361236572266,
-23.1535320281982,2.35931634902954,
-0.340327024459839,15.8665819168091,
18.3412151336670,-7.78828620910645,
26.7010021209717,-28.4487953186035,
24.8547058105469,-21.2477378845215,
12.7982606887817,3.74085950851440,
0.424340546131134,20.5501594543457,
2.30339789390564,22.2267570495605,
22.8925514221191,17.2179832458496,
35.1896705627441,17.7550220489502,
13.0411615371704,25.8334751129150,
-23.8376522064209,37.4775352478027,
-31.5128936767578,44.9699134826660,
0.376791477203369,44.5265846252441,
32.9933547973633,33.9844589233398,
29.4728202819824,18.0507335662842,
4.70009040832520,-0.244354113936424,
-5.60318756103516,-22.7359352111816,
8.84652423858643,-39.7342300415039,
24.3694286346436,-37.4549674987793,
26.9964790344238,-24.5465908050537,
29.5044136047363,-23.6351909637451,
42.8946914672852,-33.6098060607910,
50.1588211059570,-23.0006141662598,
33.5162239074707,26.0048217773438,
6.80443191528320,79.6778717041016,
-3.06148576736450,83.9758605957031,
6.24821662902832,39.9127464294434,
10.9633769989014,8.94492626190186,
-3.54217362403870,28.2203865051270,
-31.9119720458984,57.7382049560547,
-53.4120864868164,44.0266189575195,
-54.1552619934082,0.373792529106140,
-33.6809387207031,-10.9158430099487,
-4.56175184249878,21.5381431579590,
5.76431608200073,43.6645355224609,
-18.3524589538574,17.1883201599121,
-55.1891288757324,-16.6236610412598,
-59.5121002197266,-6.83433151245117,
-24.2536277770996,30.8359737396240,
10.1021642684937,34.0087585449219,
9.34173679351807,-10.4282274246216,
-5.58185386657715,-45.9523773193359,
-2.40336084365845,-28.2663822174072,
9.93913841247559,15.5330390930176,
-5.61755275726318,30.4056568145752,
-49.0551872253418,12.4824237823486,
-71.3802108764648,-6.75626850128174,
-40.7692070007324,-9.85804748535156,
8.24182510375977,-8.46029090881348,
27.2608699798584,-16.9452171325684,
19.4172248840332,-32.2983741760254,
19.1904354095459,-42.7737159729004,
30.4427623748779,-42.7159233093262,
27.5065193176270,-26.9080638885498,
6.38106060028076,4.48077964782715,
-1.53225505352020,32.5707664489746,
12.3380517959595,30.2019996643066,
27.2907924652100,4.58159923553467,
26.3145885467529,-3.42356300354004,
21.7405319213867,15.8953790664673,
26.8273677825928,23.7600269317627,
25.9431762695313,-2.70735836029053,
-1.83879971504211,-29.2602462768555,
-32.8220367431641,-7.10265874862671,
-30.4026947021484,49.2998199462891,
-0.222095608711243,70.5083312988281,
16.8963127136230,27.2541351318359,
9.50231456756592,-27.2476749420166,
-0.381575465202332,-40.5994949340820,
-7.15461587905884,-29.6156768798828,
-29.2450981140137,-31.5947589874268,
-57.8775672912598,-36.1772613525391,
-56.7339859008789,-7.54492092132568,
-13.9001674652100,36.7497825622559,
23.0487995147705,40.5952339172363,
12.7354869842529,-4.19760894775391,
-13.3765077590942,-38.1340789794922,
6.48242378234863,-19.5193939208984,
60.6828994750977,13.3320512771606,
76.9151458740234,7.33680534362793,
31.3886318206787,-19.4207038879395,
-17.1997718811035,-8.69765949249268,
-22.7594928741455,38.6148796081543,
-10.6119155883789,60.0033569335938,
-15.9711685180664,27.5145587921143,
-19.0700092315674,-10.1751985549927,
14.9973201751709,-8.99016094207764,
60.6980857849121,7.68819427490234,
61.2828750610352,-8.04803085327148,
17.9326725006104,-46.2893524169922,
-8.60369586944580,-54.6446723937988,
9.20892047882080,-16.1448993682861,
27.8648471832275,27.4273433685303,
8.03907394409180,37.5840606689453,
-19.6249732971191,31.0502147674561,
-12.1218433380127,32.8710479736328,
12.3028135299683,30.2517604827881,
8.76789188385010,4.66014337539673,
-19.5666065216064,-26.7361011505127,
-32.9350852966309,-26.7371807098389,
-11.3299570083618,5.83350086212158,
16.6038074493408,33.3952636718750,
22.4525852203369,33.3174209594727,
17.7538547515869,17.8684921264648,
21.6922569274902,6.85099029541016,
32.0963401794434,-0.895011067390442,
39.0697860717773,-11.0753393173218,
47.2121315002441,-8.30164909362793,
52.8516273498535,21.0510158538818,
31.6064243316650,50.7153587341309,
-18.2623825073242,42.8602294921875,
-54.8044509887695,-0.567888200283051,
-37.8944664001465,-34.2172164916992,
8.83664703369141,-23.9629039764404,
22.7440681457520,11.2609939575195,
-16.0622348785400,29.0410575866699,
-53.6488265991211,8.37906455993652,
-36.2797470092773,-24.3887367248535,
15.6751003265381,-31.0410594940186,
37.9209632873535,-3.71278476715088,
13.6269693374634,30.7125129699707,
-19.2573852539063,41.2160186767578,
-25.4907531738281,22.6105003356934,
-22.1937618255615,-0.565328836441040,
-35.2438507080078,-4.87642574310303,
-55.4789543151856,0.114431500434875,
-52.7739143371582,-10.3827629089355,
-28.4303722381592,-33.4499130249023,
-8.75618076324463,-37.6392211914063,
-7.44113922119141,-16.5929031372070,
-7.70612335205078,-2.01771473884583,
7.81654167175293,-22.2121772766113,
20.0898532867432,-56.3716163635254,
9.15402126312256,-57.5195236206055,
-11.5052623748779,-21.6995754241943,
-4.48556566238403,6.91832256317139,
38.1766548156738,-1.39601469039917,
79.0842514038086,-19.1768760681152,
79.1981811523438,-9.93603515625000,
38.2698860168457,19.8777961730957,
-5.44310283660889,31.1198291778564,
-18.7696380615234,9.58980560302734,
-0.496249437332153,-12.7705125808716,
26.0391998291016,-8.84232330322266,
33.5805740356445,15.7322139739990,
5.63239097595215,34.9310340881348,
-42.9028472900391,26.5763206481934,
-70.9459686279297,-9.96929359436035,
-47.3392028808594,-52.0806808471680,
10.6560220718384,-68.3643569946289,
50.5964202880859,-41.7003326416016,
35.6671867370606,8.05042648315430,
-14.6088781356812,42.0897674560547,
-50.5832214355469,36.5858459472656,
-48.1726760864258,14.1925306320190,
-21.2599372863770,-4.21713638305664,
6.13624572753906,-25.3592510223389,
24.3465480804443,-59.8629951477051,
29.0193386077881,-79.6055297851563,
20.6977920532227,-46.0289077758789,
11.1508798599243,23.9083080291748,
13.4568433761597,67.5697479248047,
22.0822620391846,50.2966308593750,
14.1468839645386,5.89422988891602,
-11.4841480255127,-11.3460721969605,
-24.0266532897949,-2.95935368537903,
-2.24123144149780,-5.28910303115845,
34.8777542114258,-17.3182067871094,
41.5034217834473,-1.54907178878784,
11.8075008392334,50.1525611877441,
-16.7939224243164,89.6924972534180,
-19.8647956848145,82.1363067626953,
-8.94511032104492,45.1560249328613,
-0.132459282875061,11.3347587585449,
6.70869207382202,-15.5403337478638,
16.9891204833984,-47.0476493835449,
19.8909301757813,-57.6696548461914,
9.13080787658691,-21.0669574737549,
2.70121002197266,36.5826492309570,
13.3003578186035,51.5292243957520,
21.6609630584717,9.94382190704346,
2.30392718315125,-27.2244224548340,
-31.8123722076416,-15.8562717437744,
-34.3444137573242,7.84203863143921,
5.64597558975220,-4.43326187133789,
41.8658027648926,-30.8532657623291,
33.7857551574707,-12.1002092361450,
-0.0114340782165527,49.0706253051758,
-15.7554235458374,75.9282455444336,
-2.60995793342590,26.9676494598389,
15.0010881423950,-46.6592330932617,
12.8046026229858,-67.5086364746094,
-8.88406372070313,-33.7751693725586,
-35.9138412475586,-3.56300973892212,
-53.2057914733887,-8.79115104675293,
-45.0488662719727,-22.3212680816650,
-5.01380634307861,-21.9655666351318,
39.4530143737793,-23.0444355010986,
49.9968566894531,-35.7715721130371,
21.7293968200684,-38.6223297119141,
-5.93527412414551,-8.77355384826660,
-2.65652489662170,33.8528938293457,
14.4841527938843,45.8719253540039,
18.3098125457764,14.5121850967407,
14.7315645217896,-21.0018043518066,
21.5535697937012,-17.8314189910889,
34.5564308166504,18.1608428955078,
24.9320087432861,46.8095054626465,
-12.3560533523560,43.2962112426758,
-37.4645233154297,12.0230283737183,
-17.5902862548828,-19.2746887207031,
23.1351833343506,-23.8058662414551,
43.9414024353027,-3.71172547340393,
35.1315383911133,11.5254459381104,
19.6775836944580,7.90748214721680,
10.3424816131592,5.31962633132935,
-2.03736996650696,27.5541267395020,
-16.7387714385986,64.7732696533203,
-21.3946800231934,77.5297470092773,
-19.2344150543213,53.3025550842285,
-31.5463771820068,27.8753166198730,
-59.0476531982422,34.7859382629395,
-64.1308746337891,47.9434509277344,
-19.1754646301270,23.9657783508301,
34.8670272827148,-18.9384727478027,
33.2041969299316,-26.4456310272217,
-23.4209041595459,3.64802956581116,
-64.1054458618164,14.9857959747314,
-39.8286247253418,-24.2023506164551,
14.0402431488037,-56.5321502685547,
36.1953849792481,-19.8527450561523,
15.6274032592773,55.6111640930176,
-9.75615596771240,88.9944610595703,
-17.7228889465332,59.6695709228516,
-19.4987239837647,28.2312221527100,
-22.8544979095459,28.8217391967773,
-13.6264991760254,22.5464363098145,
6.81240749359131,-24.9492969512939,
8.58961105346680,-63.3736877441406,
-15.7312974929810,-37.0116271972656,
-32.7449913024902,26.8956775665283,
-8.11166572570801,42.7002067565918,
34.0366249084473,-11.3801097869873,
49.0393981933594,-68.6682891845703,
28.9631500244141,-67.5623245239258,
1.06823062896729,-22.6785011291504,
-12.6606788635254,17.0132980346680,
-18.1630268096924,34.5627975463867,
-20.7702789306641,44.0972938537598,
-6.32448387145996,39.0882186889648,
26.3885002136230,11.6526832580566,
45.0329475402832,-8.90652656555176,
25.1113662719727,5.84694766998291,
-18.0173339843750,34.7634315490723,
-49.0927162170410,28.3212223052979,
-50.7366218566895,-19.3721313476563,
-28.3862857818604,-55.6620407104492,
9.52180194854736,-42.8249053955078,
44.0080490112305,-5.70424222946167,
44.8279457092285,9.63240432739258,
4.31892204284668,1.90598368644714,
-42.1291084289551,-0.772432625293732,
-45.9452819824219,0.574609994888306,
-7.51479530334473,-20.8108348846436,
16.2638740539551,-52.7195816040039,
-6.84231090545654,-54.1016540527344,
-40.9405555725098,-18.8633594512939,
-37.8588752746582,3.38160324096680,
0.738304138183594,-20.8137416839600,
33.4375190734863,-58.9770469665527,
43.7257270812988,-55.2529830932617,
44.7017135620117,-9.02207660675049,
39.9007835388184,27.4794273376465,
19.0120964050293,21.0405597686768,
-13.4079446792603,-5.40794134140015,
-19.8479881286621,-13.2806053161621,
14.0758161544800,-0.909968852996826,
46.9367637634277,15.1288576126099,
32.2688369750977,24.5657482147217,
-17.3269367218018,26.1548175811768,
-41.0416831970215,15.7759418487549,
-7.84331226348877,-4.70641756057739,
43.8351974487305,-18.6288757324219,
62.4712295532227,-15.2226486206055,
42.3248291015625,2.96503782272339,
10.9127016067505,16.8587722778320,
-10.4113044738770,12.4787425994873,
-26.4773368835449,-5.91894006729126,
-43.2219276428223,-21.9451007843018,
-50.0345840454102,-26.6066379547119,
-41.2420616149902,-12.1886329650879,
-25.8726348876953,18.1356697082520,
-19.1224536895752,38.2534751892090,
-19.4359111785889,30.1979064941406,
-11.6782236099243,11.0181274414063,
5.49177026748657,8.51230430603027,
20.2237968444824,22.9756393432617,
21.8819141387939,17.8652896881104,
4.72172117233276,-22.6414985656738,
-20.1507530212402,-57.8546066284180,
-33.7347335815430,-37.7607994079590,
-29.2069072723389,16.7507476806641,
-16.2503414154053,33.7763595581055,
-9.93493270874023,-10.7196445465088,
-9.59701538085938,-50.5771408081055,
-1.77070975303650,-21.2463436126709,
10.2547922134399,47.2620506286621,
3.48574066162109,70.3035049438477,
-33.5921821594238,22.8504447937012,
-66.1827850341797,-23.4619636535645,
-53.7559509277344,-5.43796157836914,
-9.08615684509277,47.3830299377441,
11.3509998321533,65.4144973754883,
-15.1196098327637,37.8045883178711,
-46.7791938781738,19.4377384185791,
-41.2140541076660,39.8287086486816,
-12.2617254257202,64.1215820312500,
-4.55718994140625,50.3682022094727,
-22.2332935333252,18.7820320129395,
-30.0865173339844,9.69357109069824,
-13.2678165435791,20.1688709259033,
0.736525654792786,13.1496953964233,
-7.51663637161255,-21.7850818634033,
-14.9310827255249,-48.1329956054688,
2.65426874160767,-40.1295928955078,
31.3433284759522,-22.3675251007080,
38.3801612854004,-35.0301094055176,
21.3177814483643,-66.6705627441406,
5.15638637542725,-73.4458312988281,
-2.34204363822937,-39.2697792053223,
-12.3531808853149,1.45093894004822,
-26.2012538909912,10.9965496063232,
-29.2688865661621,-17.5760955810547,
-12.7116718292236,-53.8914756774902,
6.00533580780029,-68.4480361938477,
9.86880588531494,-50.1784400939941,
6.07281684875488,-11.1773719787598,
11.8124132156372,27.3275604248047,
25.6646595001221,45.3805770874023,
34.6904182434082,38.4304504394531,
36.4356040954590,24.9455928802490,
33.3739242553711,20.1681613922119,
15.2118787765503,20.8450794219971,
-22.7387123107910,19.5527534484863,
-60.4329986572266,12.7014350891113,
-70.8435516357422,2.49523305892944,
-48.9618682861328,-14.5417871475220,
-28.0596694946289,-32.2855987548828,
-34.9034423828125,-39.1632194519043,
-55.6474456787109,-27.2003116607666,
-60.9650421142578,-12.1057357788086,
-44.9128456115723,-20.0486850738525,
-24.0442314147949,-42.7949180603027,
-5.80477046966553,-40.6605911254883,
15.1929111480713,1.12317085266113,
27.3866558074951,49.0261497497559,
8.46081256866455,55.4674301147461,
-33.4358329772949,22.3353385925293,
-50.0030097961426,-11.0614452362061,
-9.13709831237793,-19.7300834655762,
54.8523597717285,-14.7028589248657,
75.9221343994141,-11.2960729598999,
36.0817565917969,-1.53841781616211,
-13.6579551696777,20.7118911743164,
-19.7383365631104,36.6234321594238,
7.73535966873169,18.5395278930664,
23.4615097045898,-24.8696556091309,
5.49299907684326,-55.0224876403809,
-22.8156909942627,-46.3325004577637,
-34.8531303405762,-12.1983375549316,
-27.4126853942871,16.8385028839111,
-17.8110046386719,25.8155593872070,
-18.5161800384522,16.6925601959229,
-28.5791530609131,1.13709223270416,
-37.0968780517578,-11.0255889892578,
-33.8201370239258,-23.0279731750488,
-13.3455162048340,-39.1380081176758,
19.3441371917725,-55.3244705200195,
42.0149955749512,-51.6997070312500,
42.2418098449707,-9.10968589782715,
29.5409336090088,55.1180534362793,
16.2245731353760,91.3579864501953,
6.84375810623169,65.6364440917969,
1.44264638423920,4.98032283782959,
1.09533715248108,-30.5747718811035,
2.47484779357910,-23.9713001251221,
-2.30636405944824,-13.4193725585938,
-18.0403461456299,-26.7326049804688,
-26.2041015625000,-45.0284919738770,
-6.62041378021240,-32.2430076599121,
26.7488098144531,6.44916343688965,
30.0837039947510,31.2318286895752,
-12.1294116973877,24.3606281280518,
-58.3940887451172,6.58026266098023,
-61.7783546447754,-5.01854896545410,
-31.5797290802002,-21.9310607910156,
-9.28285884857178,-41.6573791503906,
-6.66633367538452,-38.1634140014648,
-3.20599555969238,0.877261221408844,
11.5016622543335,40.1446723937988,
12.5194244384766,33.9532928466797,
-13.4757452011108,-0.331747770309448,
-41.6615142822266,-11.7802009582520,
-44.8728446960449,12.5194425582886,
-36.4765739440918,30.0037956237793,
-39.4248161315918,8.06127452850342,
-39.1538810729981,-20.4198188781738,
-8.39534568786621,-11.1431293487549,
35.3069267272949,18.7194843292236,
40.8477859497070,17.6636543273926,
1.32360100746155,-18.0130481719971,
-31.8006076812744,-42.5791511535645,
-18.7840080261230,-22.9149169921875,
20.0637989044189,16.7088394165039,
37.4601211547852,35.2671127319336,
27.2054786682129,28.8577976226807,
14.1165266036987,15.7253789901733,
8.05840396881104,2.54153037071228,
-3.36562061309814,-12.4753217697144,
-21.0195159912109,-14.9906711578369,
-23.2628822326660,9.57715892791748,
-5.19173431396484,37.9940109252930,
7.61518812179565,27.2488536834717,
4.00318002700806,-19.6379547119141,
-3.29103302955627,-44.5319099426270,
3.52828526496887,-8.22153663635254,
17.6892738342285,49.8733139038086,
23.8959960937500,62.4796066284180,
15.8113775253296,23.7403030395508,
-1.46483898162842,-10.7771692276001,
-19.2664108276367,-2.94909715652466,
-27.4483451843262,16.9507217407227,
-13.8126802444458,7.91512870788574,
18.3823432922363,-13.5991210937500,
37.0271949768066,-6.09978437423706,
18.4281349182129,33.0580596923828,
-14.0481595993042,53.4974822998047,
-16.1242923736572,29.5961933135986,
22.8023891448975,-1.60658490657806,
59.0314025878906,2.76758241653442,
51.9475593566895,34.1651840209961,
12.2156152725220,41.2558174133301,
-17.7933101654053,3.84094905853272,
-18.1022624969482,-39.4305763244629,
-7.36180400848389,-44.2618293762207,
-7.03237533569336,-18.4106178283691,
-9.19503593444824,-1.15941321849823,
1.92813992500305,0.193081334233284,
16.1507244110107,14.4372177124023,
7.15172863006592,53.4685935974121,
-27.2496528625488,80.6384887695313,
-53.2559356689453,50.6535148620606,
-37.7866477966309,-21.4024047851563,
7.34074687957764,-60.0201606750488,
40.4216995239258,-19.2471332550049,
35.4604110717773,55.1032409667969,
6.20508241653442,86.7241210937500,
-15.2908535003662,57.5758323669434,
-16.1638851165772,16.9411163330078,
-5.04724836349487,3.82467412948608,
5.63849878311157,-5.97498703002930,
5.76554870605469,-44.0120773315430,
-4.53649187088013,-80.4953689575195,
-13.7870292663574,-59.2569808959961,
-4.52098035812378,7.53527927398682,
20.5252342224121,43.6029357910156,
39.2311935424805,12.3202800750732,
32.2392005920410,-34.5981903076172,
7.35298585891724,-33.0182991027832,
-6.90774297714233,0.953099787235260,
-1.55376744270325,-1.66233348846436,
6.32336425781250,-46.8146018981934,
10.4159431457520,-67.8159942626953,
20.8307571411133,-26.1388854980469,
36.8979377746582,37.1774826049805,
40.3468437194824,57.8919448852539,
23.1588745117188,34.7243309020996,
3.12501788139343,22.4126739501953,
-4.17140007019043,43.8729438781738,
-12.8631620407105,64.4485168457031,
-41.1009826660156,43.9184455871582,
-64.1948623657227,-8.40529251098633,
-37.0229721069336,-57.0321922302246,
32.4564018249512,-67.8352050781250,
76.1631851196289,-32.3728256225586,
51.9687843322754,19.9394855499268,
0.654906749725342,43.9583129882813,
-13.3926143646240,23.8988647460938,
11.6475000381470,-6.44243240356445,
28.5092926025391,0.369956731796265,
16.9669742584229,42.6601600646973,
7.49519062042236,68.0537719726563,
18.3136119842529,42.5939826965332,
21.0884857177734,3.47417426109314,
-8.26653385162354,0.0784718692302704,
-40.1006393432617,14.1667785644531,
-28.3188285827637,-3.54787635803223,
13.7810211181641,-47.2471618652344,
29.7362823486328,-58.2526588439941,
0.837424039840698,-14.5365781784058,
-32.2568244934082,31.0919837951660,
-35.6415100097656,27.3524246215820,
-23.3984947204590,-1.94782876968384,
-23.6346263885498,-5.23109197616577,
-35.1747283935547,18.1404190063477,
-35.1914558410645,19.5803298950195,
-18.1254158020020,-15.2807426452637,
1.42763066291809,-43.7693824768066,
16.8452816009522,-37.3242797851563,
31.7881317138672,-16.1689224243164,
35.4133796691895,-10.4575567245483,
12.6658697128296,-11.6929216384888,
-16.3076133728027,-7.92771863937378,
-12.6206007003784,-10.4501581192017,
25.5059719085693,-23.8887901306152,
51.1838417053223,-24.5122280120850,
30.5150203704834,9.02607345581055,
-14.2369384765625,44.0445213317871,
-40.7997093200684,23.4751567840576,
-36.9767608642578,-46.4571075439453,
-23.9244766235352,-85.0022735595703,
-15.1685733795166,-44.5335884094238,
-3.97763538360596,24.2285614013672,
9.58637714385986,44.5919494628906,
12.4012002944946,10.3142004013062,
8.86141014099121,-24.4533786773682,
19.1204357147217,-29.0508975982666,
43.0311088562012,-21.7602863311768,
55.0306549072266,-16.1225719451904,
38.6259269714356,8.67032718658447,
9.36500740051270,60.9746017456055,
-15.5001077651978,95.0301742553711,
-37.8675918579102,70.8820724487305,
-53.3666572570801,14.2566013336182,
-43.9849128723145,-9.45554828643799,
0.451535224914551,11.2088851928711,
50.0288543701172,23.2810363769531,
59.2222671508789,-6.11327791213989,
27.9018363952637,-40.1396827697754,
-3.40889382362366,-33.6515502929688,
-10.4015989303589,6.17798995971680,
-10.0061931610107,29.8003826141357,
-18.3980751037598,16.0385208129883,
-22.9029407501221,-8.06412124633789,
-11.3104419708252,-18.1151504516602,
0.892352759838104,-25.3435802459717,
-2.27102756500244,-44.0680313110352,
-4.72458934783936,-62.1629905700684,
11.0293588638306,-60.2133827209473,
33.6453247070313,-42.7776947021484,
30.4271774291992,-28.2925453186035,
1.32767486572266,-21.2825202941895,
-16.6908073425293,-18.1639385223389,
-1.92025232315063,-13.1295185089111,
19.0420589447022,-10.2966842651367,
16.5000209808350,-12.3192462921143,
-1.61233234405518,-16.0358657836914,
-12.3286323547363,-19.4350738525391,
-13.6569890975952,-25.6788272857666,
-17.9757270812988,-29.0903644561768,
-18.4201011657715,-21.2278614044189,
-3.10960841178894,-13.4800662994385,
14.7417898178101,-19.0982780456543,
5.68849182128906,-28.1872310638428,
-28.7742938995361,-15.7275800704956,
-47.5491180419922,19.2968883514404,
-22.3723583221436,36.3787651062012,
17.3195915222168,7.09958887100220,
23.3784389495850,-42.1679916381836,
-12.4682979583740,-55.9534797668457,
-52.4332008361816,-24.5790748596191,
-62.7677650451660,3.85975098609924,
-38.8888931274414,-3.40688896179199,
4.85984373092651,-18.9536075592041,
45.8398437500000,-0.444292545318604,
55.4689025878906,39.9526557922363,
21.3465385437012,53.5353050231934,
-35.0716857910156,21.4342765808105,
-66.6197814941406,-12.9752988815308,
-50.0844497680664,-11.9793100357056,
-14.6867218017578,11.4867115020752,
-3.35036587715149,18.7909870147705,
-20.5840911865234,1.90994608402252,
-37.7792968750000,-12.1693792343140,
-35.3092041015625,-4.91214752197266,
-26.1907825469971,6.78179311752319,
-20.7087612152100,3.09155678749084,
-13.6674613952637,-8.55159473419190,
-4.42833280563355,-9.52786827087402,
-4.79157733917236,0.513097524642944,
-27.1379890441895,-1.94040238857269,
-49.4176406860352,-30.5116653442383,
-36.5949592590332,-68.5943222045898,
10.5519447326660,-79.8641433715820,
53.8011703491211,-46.0096740722656,
60.4562492370606,4.21473026275635,
40.9432754516602,26.9565429687500,
27.2838706970215,9.37577342987061,
28.7268848419189,-16.7984199523926,
32.4944534301758,-16.9137935638428,
30.3994331359863,9.65402984619141,
30.2310314178467,33.2522048950195,
31.2978343963623,36.3206291198731,
15.4197521209717,27.3055152893066,
-20.3885135650635,13.7699375152588,
-43.8369178771973,-12.6420469284058,
-25.8812751770020,-40.5705604553223,
12.7874279022217,-36.6955451965332,
24.2010955810547,3.13358402252197,
-1.76474118232727,36.7598266601563,
-21.4004688262939,27.9826889038086,
-4.46535587310791,-2.71746635437012,
22.4656963348389,0.124127864837646,
20.1274242401123,32.0029716491699,
-6.62617206573486,33.4077873229981,
-15.5021276473999,-18.1088695526123,
1.47744798660278,-59.0051727294922,
9.27207565307617,-30.9031162261963,
-14.0131731033325,25.7439708709717,
-37.7203102111816,22.3467235565186,
-30.0371456146240,-46.5199851989746,
-0.310748517513275,-84.3730850219727,
13.6255159378052,-28.4919223785400,
2.89487195014954,58.6630897521973,
-7.43331289291382,73.3578491210938,
-0.457064867019653,7.47663068771362,
15.2223300933838,-50.3802070617676,
22.5092639923096,-43.8674163818359,
17.9921360015869,-10.2928428649902,
8.27569484710693,-13.9411239624023,
-2.40893220901489,-47.2368202209473,
-14.8761901855469,-53.9360847473145,
-22.0371723175049,-17.6626205444336,
-19.0993518829346,15.3020334243774,
-14.9055423736572,7.93531990051270,
-20.5575847625732,-19.5936889648438,
-36.9679603576660,-26.8465766906738,
-49.7952575683594,-11.3129549026489,
-36.7017097473145,2.39819979667664,
8.68070888519287,4.85584831237793,
54.6842308044434,14.6954298019409,
58.0027008056641,42.5026245117188,
12.6071481704712,63.9053421020508,
-28.5592155456543,56.7177047729492,
-12.7911071777344,32.2293548583984,
44.0046463012695,13.8631114959717,
70.6598739624023,10.9763031005859,
33.0559959411621,12.9704198837280,
-24.7065086364746,14.2078828811646,
-36.7936477661133,18.6409492492676,
-4.92289972305298,23.1070499420166,
15.5853738784790,7.73115491867065,
1.44171404838562,-32.8503532409668,
-18.3253936767578,-65.7299957275391,
-14.0245008468628,-61.3322181701660,
3.38153266906738,-23.1761722564697,
11.5390548706055,14.0461168289185,
12.9509840011597,17.4001445770264,
22.3767395019531,-12.0929956436157,
25.7041873931885,-46.4098663330078,
9.53046607971191,-52.7957458496094,
-8.16859340667725,-25.9341144561768,
6.19410419464111,12.4472246170044,
48.3276443481445,25.0036067962647,
67.8805236816406,5.73165035247803,
34.1793403625488,-5.42928457260132,
-12.4562339782715,24.2839946746826,
-15.6666021347046,67.6153945922852,
20.4747467041016,61.2329063415527,
43.4170875549316,-9.86147689819336,
22.1246719360352,-77.1092910766602,
-21.5760154724121,-70.1258392333984,
-39.4671936035156,-6.34015178680420,
-16.3942832946777,39.2991638183594,
23.5797939300537,27.6162796020508,
49.7116127014160,-2.34856009483337,
43.2219047546387,1.59269082546234,
10.0356626510620,32.3409233093262,
-22.7700691223145,39.6606216430664,
-27.9460716247559,4.60496711730957,
-8.06032943725586,-41.7569160461426,
3.24496912956238,-59.2027244567871,
-11.2060718536377,-37.4231796264648,
-19.8591403961182,3.35784125328064,
4.28954744338989,34.6447792053223,
36.2374992370606,41.3793678283691,
23.8847827911377,29.1062049865723,
-39.5816802978516,22.1679229736328,
-89.4575195312500,22.8942489624023,
-66.5798797607422,12.4234495162964,
3.47915935516357,-16.6012248992920,
47.8984680175781,-39.5330123901367,
38.9539337158203,-16.0460700988770,
7.14015483856201,47.5413932800293,
-14.4429426193237,90.8251953125000,
-24.5886287689209,69.5008773803711,
-27.5335941314697,11.3794307708740,
-10.8276882171631,-28.4601688385010,
20.6221771240234,-27.6309661865234,
32.6747932434082,-5.39851665496826,
-0.968341886997223,15.3325462341309,
-46.4964752197266,29.8009395599365,
-49.4337310791016,26.8169479370117,
-9.97804069519043,-4.86238622665405,
18.1569824218750,-44.4703788757324,
6.24553966522217,-52.5479202270508,
-13.2443046569824,-15.2487001419067,
-0.916551947593689,27.8128852844238,
19.0224666595459,35.4321594238281,
7.13313674926758,15.7065582275391,
-28.6641540527344,10.1230764389038,
-42.4814300537109,28.7493228912354,
-21.0575523376465,44.5628776550293,
-9.75876808166504,40.5690116882324,
-37.6777839660645,21.7231025695801,
-69.8244628906250,-0.0473346188664436,
-55.3541450500488,-18.2364139556885,
-3.36896657943726,-23.7968006134033,
24.9732055664063,-6.99308490753174,
4.76658439636231,21.7527160644531,
-23.2825450897217,29.5894947052002,
-16.3477077484131,5.47373771667481,
22.5408458709717,-19.1254844665527,
51.6301689147949,-14.3256397247314,
48.7502212524414,3.03265213966370,
26.5914402008057,-8.92504882812500,
7.70451116561890,-49.1012687683106,
-3.12634992599487,-67.2748870849609,
-10.3910989761353,-40.9600753784180,
-15.3694610595703,-1.82010078430176,
-13.5475387573242,9.50278091430664,
1.22091126441956,-2.25945544242859,
24.7827453613281,0.877136707305908,
41.9511566162109,24.9909515380859,
27.8093395233154,37.3095245361328,
-11.6752099990845,15.2294864654541,
-39.1724815368652,-20.9703407287598,
-21.8693695068359,-37.6604118347168,
29.9295272827148,-27.8020858764648,
69.2234725952148,-12.3463163375855,
63.7854003906250,-6.09248733520508,
32.4527206420898,-11.5419397354126,
14.7439994812012,-26.8586959838867,
20.5133514404297,-47.6652488708496,
32.2355918884277,-58.5535850524902,
31.9117908477783,-45.4757575988770,
18.1292324066162,-14.0669612884521,
-5.94130325317383,13.4900083541870,
-35.4784851074219,21.2480831146240,
-54.8876991271973,16.8726692199707,
-44.9275627136231,16.3932571411133,
-9.52771472930908,22.1311111450195,
18.3949527740479,27.4495449066162,
14.2689332962036,29.1837673187256,
-11.0459508895874,25.8233318328857,
-26.9367942810059,7.65787792205811,
-17.5995216369629,-27.7820358276367,
0.527679085731506,-64.5544586181641,
6.02891063690186,-77.3220825195313,
3.36999106407166,-59.0360221862793,
-0.264884918928146,-31.2886085510254,
-1.09886848926544,-20.5710659027100,
-0.672888994216919,-24.1919498443604,
0.949254512786865,-28.9341335296631,
-0.560918688774109,-24.5069484710693,
-7.54650831222534,-18.1201343536377,
-17.7740707397461,-15.2234582901001,
-15.1439781188965,-17.6762123107910,
1.02359318733215,-29.1162948608398,
8.57430171966553,-45.6653976440430,
-12.1491928100586,-46.7206344604492,
-38.0956459045410,-20.7313652038574,
-22.1000232696533,14.5977010726929,
33.0072822570801,20.8398571014404,
67.3583908081055,-9.81964683532715,
38.4319229125977,-38.6794204711914,
-18.3230419158936,-26.7533645629883,
-34.8453025817871,22.1546497344971,
-3.45687842369080,61.7556533813477,
18.2059364318848,68.8155975341797,
-8.02065563201904,51.7020606994629,
-47.7766685485840,21.2365722656250,
-50.8455505371094,-15.3394088745117,
-21.7217826843262,-39.2752609252930,
-4.07147789001465,-30.1236495971680,
-10.6024770736694,7.11635780334473,
-6.98465633392334,35.7203407287598,
24.2934494018555,29.4457073211670,
56.5713500976563,10.0418128967285,
58.5426750183106,6.39252185821533,
33.3148994445801,11.1628522872925,
7.10017013549805,-0.732109785079956,
-1.79194223880768,-17.7368507385254,
6.87291717529297,-1.10615420341492,
18.0191307067871,42.6075096130371,
24.3633441925049,51.1133270263672,
20.1605415344238,-5.34563541412354,
11.8250560760498,-67.4880523681641,
13.7262973785400,-62.2692756652832,
20.2707729339600,5.73504590988159,
8.32880210876465,51.7248268127441,
-28.6291160583496,28.5629634857178,
-52.6065979003906,-19.6534786224365,
-27.5817432403564,-30.0054378509522,
20.6449699401855,-3.77961206436157,
35.9139633178711,10.2784204483032,
7.79860019683838,1.20231330394745,
-12.7355718612671,-1.62933015823364,
11.8982801437378,18.1535034179688,
45.3973617553711,40.0475502014160,
29.6826477050781,42.2152214050293,
-32.3214454650879,30.4164829254150,
-74.7244796752930,16.1395912170410,
-53.4031791687012,-7.55019569396973,
6.39132690429688,-41.3868789672852,
51.2712249755859,-58.5439491271973,
56.4757766723633,-34.1561279296875,
27.8310279846191,12.4597482681274,
-11.7661266326904,34.2691040039063,
-38.3989143371582,28.0397739410400,
-39.0756912231445,27.4232711791992,
-29.0707817077637,44.6929244995117,
-31.1225357055664,46.5946998596191,
-40.2913589477539,10.3244743347168,
-30.7184028625488,-30.8596305847168,
5.74999380111694,-25.9690647125244,
38.2325172424316,15.2749519348145,
35.0897979736328,34.8323097229004,
15.7001609802246,9.86857223510742,
21.9888954162598,-16.6697635650635,
45.3195571899414,-8.01306724548340,
39.0984992980957,14.5918216705322,
-3.95382642745972,13.2360830307007,
-38.2093544006348,-3.91962099075317,
-31.9990730285645,-2.23137116432190,
-9.35083484649658,21.8155994415283,
-6.35036420822144,34.6032791137695,
-8.22600460052490,21.4780788421631,
13.6913166046143,10.9240865707397,
41.4386520385742,24.2039699554443,
24.0663509368897,42.9980087280273,
-35.5734405517578,32.3051567077637,
-69.5143508911133,-1.61954832077026,
-35.2171707153320,-23.4624042510986,
20.3258094787598,-14.2590608596802,
28.5973472595215,14.4462337493896,
-10.5926532745361,44.4220199584961,
-41.1418457031250,58.4636268615723,
-34.0288314819336,41.4988441467285,
-15.3195190429688,-6.38483142852783,
-12.0941143035889,-59.5775032043457,
-14.8826065063477,-78.8130722045898,
-6.20830726623535,-51.1752929687500,
4.83267879486084,-5.82069396972656,
-1.16130065917969,24.6063003540039,
-11.4895439147949,35.0954513549805,
-2.08642292022705,38.0545425415039,
20.8579082489014,37.1404151916504,
19.4693565368652,28.6744155883789,
-15.8098573684692,22.3856678009033,
-50.1960639953613,25.1949806213379,
-51.8666114807129,23.8131561279297,
-23.0411148071289,5.29708862304688,
9.16360473632813,-17.9333972930908,
26.7596740722656,-19.4150791168213,
32.1400375366211,7.87032794952393,
32.2820053100586,32.9279212951660,
23.0311717987061,28.6763381958008,
12.1477222442627,1.72828149795532,
10.2318201065063,-24.6765842437744,
15.9227390289307,-38.0867843627930,
23.7238254547119,-39.4201812744141,
31.3273735046387,-21.1645717620850,
39.0748138427734,12.3858032226563,
35.6485519409180,30.7319755554199,
12.4935760498047,5.71311855316162,
-13.1381721496582,-39.7103195190430,
-13.6982250213623,-45.3774261474609,
8.13938045501709,7.62613630294800,
15.7594461441040,65.0998001098633,
-13.0126953125000,62.1466064453125,
-39.5262031555176,8.39573764801025,
-14.4931707382202,-28.4674434661865,
45.3090667724609,-10.5135593414307,
71.6028671264648,27.4490890502930,
25.1813869476318,32.7528800964356,
-47.7351760864258,7.63719272613525,
-76.6218032836914,-10.3965673446655,
-50.7934799194336,-3.61025738716126,
-14.7180986404419,7.08384275436401,
-2.59220862388611,-4.06951045989990,
-4.14151144027710,-28.3187561035156,
2.48150539398193,-44.0680236816406,
12.2617607116699,-43.2515220642090,
5.06736946105957,-41.6096343994141,
-14.3020429611206,-51.0902366638184,
-19.3489742279053,-54.0618972778320,
-0.112409710884094,-30.5205345153809,
18.7155303955078,13.6353759765625,
7.63909912109375,49.1238975524902,
-29.3713455200195,42.5251007080078,
-57.1560859680176,-1.12958920001984,
-42.2214469909668,-41.9837684631348,
7.89427280426025,-46.1563835144043,
51.7584037780762,-18.2901134490967,
52.0135116577148,13.6165838241577,
12.7733802795410,32.7563629150391,
-27.9455528259277,42.6758918762207,
-33.3384017944336,48.7131462097168,
-4.67691516876221,39.1914978027344,
25.9749927520752,2.25178670883179,
28.5682296752930,-41.4474983215332,
8.14391422271729,-55.2869796752930,
-6.24791336059570,-21.7938861846924,
-1.80717968940735,31.9289016723633,
2.93277883529663,59.7563514709473,
-13.3698482513428,40.9065933227539,
-41.5003356933594,-3.70902609825134,
-41.5069770812988,-35.4443359375000,
5.40735149383545,-38.0508041381836,
62.1306686401367,-19.3856315612793,
72.9030151367188,2.20252370834351,
25.4380798339844,18.1243019104004,
-30.6917743682861,28.6297264099121,
-38.0525512695313,29.5949573516846,
3.74767684936523,12.3850126266480,
39.8765487670898,-16.9559211730957,
28.2580280303955,-31.0899181365967,
-12.0430049896240,-10.7865810394287,
-28.1712265014648,30.3428230285645,
0.341256767511368,56.4758567810059,
42.4400138854981,43.8805389404297,
53.5325393676758,14.9056434631348,
27.1377182006836,9.15985393524170,
0.245900273323059,30.6106719970703,
-1.47448468208313,48.0219230651856,
6.99275875091553,35.3092994689941,
-4.97516536712647,-0.840509474277496,
-31.5295047760010,-30.3789672851563,
-29.7415657043457,-39.1193161010742,
15.4371194839478,-34.6473846435547,
66.8628921508789,-22.4604167938232,
67.2491912841797,1.29206728935242,
17.4654731750488,27.4880714416504,
-24.2029380798340,27.1598548889160,
-15.2679405212402,-5.99425601959229,
19.6679706573486,-37.2171592712402,
26.0295391082764,-26.9235267639160,
-11.2127447128296,12.7589092254639,
-50.5909309387207,23.4871692657471,
-49.5076713562012,-20.0849475860596,
-10.8515262603760,-69.0814056396484,
33.0846176147461,-65.9193420410156,
52.7703399658203,-22.2132549285889,
40.4890747070313,2.19275617599487,
9.00458145141602,-17.2017688751221,
-22.9192333221436,-35.3320350646973,
-41.4252090454102,-12.5893802642822,
-44.8595199584961,21.7466659545898,
-41.5346527099609,17.9618968963623,
-32.2536201477051,-19.0053558349609,
-17.8864784240723,-34.1336898803711,
-2.86662173271179,-4.02794075012207,
-3.96726799011230,25.6631679534912,
-20.7233867645264,7.15898323059082,
-26.8871974945068,-47.2187728881836,
-10.2097511291504,-76.8079528808594,
7.29812860488892,-52.4613647460938,
-0.134490936994553,-5.07082176208496,
-21.4961357116699,22.2388439178467,
-18.9778366088867,19.3952941894531,
16.5148639678955,2.95926904678345,
42.0024490356445,-2.97299861907959,
21.1200714111328,6.35259914398193,
-29.0118522644043,17.0057868957520,
-60.7481994628906,11.9225549697876,
-59.0810661315918,-6.12904262542725,
-45.2987174987793,-21.3183631896973,
-30.3504104614258,-27.1183242797852,
-5.72690820693970,-29.5608234405518,
26.8177051544189,-42.0122413635254,
40.0159835815430,-51.0712318420410,
22.3428955078125,-31.6839828491211,
4.08639574050903,10.8349189758301,
15.8844795227051,34.4297676086426,
41.5192642211914,19.9871692657471,
38.1632881164551,-8.02639770507813,
2.98505377769470,-13.2439966201782,
-20.0615787506104,3.12590837478638,
-3.49183320999146,14.8276958465576,
18.4389915466309,17.4196376800537,
5.02376127243042,27.2508335113525,
-28.8571796417236,38.2409782409668,
-40.0531044006348,16.5960826873779,
-16.4247398376465,-41.7412452697754,
12.6578178405762,-87.8122024536133,
19.3355579376221,-76.2512435913086,
13.5836544036865,-29.3959045410156,
9.73003387451172,-6.59545183181763,
6.40892791748047,-20.8684844970703,
-2.10963082313538,-33.8436927795410,
-7.46479892730713,-20.7311286926270,
-5.41543865203857,-0.453907936811447,
-13.9308414459229,1.46543192863464,
-41.3392562866211,-10.5600194931030,
-56.8299636840820,-23.2469387054443,
-34.4103507995606,-36.8783149719238,
1.87222015857697,-55.4967231750488,
5.68178510665894,-60.9403800964356,
-27.6793422698975,-35.5578689575195,
-50.6126480102539,-3.61624765396118,
-28.5957965850830,-1.58720159530640,
11.7708740234375,-22.6033916473389,
25.6630992889404,-17.8843784332275,
13.6211919784546,22.8005504608154,
0.845016121864319,51.4972419738770,
-11.5988454818726,35.6313018798828,
-33.9477043151856,-4.10374069213867,
-46.2664566040039,-28.9448490142822,
-22.3047790527344,-35.8614997863770,
18.1009654998779,-45.3609733581543,
25.7784652709961,-54.9575233459473,
-4.85190057754517,-39.5116653442383,
-21.0639114379883,-7.10218524932861,
5.63304901123047,5.43213462829590,
34.4789848327637,-4.15225458145142,
12.2311925888062,-6.03166723251343,
-34.7074165344238,3.53566288948059,
-39.0134239196777,-11.7619524002075,
2.83380866050720,-56.4185676574707,
25.8462982177734,-70.7154159545898,
4.70761394500732,-17.2392368316650,
-14.7853136062622,49.3244590759277,
4.83842086791992,51.9821357727051,
30.2630786895752,2.84841322898865,
15.6033735275269,-9.66385555267334,
-15.1658229827881,44.3483505249023,
-10.6719274520874,84.7118453979492,
20.9922809600830,48.4245605468750,
18.2021293640137,-22.6510486602783,
-36.4696502685547,-41.2718238830566,
-79.3240051269531,-7.26383209228516,
-61.0077819824219,8.91792678833008,
-17.9142875671387,-24.8582477569580,
-9.13640880584717,-64.9667587280273,
-27.4539089202881,-68.8067398071289,
-20.1803474426270,-46.2893218994141,
21.5044689178467,-28.5627021789551,
52.8601570129395,-12.3744010925293,
39.2952079772949,14.4071865081787,
0.980945825576782,37.9472961425781,
-21.9804210662842,24.0137100219727,
-22.4649753570557,-22.7725868225098,
-12.1566486358643,-63.8225326538086,
4.05358934402466,-73.3641128540039,
23.7019729614258,-57.2147521972656,
31.0230731964111,-29.0057334899902,
12.9228267669678,-5.03534936904907,
-9.30178070068359,2.52018141746521,
-4.40096426010132,-7.72553396224976,
22.7695903778076,-16.0298175811768,
41.7698783874512,0.727855324745178,
35.1385192871094,36.9515991210938,
20.8295898437500,58.7772865295410,
21.8043899536133,44.7038116455078,
27.2180290222168,23.0572700500488,
10.2419157028198,24.6228446960449,
-32.6052398681641,40.8641433715820,
-68.4347381591797,34.7016372680664,
-66.4779739379883,1.28595483303070,
-26.3207950592041,-23.9079113006592,
22.2744941711426,-16.1972656250000,
48.6678047180176,13.5137929916382,
39.1934394836426,33.2316398620606,
10.0569286346436,34.8594703674316,
-6.59529733657837,32.0799026489258,
1.76050436496735,31.8214035034180,
18.6929664611816,29.0811271667480,
16.8719425201416,26.0821971893311,
-8.24802780151367,32.7833023071289,
-39.9484672546387,44.8168907165527,
-54.4925727844238,44.1799545288086,
-48.6032600402832,25.4621543884277,
-27.6794242858887,12.7918481826782,
-1.94487428665161,23.1005935668945,
13.9821701049805,38.7085456848145,
3.30628395080566,25.1632061004639,
-31.1761493682861,-11.0035114288330,
-57.1435813903809,-25.0471801757813,
-47.1570892333984,4.45678520202637,
-9.07997512817383,41.1799278259277,
23.7269821166992,37.6297607421875,
36.6325912475586,2.87701630592346,
39.8068733215332,-13.4368162155151,
37.0431671142578,11.5547485351563,
15.4943923950195,39.2158088684082,
-26.8508739471436,34.3270339965820,
-62.2342567443848,11.8641157150269,
-61.2780113220215,7.28267145156860,
-31.5973854064941,19.8934822082520,
-8.71570682525635,16.3077583312988,
-3.72902870178223,-14.9842863082886,
2.97937512397766,-36.1681251525879,
21.1465682983398,-15.1171302795410,
35.4755859375000,29.3309516906738,
26.9843692779541,46.8797264099121,
3.70842719078064,23.0377082824707,
-13.0361480712891,-8.96564674377441,
-17.1845798492432,-7.56778287887573,
-17.1746520996094,29.5147953033447,
-16.6187095642090,54.2143440246582,
-7.50888729095459,28.7878265380859,
0.0585557594895363,-30.4340209960938,
-8.14526557922363,-67.8264923095703,
-29.6455383300781,-50.8498420715332,
-38.1619987487793,-2.62088537216187,
-22.5965194702148,20.6650543212891,
-13.0631484985352,2.50195479393005,
-36.6666908264160,-23.0001277923584,
-75.4894256591797,-23.4062442779541,
-77.7430801391602,-10.9954891204834,
-26.6550064086914,-16.2818717956543,
31.8257923126221,-31.9510974884033,
47.4302444458008,-20.5075759887695,
27.0335712432861,25.4762649536133,
17.2768363952637,60.9775314331055,
39.1111717224121,47.5923194885254,
61.8852424621582,5.22612380981445,
55.8109016418457,-11.1273965835571,
31.6798591613770,17.8504905700684,
17.2846755981445,56.2157821655273,
19.1674594879150,55.9949836730957,
20.1389904022217,14.7341585159302,
12.8264074325562,-23.4789237976074,
8.16817855834961,-24.1755104064941,
13.6282176971436,9.19165802001953,
15.0696086883545,38.6548461914063,
2.61739730834961,28.0901260375977,
-15.9367656707764,-15.7137832641602,
-20.1153488159180,-42.5402183532715,
-4.40727424621582,-19.1586055755615,
26.6749858856201,27.8986797332764,
55.0059585571289,38.8833312988281,
57.0006179809570,-0.121128559112549,
24.8445701599121,-33.8073539733887,
-17.1176986694336,-7.56511878967285,
-34.5262336730957,47.7291374206543,
-14.0391883850098,51.6854591369629,
15.6405744552612,-6.04704761505127,
24.4014377593994,-46.6217269897461,
17.9335842132568,-12.9203643798828,
22.5021800994873,49.6091537475586,
36.5033111572266,58.0662918090820,
36.0384750366211,8.92488670349121,
17.3597202301025,-19.4735050201416,
6.19387578964233,12.7351160049438,
7.37067222595215,51.4719963073731,
-2.37423086166382,37.9202041625977,
-30.0538501739502,-5.08978939056397,
-45.6173019409180,-17.5330295562744,
-18.4953765869141,5.26607847213745,
24.1478271484375,8.87271881103516,
32.1321372985840,-28.8549957275391,
3.33600926399231,-64.9407043457031,
-16.0296993255615,-59.1488800048828,
-2.21361875534058,-29.2865142822266,
13.8521709442139,-8.49404716491699,
3.29071593284607,1.03539311885834,
-15.9364728927612,17.6041011810303,
-16.8048000335693,38.5822296142578,
-12.3858041763306,39.2789306640625,
-31.2376842498779,14.6453456878662,
-54.4315567016602,-4.74070167541504,
-39.0627746582031,-1.00502598285675,
18.5992202758789,8.06438541412354,
62.4651679992676,5.31568527221680,
45.1355628967285,-2.79172945022583,
-10.0380640029907,-5.95977258682251,
-40.0563392639160,-0.677882671356201,
-24.0082626342773,11.4310569763184,
6.62968730926514,25.4014415740967,
17.5805950164795,32.1878814697266,
2.29208898544312,21.0253505706787,
-23.4806766510010,-4.29022216796875,
-31.9781475067139,-13.4721851348877,
-8.76106739044190,8.87135505676270,
31.7127628326416,35.9815788269043,
47.1870918273926,31.1879272460938,
12.2261581420898,6.82022094726563,
-38.0433425903320,8.41809368133545,
-42.9397850036621,39.8882675170898,
7.67133808135986,52.0737953186035,
50.4412536621094,14.9339170455933,
29.1599388122559,-28.5270671844482,
-27.7981586456299,-21.9989814758301,
-45.5333938598633,27.9281940460205,
-12.3127441406250,57.7601547241211,
14.9763669967651,37.4914245605469,
-9.53082847595215,3.26043343544006,
-59.1057586669922,-7.62193918228149,
-77.0966567993164,-6.75602102279663,
-44.4336242675781,-21.8556156158447,
5.21446180343628,-43.6482315063477,
35.5192146301270,-37.8996543884277,
34.4708976745606,-4.20938491821289,
2.85005879402161,21.0281276702881,
-42.1323127746582,18.6059989929199,
-69.5760574340820,-1.52141904830933,
-57.0849952697754,-18.6237564086914,
-22.9409503936768,-32.0650634765625,
-8.66147327423096,-45.6594886779785,
-23.1561298370361,-50.4000663757324,
-30.4051113128662,-34.5219688415527,
-13.2743225097656,-7.69302988052368,
-0.176752254366875,6.84474706649780,
-26.5299797058105,0.754386603832245,
-68.1373367309570,-19.1892757415772,
-63.2117271423340,-38.3541526794434,
3.87836837768555,-43.3750991821289,
70.8211975097656,-24.4356174468994,
80.1800460815430,6.16259956359863,
44.4513092041016,14.9619560241699,
17.0222930908203,-16.2023010253906,
16.7841854095459,-61.5713500976563,
15.9618835449219,-73.7935333251953,
-5.89255619049072,-37.6344909667969,
-25.8214893341064,11.0344371795654,
-24.0646915435791,28.1368255615234,
-10.7833757400513,13.5801773071289,
-13.0630865097046,-4.76206016540527,
-27.4083271026611,-8.91723918914795,
-31.5437049865723,-2.39764237403870,
-16.1534576416016,13.8905153274536,
1.13036417961121,33.6653366088867,
3.88158631324768,44.3733863830566,
1.54700493812561,37.8733177185059,
-2.85631847381592,24.9447917938232,
-12.9567108154297,22.4545974731445,
-25.7944774627686,20.7536582946777,
-29.5456199645996,-6.10637807846069,
-11.1454696655273,-50.3408203125000,
19.9017791748047,-61.8075218200684,
40.0791397094727,-13.3199005126953,
37.1824188232422,48.6571998596191,
24.2291660308838,53.6176452636719,
23.2179260253906,3.94559812545776,
38.9254226684570,-24.5978107452393,
57.4047012329102,9.15850925445557,
50.5231704711914,60.1800231933594,
2.09479904174805,60.1589317321777,
-59.4066848754883,16.2366809844971,
-81.0393600463867,-7.94458913803101,
-44.6998443603516,12.9206485748291,
3.98269653320313,36.8216934204102,
11.8883476257324,24.2042598724365,
-19.6356906890869,-0.901028633117676,
-41.8150749206543,3.61271309852600,
-30.2323303222656,28.5226650238037,
-13.5776033401489,27.8787097930908,
-19.4468727111816,-11.1515293121338,
-21.6559333801270,-49.7789726257324,
10.3486995697021,-56.1157493591309,
50.5245056152344,-41.5031433105469,
44.8897056579590,-32.2518081665039,
-4.28115797042847,-35.0432090759277,
-34.5844078063965,-37.5663375854492,
-14.1680202484131,-32.4649810791016,
11.4239311218262,-26.3745365142822,
-11.4267292022705,-18.9712543487549,
-55.0501174926758,-9.75177574157715,
-54.1743469238281,-7.36449718475342,
2.68566560745239,-17.3859176635742,
45.0015792846680,-25.2261886596680,
20.7790451049805,-14.6275529861450,
-33.2075691223145,3.50857734680176,
-46.6741218566895,7.30721759796143,
-8.79189109802246,-9.01955699920654,
34.2018356323242,-27.1201038360596,
47.2732734680176,-28.8901672363281,
39.7578926086426,-14.8022127151489,
32.8526458740234,3.90572261810303,
28.9422454833984,25.2484416961670,
22.0794563293457,40.5060005187988,
14.1031799316406,35.1590881347656,
3.70591402053833,10.6217451095581,
-17.5448970794678,-4.23583412170410,
-46.1351356506348,4.37267875671387,
-57.2558479309082,7.35565185546875,
-31.4103279113770,-24.1107330322266,
5.59466648101807,-69.4843597412109,
21.2541503906250,-81.0139846801758,
20.4266166687012,-55.0081405639648,
27.4216346740723,-31.4887733459473,
41.1419944763184,-35.2521362304688,
34.4401702880859,-36.9127960205078,
1.56253397464752,-7.26158142089844,
-23.6446590423584,27.2513675689697,
-6.98784685134888,20.6774177551270,
31.2357158660889,-10.5892219543457,
49.4665451049805,-15.8066473007202,
37.4763832092285,14.6371603012085,
15.2438058853149,32.5281066894531,
-10.7435369491577,11.9336118698120,
-39.2901458740234,-13.4222354888916,
-55.1745605468750,-9.51152801513672,
-36.3125038146973,0.469884783029556,
0.0727952718734741,-22.8961238861084,
18.0782566070557,-61.3933906555176,
10.2755298614502,-61.6401176452637,
14.8897027969360,-14.2007808685303,
48.2673187255859,21.6520748138428,
66.6009750366211,14.6616983413696,
31.7327117919922,1.63113296031952,
-24.7182407379150,25.3868999481201,
-32.1348152160645,64.7467498779297,
13.7356729507446,69.7607803344727,
40.2812576293945,45.1277847290039,
4.98237991333008,34.2969131469727,
-48.2752685546875,49.7854995727539,
-57.6593780517578,54.7123756408691,
-25.9183197021484,24.0849628448486,
-10.6359491348267,-9.59031009674072,
-37.5938835144043,-10.0616903305054,
-74.7923126220703,6.86690998077393,
-76.7595214843750,-1.54341816902161,
-40.9597091674805,-34.2897071838379,
4.18109512329102,-46.5035896301270,
32.7845764160156,-17.0351581573486,
33.6963043212891,23.6143817901611,
12.1405057907105,34.0611534118652,
-11.0068225860596,6.16582393646240,
-6.11264801025391,-33.6610260009766,
21.2407493591309,-57.2069511413574,
37.5433311462402,-50.6542892456055,
22.2579936981201,-22.8273239135742,
-3.69104480743408,13.4337320327759,
-9.10742950439453,39.4501647949219,
3.76280856132507,46.5597343444824,
3.11755275726318,42.4705924987793,
-19.1520271301270,36.1260643005371,
-34.7309913635254,28.2694797515869,
-24.6949996948242,23.4506454467773,
-11.9189434051514,30.7948760986328,
-12.3835439682007,41.6033096313477,
-9.28884315490723,34.5599746704102,
21.2843418121338,13.8228578567505,
58.4448471069336,8.16342735290527,
51.1798782348633,34.1487998962402,
-4.01277923583984,59.6677055358887,
-50.4758644104004,35.5413208007813,
-41.8645095825195,-25.6331882476807,
-1.90483343601227,-53.9275283813477,
14.9513864517212,-17.5608940124512,
-0.992176711559296,33.0950660705566,
-9.43707370758057,28.4370574951172,
7.52277803421021,-16.5703182220459,
20.2964820861816,-28.9060802459717,
1.34795558452606,16.0231056213379,
-30.3957118988037,53.0095596313477,
-37.2223739624023,23.8991165161133,
-12.5252332687378,-41.0296783447266,
12.8260421752930,-62.4760513305664,
18.4020252227783,-20.9354324340820,
7.92317581176758,23.5274505615234,
-7.36025667190552,15.3381090164185,
-20.1320972442627,-29.8840866088867,
-28.5733394622803,-54.2211837768555,
-21.2896251678467,-33.7089080810547,
-1.39237022399902,3.56863617897034,
7.50241279602051,28.3015747070313,
-6.08387470245361,36.9124603271484,
-25.6180095672607,41.6867332458496,
-25.6731929779053,47.5050506591797,
-2.97075867652893,45.0671348571777,
19.4546527862549,28.0917968750000,
13.0109577178955,5.44479846954346,
-22.2458381652832,-7.65845537185669,
-52.2521858215332,-13.8914375305176,
-44.7217559814453,-22.2531719207764,
0.985440254211426,-37.8481750488281,
44.8478889465332,-49.1936302185059,
39.6697616577148,-30.9153575897217,
-13.8719072341919,19.7131900787354,
-58.8764114379883,61.2449684143066,
-47.3675117492676,48.0635108947754,
0.814372062683106,-10.9974231719971,
23.2530269622803,-58.6335220336914,
-0.781584501266480,-46.9068679809570,
-22.4968986511230,3.54434967041016,
-2.08946561813355,34.6761627197266,
35.5403327941895,30.1845893859863,
35.8524246215820,24.3677387237549,
-7.06651973724365,45.4247741699219,
-39.6663894653320,64.1984100341797,
-24.0613174438477,45.3911209106445,
8.06074428558350,6.85869359970093,
10.2578973770142,-4.38661766052246,
-14.2168426513672,15.4599037170410,
-25.2060546875000,26.6299686431885,
-1.81837654113770,6.65269422531128,
36.5121955871582,-13.5650196075439,
61.3338508605957,-0.277708530426025,
51.7114562988281,27.2091007232666,
4.84289407730103,31.2571220397949,
-55.7097167968750,11.0458354949951,
-81.7584304809570,-3.80373334884644,
-45.1300201416016,-9.11264991760254,
11.9138088226318,-27.2894115447998,
18.0001144409180,-52.4137191772461,
-33.3287811279297,-46.5123405456543,
-67.2063217163086,-6.53262710571289,
-26.1453208923340,18.8790893554688,
41.2477340698242,-0.0504510402679443,
51.2044258117676,-27.3034553527832,
5.68957996368408,-9.15103244781494,
-15.3063287734985,38.6498489379883,
20.0006237030029,51.8117790222168,
49.5665550231934,12.9385404586792,
12.0580482482910,-23.8742427825928,
-63.0602149963379,-19.0153102874756,
-85.9484558105469,-1.52687156200409,
-29.3965873718262,-11.9845237731934,
46.6123657226563,-34.3954315185547,
70.1707916259766,-32.9161376953125,
29.5614147186279,-13.2851915359497,
-32.6321716308594,-11.2162170410156,
-64.5815887451172,-30.1232738494873,
-44.9874114990234,-31.9302043914795,
4.63156366348267,-0.614615678787231,
24.8396339416504,28.4906826019287,
-9.09918594360352,23.6186370849609,
-47.3839607238770,3.29884815216064,
-26.6588935852051,-1.92108678817749,
46.2525520324707,2.64291357994080,
95.3600616455078,1.62884712219238,
67.0818862915039,9.81633472442627,
0.424278497695923,41.4491271972656,
-30.5311870574951,68.5837707519531,
-15.4431152343750,52.0150032043457,
-8.35664367675781,3.35899424552918,
-29.4742317199707,-16.9402160644531,
-51.9583168029785,11.3978023529053,
-58.4301376342773,33.5830688476563,
-61.7168884277344,-0.364551305770874,
-67.3072357177734,-52.2017440795898,
-46.1654548645020,-50.1777763366699,
7.71780776977539,0.127034664154053,
42.5375938415527,28.6629829406738,
14.2742424011230,4.57423686981201,
-48.1036720275879,-25.4377899169922,
-72.9616622924805,-17.7979564666748,
-44.0363082885742,2.93753671646118,
-19.5627670288086,-7.76694059371948,
-38.4251785278320,-40.3595161437988,
-58.9957847595215,-47.8122215270996,
-35.8077888488770,-22.3733596801758,
11.9221572875977,1.57960641384125,
32.2089424133301,-0.250880241394043,
12.4000787734985,-6.17386627197266,
-14.9166460037231,1.38267111778259,
-25.5199794769287,4.06091499328613,
-24.9739418029785,-15.3304595947266,
-14.4659423828125,-38.9687881469727,
18.0747871398926,-42.9519424438477,
59.1281356811523,-27.3261299133301,
62.6565628051758,-10.5228700637817,
9.90793037414551,-2.16755867004395,
-47.2103309631348,1.77950835227966,
-44.8830604553223,7.81443309783936,
5.81410169601440,15.3769178390503,
35.9684486389160,25.5618133544922,
7.97187089920044,39.2837028503418,
-42.0057563781738,43.3045272827148,
-63.1459884643555,26.8381366729736,
-49.6563835144043,7.10041570663452,
-36.3923301696777,9.25691986083984,
-42.3743019104004,24.5930347442627,
-51.7537269592285,20.5657501220703,
-51.8434829711914,-14.0401134490967,
-50.7690887451172,-45.0165596008301,
-50.3564720153809,-46.5398674011231,
-41.2390670776367,-32.6240348815918,
-16.6931247711182,-31.4803504943848,
10.8452806472778,-39.0661468505859,
28.3957405090332,-24.5066509246826,
34.0422744750977,19.0434360504150,
29.3496303558350,53.8876647949219,
13.6966314315796,51.7849235534668,
-9.92716407775879,26.7971858978272,
-30.3274555206299,4.69479131698608,
-34.9527816772461,-7.29196262359619,
-30.5740108489990,-19.3940620422363,
-33.3679885864258,-31.4920692443848,
-32.3355979919434,-40.7728004455566,
-7.49210166931152,-55.4895324707031,
32.5218162536621,-74.3054962158203,
49.6423683166504,-71.4801635742188,
28.3457641601563,-26.2031497955322,
-5.99806833267212,33.0627098083496,
-19.8429870605469,45.7831764221191,
-11.6937799453735,-5.86113643646240,
-3.87619900703430,-65.2339935302734,
5.05203866958618,-64.5231094360352,
29.2249908447266,-9.58906459808350,
50.5589179992676,36.4524726867676,
33.6287307739258,38.3643302917481,
-14.5213356018066,7.81279468536377,
-34.8758621215820,-19.0171356201172,
3.92762088775635,-21.6037845611572,
49.8767356872559,-1.49676775932312,
38.1825523376465,28.9954223632813,
-16.0966606140137,45.3208999633789,
-37.1525955200195,33.0493087768555,
1.59091401100159,6.97088003158569,
37.1800880432129,4.59916353225708,
12.5246229171753,26.9097385406494,
-47.2599563598633,34.2304420471191,
-69.8825683593750,-0.902631759643555,
-38.3980255126953,-32.5812911987305,
0.648930788040161,-4.54759025573731,
9.56220436096191,60.1879997253418,
-1.73436617851257,86.4555435180664,
-6.45793294906616,37.0401229858398,
-1.66755998134613,-34.3622016906738,
10.8137531280518,-54.1176338195801,
29.2217063903809,-19.5865192413330,
46.0718154907227,17.2341175079346,
41.8642311096191,28.9847297668457,
6.37647485733032,27.6532325744629,
-38.2634506225586,25.3746051788330,
-57.8973770141602,15.0436353683472,
-47.4429168701172,3.10475325584412,
-28.9470977783203,16.1531696319580,
-13.9571723937988,51.9941825866699,
0.915872097015381,63.5121803283691,
9.90536117553711,19.1443004608154,
9.03884792327881,-49.6270828247070,
7.51217460632324,-77.5069885253906,
25.4171657562256,-47.0907859802246,
56.4703369140625,-4.93431472778320,
68.2328033447266,2.96861386299133,
47.8165016174316,-16.5538406372070,
23.5279846191406,-27.2473506927490,
30.6607093811035,-17.5902996063232,
53.6104469299316,2.20358753204346,
51.8794174194336,23.6910934448242,
17.2310104370117,40.1490402221680,
-10.1446084976196,40.3907546997070,
-0.446153044700623,17.8968715667725,
22.7517871856689,-6.14678287506104,
25.9741783142090,-0.0302776694297791,
2.79848003387451,35.9202308654785,
-23.4957351684570,62.1662254333496,
-37.5664634704590,41.5963211059570,
-38.3809509277344,-15.8920869827271,
-21.7248649597168,-63.4952316284180,
13.8399095535278,-74.6627502441406,
54.9244384765625,-52.1227302551270,
74.5519332885742,-14.4764347076416,
59.3895835876465,19.3336238861084,
30.8191566467285,32.8826293945313,
12.7545318603516,26.4842319488525,
9.89733409881592,13.2371168136597,
15.5167417526245,7.95414113998413,
28.2515907287598,11.7458648681641,
42.2829055786133,9.45347499847412,
44.6583480834961,3.94277715682983,
32.0474052429199,14.8785209655762,
14.8621139526367,40.3549804687500,
-1.29740476608276,45.7119102478027,
-21.1716442108154,10.3598213195801,
-50.8304901123047,-28.5891075134277,
-70.1804656982422,-22.4354362487793,
-52.9894714355469,14.9003391265869,
-10.2911024093628,20.8654670715332,
12.0688276290894,-28.8652305603027,
-6.21953821182251,-70.4201278686523,
-30.8549537658691,-42.6669502258301,
-29.7856979370117,25.5160751342773,
-10.7401180267334,48.7464561462402,
1.09752869606018,2.51328325271606,
8.51966667175293,-43.0291213989258,
28.1501522064209,-25.1176471710205,
43.3120117187500,29.3036918640137,
16.5947933197022,52.0934677124023,
-40.1509857177734,26.0508594512939,
-64.8919296264648,-9.47779273986816,
-24.3497581481934,-17.4728832244873,
32.3153800964356,-5.49992227554321,
34.3308105468750,4.46234416961670,
-14.2806634902954,2.58639287948608,
-42.0208702087402,-9.77432441711426,
-19.0390548706055,-31.2771739959717,
14.5204124450684,-48.7853546142578,
10.8027572631836,-41.1685676574707,
-22.1027622222900,-8.33731365203857,
-40.6267166137695,16.1293392181397,
-23.8095092773438,16.5101165771484,
5.77843284606934,16.1829566955566,
19.0513858795166,33.0848464965820,
8.95492935180664,43.2443695068359,
-8.60957241058350,13.8657484054565,
-9.42651081085205,-39.2886924743652,
14.1275215148926,-57.0593605041504,
44.8130035400391,-16.9630279541016,
46.9410095214844,25.4646244049072,
4.31888771057129,17.5335636138916,
-43.7432746887207,-17.9946498870850,
-52.1052131652832,-25.9472675323486,
-22.4436416625977,1.29180324077606,
6.03300714492798,14.0784091949463,
6.91764354705811,-15.3546028137207,
-7.42971992492676,-41.5004730224609,
-8.94575595855713,-21.9817161560059,
8.48079109191895,22.6234054565430,
28.7369480133057,40.0859680175781,
40.6441802978516,21.4519138336182,
35.9857673645020,8.62810230255127,
7.79217433929443,25.3408660888672,
-31.2689838409424,35.9207496643066,
-44.5715446472168,3.96569204330444,
-12.2261543273926,-41.4214897155762,
33.8285560607910,-37.7240562438965,
41.4723930358887,24.1752815246582,
3.73464465141296,80.1425476074219,
-25.2772884368897,62.9749107360840,
-3.94098043441772,-19.9546527862549,
39.9990158081055,-88.5934066772461,
44.5122947692871,-76.1828613281250,
1.21797871589661,-8.19653320312500,
-35.0148811340332,34.2881469726563,
-22.7670612335205,7.22426605224609,
10.0002574920654,-47.4928588867188,
17.0008869171143,-56.4282073974609,
2.00536394119263,-6.61438417434692,
1.84253025054932,42.4796791076660,
23.6683082580566,36.5984191894531,
27.0499134063721,-4.35085391998291,
-6.94693660736084,-26.2121658325195,
-35.2773361206055,-18.1626834869385,
-13.7033882141113,-10.2844791412354,
35.5997734069824,-11.0143728256226,
52.4417648315430,3.16016101837158,
20.6857872009277,42.7607803344727,
-16.9579181671143,74.0645446777344,
-26.6530818939209,65.9335327148438,
-21.6162414550781,36.6513023376465,
-24.8918819427490,16.3663921356201,
-25.0719871520996,1.38516366481781,
-7.39738082885742,-31.3679428100586,
10.8974885940552,-66.1548309326172,
4.30667304992676,-59.2330818176270,
-15.3826818466187,-8.06166648864746,
-13.7807874679565,31.7850914001465,
11.1413335800171,25.3180580139160,
18.9727268218994,1.89222252368927,
-6.69890785217285,4.24002695083618,
-27.3744640350342,19.2991485595703,
-8.27128028869629,6.42411994934082,
27.7249469757080,-26.9573993682861,
30.3228626251221,-31.8021812438965,
-17.5078315734863,6.61608886718750,
-71.6987152099609,34.7028694152832,
-79.1436538696289,7.30472135543823,
-33.3371734619141,-40.3830299377441,
20.5958843231201,-44.0839576721191,
33.6002731323242,-0.116452753543854,
-2.01301765441895,27.6691093444824,
-45.6634292602539,1.15824794769287,
-46.4444541931152,-37.7513847351074,
0.539086818695068,-32.5775184631348,
45.5319862365723,15.8384494781494,
38.4606971740723,51.2458190917969,
-8.54495811462402,35.8430252075195,
-37.9372787475586,-8.71928596496582,
-21.1704978942871,-40.7285537719727,
14.8536520004272,-50.3235054016113,
31.4958419799805,-53.9902458190918,
25.6407184600830,-54.8256378173828,
24.9228935241699,-41.8387756347656,
40.0530319213867,-10.1149187088013,
46.0908164978027,23.3355808258057,
29.9294872283936,32.0166549682617,
2.78028225898743,9.99863910675049,
-13.9747447967529,-15.8046388626099,
-14.1601181030273,-17.1899986267090,
-3.82883310317993,3.04530572891235,
10.4183263778687,18.5046920776367,
24.4825935363770,13.8211927413940,
22.8024215698242,0.811300694942474,
-1.67135882377625,5.70478010177612,
-27.6569633483887,27.0584449768066,
-25.6436405181885,27.7217674255371,
3.33986330032349,-5.88566923141480,
27.8572139739990,-40.3661079406738,
14.5530872344971,-37.3434944152832,
-22.1999778747559,-5.45751190185547,
-45.5954780578613,12.7730684280396,
-38.7937469482422,-0.943095266819000,
-20.2675209045410,-13.7447729110718,
-13.8044471740723,4.97103929519653,
-25.0348758697510,26.7265243530273,
-38.8689422607422,8.30001926422119,
-35.5020446777344,-42.6463546752930,
-7.96148061752319,-71.7551956176758,
31.3779640197754,-54.9695701599121,
55.7330780029297,-31.0827655792236,
49.2880973815918,-42.0857315063477,
29.2088184356689,-66.4098434448242,
31.9642429351807,-52.8314590454102,
63.8003654479981,-1.34493494033813,
89.1152725219727,33.5285224914551,
69.1623153686523,15.8580827713013,
15.5148992538452,-21.8777847290039,
-22.1206378936768,-23.9798469543457,
-22.1746425628662,15.4434719085693,
-4.72972631454468,51.2271308898926,
0.386892884969711,49.8501014709473,
-6.72440528869629,27.1812229156494,
-8.86604404449463,15.5868606567383,
-3.75962901115418,17.7688560485840,
-2.82030701637268,13.1512861251831,
-5.10542726516724,-12.1275758743286,
3.50430440902710,-46.5725860595703,
25.7911491394043,-54.8065872192383,
45.3768234252930,-24.8237762451172,
47.4816436767578,25.4204730987549,
35.6863670349121,54.4015579223633,
16.8227825164795,42.7251167297363,
-5.18884658813477,5.67910671234131,
-27.5725593566895,-20.6856594085693,
-33.2420272827148,-23.2987518310547,
-16.3531284332275,-19.6176376342773,
8.83024978637695,-19.0236968994141,
20.4376697540283,-7.77090597152710,
20.9673900604248,20.6009769439697,
26.4345912933350,41.9060897827148,
35.7484054565430,23.0487937927246,
26.3832855224609,-25.2925243377686,
-7.46172237396240,-49.1652259826660,
-35.2164688110352,-16.3952598571777,
-21.8235263824463,41.7244529724121,
19.6822643280029,67.1146316528320,
39.3091583251953,45.4728088378906,
14.2462863922119,14.9582843780518,
-28.7616691589355,11.9980459213257,
-41.7132301330566,29.0598144531250,
-16.7918643951416,30.5444316864014,
7.45704174041748,6.50444030761719,
-0.277896881103516,-17.8081417083740,
-28.4813365936279,-19.2715053558350,
-37.9751091003418,-4.15793704986572,
-16.3464469909668,2.61948704719543,
9.34628868103027,-13.3053388595581,
4.14025592803955,-34.0361328125000,
-26.4858551025391,-34.8431015014648,
-47.5479278564453,-12.1359519958496,
-35.1859855651856,14.9447364807129,
-13.3338041305542,25.1451072692871,
-17.4307689666748,11.3216991424561,
-44.9926223754883,-12.6346683502197,
-57.0357513427734,-28.0340118408203,
-28.6465778350830,-27.5603542327881,
20.2287387847900,-11.3055000305176,
48.1026535034180,12.7321052551270,
40.8148651123047,34.1594238281250,
24.8997249603272,36.1397781372070,
21.6496868133545,10.8077554702759,
25.9054794311523,-36.0562171936035,
23.1371974945068,-72.5088119506836,
17.0119857788086,-68.6730575561523,
24.9075241088867,-26.7773933410645,
48.1544952392578,14.7552928924561,
62.4356307983398,18.5378208160400,
46.5456199645996,-13.7491569519043,
12.0931491851807,-42.2142829895020,
-15.7817707061768,-37.4943885803223,
-21.1687164306641,-9.84360980987549,
-10.8659162521362,10.9655227661133,
-0.378482401371002,8.64523983001709,
6.17681789398193,-6.87189722061157,
16.2316589355469,-22.0025329589844,
26.8737926483154,-35.8628425598145,
32.4516487121582,-48.7199974060059,
27.6649303436279,-54.9281921386719,
15.7124872207642,-46.4229354858398,
9.25314998626709,-22.2920646667480,
13.1331777572632,4.43368148803711,
15.9734792709351,21.8638038635254,
2.42282915115356,15.1383428573608,
-25.2424736022949,-8.28179168701172,
-36.9958457946777,-22.8654174804688,
-8.32366275787354,-12.3925638198853,
45.1907615661621,13.8618335723877,
73.4424133300781,25.7459278106689,
48.7458038330078,4.70826721191406,
6.37867927551270,-23.2980308532715,
5.62954521179199,-25.8153057098389,
50.8708305358887,-4.29535675048828,
86.4223098754883,15.7599802017212,
65.7485046386719,21.5912094116211,
8.56275653839111,22.6505508422852,
-29.0975589752197,15.6255970001221,
-24.6389961242676,-17.7277317047119,
-2.35231399536133,-64.9542388916016,
6.16663408279419,-74.0734863281250,
-1.36383819580078,-13.5034523010254,
-14.9487085342407,63.3532714843750,
-31.9987220764160,72.3575134277344,
-40.9542655944824,2.92973232269287,
-26.3146114349365,-65.5822601318359,
5.79441165924072,-58.9538192749023,
20.0805530548096,0.278109550476074,
-6.72291183471680,37.0049133300781,
-44.2960472106934,21.5103778839111,
-48.6753692626953,-17.0928783416748,
-15.9066429138184,-43.9273109436035,
13.6439609527588,-49.7992401123047,
21.7842578887939,-39.5296478271484,
28.7857074737549,-14.5345325469971,
52.4029769897461,19.0689163208008,
55.7918052673340,43.3526496887207,
10.9125919342041,49.7928733825684,
-48.0855903625488,40.4519882202148,
-59.4187355041504,17.5147533416748,
-18.9945583343506,-23.9134941101074,
15.4242897033691,-64.7585067749023,
5.51620244979858,-62.2304229736328,
-17.0197849273682,-8.19867610931397,
-12.1989622116089,43.0286178588867,
4.97525119781494,43.4495468139648,
-5.52955055236816,9.65311622619629,
-36.0874748229981,-5.27777814865112,
-41.4335136413574,12.7946186065674,
-15.4165477752686,25.4963665008545,
-8.33368206024170,6.53328561782837,
-42.3357772827148,-18.7013397216797,
-73.6946945190430,-18.3184528350830,
-55.3094367980957,-2.77511477470398,
-9.95658779144287,-2.63223242759705,
10.1763715744019,-16.1909847259522,
-6.21298027038574,-25.7981681823730,
-19.3386859893799,-28.9543151855469,
-3.82560205459595,-37.1974067687988,
12.0388736724854,-38.9195632934570,
1.02586698532105,-15.0146112442017,
-20.3290882110596,20.9834022521973,
-27.1417713165283,41.2898330688477,
-24.7059955596924,41.2060661315918,
-26.1888103485107,39.7597160339356,
-22.4973430633545,42.4778099060059,
-1.44607329368591,24.2844944000244,
21.9341106414795,-21.3304519653320,
30.3701477050781,-52.7983398437500,
33.4203033447266,-36.2097167968750,
55.3851585388184,1.93645298480988,
81.6165542602539,15.8233270645142,
65.9775161743164,10.3284368515015,
4.94718742370606,25.8709945678711,
-39.3222999572754,58.5889968872070,
-21.8662757873535,58.4535903930664,
21.7342777252197,8.59586906433106,
30.0829696655273,-39.9235992431641,
1.67666554450989,-33.0700492858887,
-13.5007572174072,14.6967287063599,
1.75709080696106,47.1134033203125,
12.1865100860596,43.8757095336914,
-3.12602066993713,35.5753898620606,
-11.4995756149292,41.8726196289063,
16.2895259857178,46.2286872863770};
