shortreal out[16384] =
'{0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1.55259199880918e-20,
2.71896480054319e-18,
1.05968205758760e-17,
3.24844679159211e-17,
7.62368496930436e-17,
1.60939026070285e-16,
3.02105523824797e-16,
5.18451979294971e-16,
8.18835114561086e-16,
1.18704764239170e-15,
1.58760084106055e-15,
1.90037156848246e-15,
1.97310205249845e-15,
1.46530781232275e-15,
-9.13225925104264e-18,
-3.18958387804900e-15,
-8.89092961173276e-15,
-1.82538107350826e-14,
-3.24263151865647e-14,
-5.29805962556224e-14,
-8.14227903308228e-14,
-1.19759115276528e-13,
-1.69548606382929e-13,
-2.32887222961081e-13,
-3.11916697982514e-13,
-4.09560325107319e-13,
-5.28508606236627e-13,
-6.71499314486290e-13,
-8.41473483774446e-13,
-1.03967355558066e-12,
-1.26806161057647e-12,
-1.52450773359403e-12,
-1.80777300681084e-12,
-2.11307685758777e-12,
-2.43611467803939e-12,
-2.76724888663427e-12,
-3.09613923041296e-12,
-3.40490548082772e-12,
-3.67242000698376e-12,
-3.86222217402255e-12,
-3.93343300639226e-12,
-3.95642936815155e-12,
-3.98897971945478e-12,
-3.99569830347724e-12,
-3.91344118569337e-12,
-3.68341598541710e-12,
-3.30984783851462e-12,
-2.85132334409965e-12,
-2.55468194342023e-12,
-2.79943234392233e-12,
-3.92436820886855e-12,
-6.28247020378892e-12,
-1.02393744524920e-11,
-1.61266052595144e-11,
-2.42408992184862e-11,
-3.47007561574131e-11,
-4.76429243279064e-11,
-6.34322733228387e-11,
-8.22911322417852e-11,
-1.04399926204035e-10,
-1.29974891960316e-10,
-1.59255469922570e-10,
-1.92513852081966e-10,
-2.29986377164870e-10,
-2.72038613857717e-10,
-3.18953891076390e-10,
-3.71116554154227e-10,
-4.28971885790830e-10,
-4.92793972295402e-10,
-5.62817181748443e-10,
-6.39252262235601e-10,
-7.22271298325694e-10,
-8.11874234507570e-10,
-9.08225050721967e-10,
-1.01161423682328e-09,
-1.12223108583720e-09,
-1.24042298654814e-09,
-1.36666400418761e-09,
-1.50136181265026e-09,
-1.64474411867843e-09,
-1.79702830394035e-09,
-1.95838345540267e-09,
-2.12894080142689e-09,
-2.30897767572458e-09,
-2.49862952550473e-09,
-2.69793898333148e-09,
-2.90698176641513e-09,
-3.12572190352967e-09,
-3.35412164709226e-09,
-3.59222585011310e-09,
-3.84000653497196e-09,
-4.09745304352782e-09,
-4.36474589804448e-09,
-4.64215688111835e-09,
-4.93011942381827e-09,
-5.22925835966248e-09,
-5.54041124090077e-09,
-5.86454840245665e-09,
-6.20256024319588e-09,
-6.55529186488479e-09,
-6.92362389642653e-09,
-7.30850668873018e-09,
-7.71096075879996e-09,
-8.13225309315158e-09,
-8.57362092432368e-09,
-9.03633345927801e-09,
-9.52186951508338e-09,
-1.00315089568426e-08,
-1.05665831640067e-08,
-1.11285398673999e-08,
-1.17189431492193e-08,
-1.23394201523297e-08,
-1.29915385116419e-08,
-1.36770559322486e-08,
-1.43976830457859e-08,
-1.51549688354180e-08,
-1.59504320862425e-08,
-1.67856235577801e-08,
-1.76622894088041e-08,
-1.85822184306517e-08,
-1.95470573061129e-08,
-2.05585699575295e-08,
-2.16185878088027e-08,
-2.27288392551372e-08,
-2.38910651262358e-08,
-2.51071323731367e-08,
-2.63790198573588e-08,
-2.77086371625046e-08,
-2.90980217698689e-08,
-3.05491880681075e-08,
-3.20640722861754e-08,
-3.36448096049935e-08,
-3.52934321767862e-08,
-3.70121071568974e-08,
-3.88030976239406e-08,
-4.06685352061231e-08,
-4.26106048223573e-08,
-4.46313599411496e-08,
-4.67328362674380e-08,
-4.89173288542588e-08,
-5.11871469655034e-08,
-5.35446140759177e-08,
-5.59921673470853e-08,
-5.85320982793292e-08,
-6.11667729799592e-08,
-6.38986961121191e-08,
-6.67304576040806e-08,
-6.96647646236670e-08,
-7.27043101278468e-08,
-7.58518012844434e-08,
-7.91099452612798e-08,
-8.24815344913077e-08,
-8.59695035160257e-08,
-8.95766305575307e-08,
-9.33058572627488e-08,
-9.71602318600162e-08,
-1.01142745734251e-07,
-1.05256596327763e-07,
-1.09504860290599e-07,
-1.13890592956523e-07,
-1.18416899397289e-07,
-1.23086721259824e-07,
-1.27902964663917e-07,
-1.32868819946452e-07,
-1.37987484549740e-07,
-1.43262056440108e-07,
-1.48695903590124e-07,
-1.54292351339791e-07,
-1.60054895559369e-07,
-1.65987046329974e-07,
-1.72092285311010e-07,
-1.78374250481284e-07,
-1.84836807193278e-07,
-1.91483763956057e-07,
-1.98318915067830e-07,
-2.05346168513643e-07,
-2.12569261748286e-07,
-2.19991818539711e-07,
-2.27617533710145e-07,
-2.35450201557796e-07,
-2.43493673224293e-07,
-2.51751856694682e-07,
-2.60228716797428e-07,
-2.68928175728433e-07,
-2.77854184105308e-07,
-2.87010692545664e-07,
-2.96401623245401e-07,
-3.06030869978713e-07,
-3.15902298098081e-07,
-3.26019744534278e-07,
-3.36387188326626e-07,
-3.47008693779571e-07,
-3.57888438884402e-07,
-3.69030715319241e-07,
-3.80439814762212e-07,
-3.92120000469731e-07,
-4.04075848337016e-07,
-4.16311905837574e-07,
-4.28832663601497e-07,
-4.41642583837165e-07,
-4.54746071909540e-07,
-4.68147817400677e-07,
-4.81852509892633e-07,
-4.95864981076011e-07,
-5.10190261593380e-07,
-5.24833410509018e-07,
-5.39799032139854e-07,
-5.55092128706747e-07,
-5.70717645587138e-07,
-5.86680357628211e-07,
-6.02985380737664e-07,
-6.19637717136357e-07,
-6.36642539575405e-07,
-6.54004793432250e-07,
-6.71729651458008e-07,
-6.89822229560377e-07,
-7.08287757333892e-07,
-7.27131521216506e-07,
-7.46358978176431e-07,
-7.65975698868715e-07,
-7.85987197104987e-07,
-8.06399214070552e-07,
-8.27217320420459e-07,
-8.48447029966337e-07,
-8.70094368110586e-07,
-8.92165189725347e-07,
-9.14665349682764e-07,
-9.37600702854979e-07,
-9.60977104114136e-07,
-9.84800635706051e-07,
-1.00907686828577e-06,
-1.03381182725570e-06,
-1.05901119695773e-06,
-1.08468134385475e-06,
-1.11082817966235e-06,
-1.13745784346975e-06,
-1.16457613330567e-06,
-1.19218918825936e-06,
-1.22030314742005e-06,
-1.24892403619015e-06,
-1.27805799365888e-06,
-1.30771138628916e-06,
-1.33789058054390e-06,
-1.36860182919918e-06,
-1.39985127134423e-06,
-1.43164527344197e-06,
-1.46399020195531e-06,
-1.49689276440768e-06,
-1.53035921357514e-06,
-1.56439625698113e-06,
-1.59901037477539e-06,
-1.63420816079451e-06,
-1.66999598150142e-06,
-1.70638043073268e-06,
-1.74336821601173e-06,
-1.78096604486200e-06,
-1.81918051112007e-06,
-1.85801832230936e-06,
-1.89748629964015e-06,
-1.93759137800953e-06,
-1.97834015125409e-06,
-2.01973989533144e-06,
-2.06179674933082e-06,
-2.10451798920985e-06,
-2.14790998143144e-06,
-2.19198000195320e-06,
-2.23673396249069e-06,
-2.28217913900153e-06,
-2.32832258006965e-06,
-2.37517065215798e-06,
-2.42273108597146e-06,
-2.47101070272038e-06,
-2.52001632361498e-06,
-2.56975545198657e-06,
-2.62023536379274e-06,
-2.67146310761746e-06,
-2.72344641416566e-06,
-2.77619210464763e-06,
-2.82970790976833e-06,
-2.88400087811169e-06,
-2.93907851300901e-06,
-2.99494854516524e-06,
-3.05161779579066e-06,
-3.10909445033758e-06,
-3.16738533001626e-06,
-3.22649771078432e-06,
-3.28643909597304e-06,
-3.34721607941901e-06,
-3.40883639182721e-06,
-3.47130685440789e-06,
-3.53463451574498e-06,
-3.59882665179612e-06,
-3.66389008377155e-06,
-3.72983208762889e-06,
-3.79665948457841e-06,
-3.86437932320405e-06,
-3.93299933421076e-06,
-4.00252702092985e-06,
-4.07296874982421e-06,
-4.14433270634618e-06,
-4.21662571170600e-06,
-4.28985504186130e-06,
-4.36402888226439e-06,
-4.43915405412554e-06,
-4.51523828814970e-06,
-4.59228931504185e-06,
-4.67031486550695e-06,
-4.74932085126056e-06,
-4.82931636724970e-06,
-4.91030823468464e-06,
-4.99230372952297e-06,
-5.07531103721703e-06,
-5.15933788847178e-06,
-5.24439246873953e-06,
-5.33048250872525e-06,
-5.41761528438656e-06,
-5.50579898117576e-06,
-5.59504223929253e-06,
-5.68535233469447e-06,
-5.77673790758126e-06,
-5.86920714340522e-06,
-5.96276822761865e-06,
-6.05742980042123e-06,
-6.15320050201262e-06,
-6.25008851784514e-06,
-6.34810294286581e-06,
-6.44725241727429e-06,
-6.54754512652289e-06,
-6.64899016555864e-06,
-6.75159571983386e-06,
-6.85536997480085e-06,
-6.96032202540664e-06,
-7.06646005710354e-06,
-7.17379316483857e-06,
-7.28232907931670e-06,
-7.39207735023228e-06,
-7.50304616303765e-06,
-7.61524370318512e-06,
-7.72867952036904e-06,
-7.84336134529440e-06,
-7.95929736341350e-06,
-8.07649848866276e-06,
-8.19497199699981e-06,
-8.31472789286636e-06,
-8.43577436171472e-06,
-8.55812231748132e-06,
-8.68177903612377e-06,
-8.80675361258909e-06,
-8.93305514182430e-06,
-9.06069453776581e-06,
-9.18967907637125e-06,
-9.32001876208233e-06,
-9.45172268984607e-06,
-9.58479904511478e-06,
-9.71925874182489e-06,
-9.85510996542871e-06,
-9.99236090137856e-06,
-1.01310215541162e-05,
-1.02711001090938e-05,
-1.04126056612586e-05,
-1.05555482150521e-05,
-1.06999341369374e-05,
-1.08457743408508e-05,
-1.09930779217393e-05,
-1.11418521555606e-05,
-1.12921088657458e-05,
-1.14438553282525e-05,
-1.15971006380278e-05,
-1.17518557090079e-05,
-1.19081278171507e-05,
-1.20659269668977e-05,
-1.22252622531960e-05,
-1.23861445899820e-05,
-1.25485812532133e-05,
-1.27125831568264e-05,
-1.28781584862736e-05,
-1.30453181554913e-05,
-1.32140703499317e-05,
-1.33844250740367e-05,
-1.35563932417426e-05,
-1.37299830385018e-05,
-1.39052053782507e-05,
-1.40820684464416e-05,
-1.42605831570108e-05,
-1.44407595144003e-05,
-1.46226066135569e-05,
-1.48061335494276e-05,
-1.49913512359490e-05,
-1.51782687680679e-05,
-1.53668952407315e-05,
-1.55572415678762e-05,
-1.57493159349542e-05,
-1.59431274369126e-05,
-1.61386888066772e-05,
-1.63360055012163e-05,
-1.65350920724450e-05,
-1.67359539773315e-05,
-1.69386039488018e-05,
-1.71430492628133e-05,
-1.73493008333026e-05,
-1.75573695742060e-05,
-1.77672627614811e-05,
-1.79789894900750e-05,
-1.81925643119030e-05,
-1.84079926839331e-05,
-1.86252873390913e-05,
-1.88444591913139e-05,
-1.90655155165587e-05,
-1.92884708667407e-05,
-1.95133306988282e-05,
-1.97401095647365e-05,
-1.99688165594125e-05,
-2.01994607778033e-05,
-2.04320549528347e-05,
-2.06666081794538e-05,
-2.09031277336180e-05,
-2.11416299862321e-05,
-2.13821185752749e-05,
-2.16246062336722e-05,
-2.18691038753605e-05,
-2.21156187762972e-05,
-2.23641636694083e-05,
-2.26147476496408e-05,
-2.28673816309311e-05,
-2.31220747082261e-05,
-2.33788377954625e-05,
-2.36376818065764e-05,
-2.38986176555045e-05,
-2.41616526182042e-05,
-2.44268030655803e-05,
-2.46940744546009e-05,
-2.49634813371813e-05,
-2.52350346272578e-05,
-2.55087434197776e-05,
-2.57846186286770e-05,
-2.60626711678924e-05,
-2.63429137703497e-05,
-2.66253573499853e-05,
-2.69100091827568e-05,
-2.71968838205794e-05,
-2.74859903584002e-05,
-2.77773397101555e-05,
-2.80709464277606e-05,
-2.83668196061626e-05,
-2.86649701592978e-05,
-2.89654071821133e-05,
-2.92681452265242e-05,
-2.95731952064671e-05,
-2.98805662168888e-05,
-3.01902728097048e-05,
-3.05023240798619e-05,
-3.08167327602860e-05,
-3.11335061269347e-05,
-3.14526623697020e-05,
-3.17742051265668e-05,
-3.20981525874231e-05,
-3.24245120282285e-05,
-3.27532980008982e-05,
-3.30845177813899e-05,
-3.34181895595975e-05,
-3.37543169735000e-05,
-3.40929218509700e-05,
-3.44340078299865e-05,
-3.47775894624647e-05,
-3.51236740243621e-05,
-3.54722797055729e-05,
-3.58234137820546e-05,
-3.61770908057224e-05,
-3.65333253284916e-05,
-3.68921246263199e-05,
-3.72535032511223e-05,
-3.76174684788566e-05,
-3.79840348614380e-05,
-3.83532169507816e-05,
-3.87250256608240e-05,
-3.90994719055016e-05,
-3.94765702367295e-05,
-3.98563315684442e-05,
-4.02387631766032e-05,
-4.06238868890796e-05,
-4.10117063438520e-05,
-4.14022324548569e-05,
-4.17954834119882e-05,
-4.21914701291826e-05,
-4.25902035203762e-05,
-4.29916944995057e-05,
-4.33959539805073e-05,
-4.38029965152964e-05,
-4.42128366557881e-05,
-4.46254816779401e-05,
-4.50409497716464e-05,
-4.54592445748858e-05,
-4.58803806395736e-05,
-4.63043725176249e-05,
-4.67312311229762e-05,
-4.71609710075427e-05,
-4.75935994472820e-05,
-4.80291309941094e-05,
-4.84675801999401e-05,
-4.89089616166893e-05,
-4.93532788823359e-05,
-4.98005501867738e-05,
-5.02507900819182e-05,
-5.07040058437269e-05,
-5.11602193000726e-05,
-5.16194340889342e-05,
-5.20816611242481e-05,
-5.25469222338870e-05,
-5.30152210558299e-05,
-5.34865721419919e-05,
-5.39609900442883e-05,
-5.44384856766555e-05,
-5.49190735910088e-05,
-5.54027647012845e-05,
-5.58895735593978e-05,
-5.63795110792853e-05,
-5.68725918128621e-05,
-5.73688230360858e-05,
-5.78682265768293e-05,
-5.83708060730714e-05,
-5.88765760767274e-05,
-5.93855511397123e-05,
-5.98977421759628e-05,
-6.04131673753727e-05,
-6.09318376518786e-05,
-6.14537639194168e-05,
-6.19789570919238e-05,
-6.25074317213148e-05,
-6.30392023595050e-05,
-6.35742908343673e-05,
-6.41126971459016e-05,
-6.46544358460233e-05,
-6.51995214866474e-05,
-6.57479758956470e-05,
-6.62998063489795e-05,
-6.68550273985602e-05,
-6.74136390443891e-05,
-6.79756703902967e-05,
-6.85411287122406e-05,
-6.91100285621360e-05,
-6.96823844918981e-05,
-7.02582037774846e-05,
-7.08375082467683e-05,
-7.14203051757067e-05,
-7.20066163921729e-05,
-7.25964418961667e-05,
-7.31897962396033e-05,
-7.37867012503557e-05,
-7.43871642043814e-05,
-7.49912069295533e-05,
-7.55988367018290e-05,
-7.62100680731237e-05,
-7.68249155953527e-05,
-7.74433865444735e-05,
-7.80655100243166e-05,
-7.86912860348821e-05,
-7.93207364040427e-05,
-7.99538756837137e-05,
-8.05907111498527e-05,
-8.12312646303326e-05,
-8.18755434011109e-05,
-8.25235547381453e-05,
-8.31753277452663e-05,
-8.38308624224737e-05,
-8.44901805976406e-05,
-8.51532895467244e-05,
-8.58202038216405e-05,
-8.64909452502616e-05,
-8.71655283845030e-05,
-8.78439459484071e-05,
-8.85262343217619e-05,
-8.92123935045674e-05,
-8.99024598766118e-05,
-9.05964188859798e-05,
-9.12943069124594e-05,
-9.19961239560507e-05,
-9.27018991205841e-05,
-9.34116251301020e-05,
-9.41253383643925e-05,
-9.48430460994132e-05,
-9.55647628870793e-05,
-9.62904960033484e-05,
-9.70202672760934e-05,
-9.77540985331871e-05,
-9.84919897746295e-05,
-9.92339701042511e-05,
-9.99800395220518e-05,
-0.000100730227131862,
-0.000101484540209640,
-0.000102242993307300,
-0.000103005600976758,
-0.000103772377769928,
-0.000104543338238727,
-0.000105318504211027,
-0.000106097875686828,
-0.000106881481769960,
-0.000107669329736382,
-0.000108461434138007,
-0.000109257802250795,
-0.000110058470454533,
-0.000110863438749220,
-0.000111672714410815,
-0.000112486333819106,
-0.000113304296974093,
-0.000114126618427690,
-0.000114953320007771,
-0.000115784408990294,
-0.000116619907203130,
-0.000117459829198197,
-0.000118304189527407,
-0.000119152995466720,
-0.000120006283395924,
-0.000120864046039060,
-0.000121726312499959,
-0.000122593090054579,
-0.000123464400530793,
-0.000124340251204558,
-0.000125220656627789,
-0.000126105631352402,
-0.000126995204482228,
-0.000127889405121095,
-0.000128788218717091,
-0.000129691659822129,
-0.000130599772091955,
-0.000131512540974654,
-0.000132429995574057,
-0.000133352179545909,
-0.000134279063786380,
-0.000135210677399300,
-0.000136147049488500,
-0.000137088194605894,
-0.000138034127303399,
-0.000138984847581014,
-0.000139940384542570,
-0.000140900767291896,
-0.000141865995828994,
-0.000142836084705777,
-0.000143811048474163,
-0.000144790930789895,
-0.000145775717101060,
-0.000146765436511487,
-0.000147760103573091,
-0.000148759732837789,
-0.000149764338857494,
-0.000150773936184123,
-0.000151788568473421,
-0.000152808206621557,
-0.000153832908836193,
-0.000154862675117329,
-0.000155897520016879,
-0.000156937443534844,
-0.000157982489326969,
-0.000159032671945170,
-0.000160087991389446,
-0.000161148476763628,
-0.000162214142619632,
-0.000163285003509372,
-0.000164361088536680,
-0.000165442397701554,
-0.000166528945555910,
-0.000167620775755495,
-0.000168717873748392,
-0.000169820268638432,
-0.000170927974977531,
-0.000172041007317603,
-0.000173159394762479,
-0.000174283137312159,
-0.000175412278622389,
-0.000176546804141253,
-0.000177686742972583,
-0.000178832109668292,
-0.000179982904228382,
-0.000181139199412428,
-0.000182300951564685,
-0.000183468189788982,
-0.000184640957741067,
-0.000185819240869023,
-0.000187003082828596,
-0.000188192483619787,
-0.000189387472346425,
-0.000190588049008511,
-0.000191794228157960,
-0.000193006068002433,
-0.000194223539438099,
-0.000195446671568789,
-0.000196675478946418,
-0.000197909990674816,
-0.000199150206753984,
-0.000200396170839667,
-0.000201647882931866,
-0.000202905357582495,
-0.000204168609343469,
-0.000205437652766705,
-0.000206712531507947,
-0.000207993245567195,
-0.000209279809496366,
-0.000210572237847373,
-0.000211870559724048,
-0.000213174789678305,
-0.000214484942262061,
-0.000215801032027230,
-0.000217123088077642,
-0.000218451110413298,
-0.000219785113586113,
-0.000221125141251832,
-0.000222471207962371,
-0.000223823299165815,
-0.000225181458517909,
-0.000226545700570568,
-0.000227916054427624,
-0.000229292520089075,
-0.000230675112106837,
-0.000232063874136657,
-0.000233458791626617,
-0.000234859908232465,
-0.000236267223954201,
-0.000237680767895654,
-0.000239100569160655,
-0.000240526613197289,
-0.000241958943661302,
-0.000243397575104609,
-0.000244842522079125,
-0.000246293784584850,
-0.000247751420829445,
-0.000249215430812910,
-0.000250685814535245,
-0.000252162630204111,
-0.000253645877819508,
-0.000255135528277606,
-0.000256631697993726,
-0.000258134299656376,
-0.000259643420577049,
-0.000261159089859575,
-0.000262681278400123,
-0.000264210015302524,
-0.000265745329670608,
-0.000267287250608206,
-0.000268835778115317,
-0.000270390941295773,
-0.000271952769253403,
-0.000273521261988208,
-0.000275096419500187,
-0.000276678270893171,
-0.000278266874374822,
-0.000279862200841308,
-0.000281464279396459,
-0.000283073110040277,
-0.000284688780084252,
-0.000286311231320724,
-0.000287940521957353,
-0.000289576651994139,
-0.000291219650534913,
-0.000292869546683505,
-0.000294526340439916,
-0.000296190031804144,
-0.000297860678983852,
-0.000299538311082870,
-0.000301222898997366,
-0.000302914471831173,
-0.000304613058688119,
-0.000306318688672036,
-0.000308031361782923,
-0.000309751107124612,
-0.000311477924697101,
-0.000313211901811883,
-0.000314952980261296,
-0.000316701189149171,
-0.000318456586683169,
-0.000320219172863290,
-0.000321988947689533,
-0.000323765969369561,
-0.000325550208799541,
-0.000327341724187136,
-0.000329140515532345,
-0.000330946641042829,
-0.000332760071614757,
-0.000334580836351961,
-0.000336408964358270,
-0.000338244484737515,
-0.000340087397489697,
-0.000341937731718645,
-0.000343795487424359,
-0.000345660751918331,
-0.000347533466992900,
-0.000349413690855727,
-0.000351301394402981,
-0.000353196664946154,
-0.000355099502485245,
-0.000357009936124086,
-0.000358927936758846,
-0.000360853562597185,
-0.000362786813639104,
-0.000364727718988434,
-0.000366676336852834,
-0.000368632638128474,
-0.000370596681023017,
-0.000372568465536460,
-0.000374548020772636,
-0.000376535346731544,
-0.000378530443413183,
-0.000380533398129046,
-0.000382544181775302,
-0.000384562852559611,
-0.000386589410481975,
-0.000388623855542392,
-0.000390666245948523,
-0.000392716581700370,
-0.000394774921005592,
-0.000396841234760359,
-0.000398915552068502,
-0.000400997902033851,
-0.000403088313760236,
-0.000405186816351488,
-0.000407293409807608,
-0.000409408094128594,
-0.000411530956625938,
-0.000413661939091980,
-0.000415801128838211,
-0.000417948525864631,
-0.000420104130171239,
-0.000422267999965698,
-0.000424440135248005,
-0.000426620536018163,
-0.000428809289587662,
-0.000431006366852671,
-0.000433211767813191,
-0.000435425579780713,
-0.000437647802755237,
-0.000439878436736763,
-0.000442117510829121,
-0.000444365083239973,
-0.000446621124865487,
-0.000448885664809495,
-0.000451158761279658,
-0.000453440414275974,
-0.000455730652902275,
-0.000458029506262392,
-0.000460336974356324,
-0.000462653115391731,
-0.000464977900264785,
-0.000467311358079314,
-0.000469653576146811,
-0.000472004525363445,
-0.000474364234833047,
-0.000476732733659446,
-0.000479110050946474,
-0.000481496215797961,
-0.000483891228213906,
-0.000486295117298141,
-0.000488707912154496,
-0.000491129583679140,
-0.000493560277391225,
-0.000495999876875430,
-0.000498448498547077,
-0.000500906200613827,
-0.000503372866660357,
-0.000505848671309650,
-0.000508333498146385,
-0.000510827463585883,
-0.000513330567628145,
-0.000515842868480831,
-0.000518364307936281,
-0.000520895002409816,
-0.000523434951901436,
-0.000525984098203480,
-0.000528542557731271,
-0.000531110214069486,
-0.000533687300048769,
-0.000536273641046137,
-0.000538869411684573,
-0.000541474553756416,
-0.000544089125469327,
-0.000546713126823306,
-0.000549346674233675,
-0.000551989709492773,
-0.000554642174392939,
-0.000557304243557155,
-0.000559975916985422,
-0.000562657136470079,
-0.000565348018426448,
-0.000568048504646868,
-0.000570758711546660,
-0.000573478522710502,
-0.000576208112761378,
-0.000578947481699288,
-0.000581696571316570,
-0.000584455556236208,
-0.000587224261835218,
-0.000590002862736583,
-0.000592791300732642,
-0.000595589634031057,
-0.000598397920839489,
-0.000601216102950275,
-0.000604044296778739,
-0.000606882444117218,
-0.000609730661381036,
-0.000612588948570192,
-0.000615457247477025,
-0.000618335674516857,
-0.000621224287897348,
-0.000624123029410839,
-0.000627031957264990,
-0.000629951013252139,
-0.000632880371995270,
-0.000635819975286722,
-0.000638769881334156,
-0.000641730090137571,
-0.000644700659904629,
-0.000647681590635330,
-0.000650672882329673,
-0.000653674651402980,
-0.000656686839647591,
-0.000659709505271167,
-0.000662742648273706,
-0.000665786326862872,
-0.000668840541038662,
-0.000671905349008739,
-0.000674980750773102,
-0.000678066804539412,
-0.000681163510307670,
-0.000684270926285535,
-0.000687389052473009,
-0.000690517888870090,
-0.000693657551892102,
-0.000696807983331382,
-0.000699969241395593,
-0.000703141326084733,
-0.000706324353814125,
-0.000709518266376108,
-0.000712723121978343,
-0.000715938920620829,
-0.000719165720511228,
-0.000722403521649540,
-0.000725652440451086,
-0.000728912418708205,
-0.000732183456420898,
-0.000735465611796826,
-0.000738759001251310,
-0.000742063508369029,
-0.000745379249565303,
-0.000748706224840134,
-0.000752044550608844,
-0.000755394168663770,
-0.000758755137212575,
-0.000762127398047596,
-0.000765511125791818,
-0.000768906204029918,
-0.000772312749177218,
-0.000775730761233717,
-0.000779160298407078,
-0.000782601360697299,
-0.000786054006312043,
-0.000789518235251308,
-0.000792994105722755,
-0.000796481617726386,
-0.000799980829469860,
-0.000803491799160838,
-0.000807014468591660,
-0.000810548895969987,
-0.000814095139503479,
-0.000817653140984476,
-0.000821223075035960,
-0.000824804883450270,
-0.000828398624435067,
-0.000832004297990352,
-0.000835621962323785,
-0.000839251617435366,
-0.000842893321532756,
-0.000846547074615955,
-0.000850212934892625,
-0.000853890902362764,
-0.000857581035234034,
-0.000861283333506435,
-0.000864997913595289,
-0.000868724717292935,
-0.000872463744599372,
-0.000876215170137584,
-0.000879978877492249,
-0.000883754983078688,
-0.000887543428689241,
-0.000891344330739230,
-0.000895157747436315,
-0.000898983620572835,
-0.000902822066564113,
-0.000906672968994826,
-0.000910536502487958,
-0.000914412725251168,
-0.000918301520869136,
-0.000922203005757183,
-0.000926117179915309,
-0.000930044159758836,
-0.000933983887080103,
-0.000937936361879110,
-0.000941901758778840,
-0.000945880019571632,
-0.000949871144257486,
-0.000953875191044062,
-0.000957892218139023,
-0.000961922283750027,
-0.000965965387877077,
-0.000970021472312510,
-0.000974090653471649,
-0.000978172989562154,
-0.000982268480584025,
-0.000986377126537263,
-0.000990499043837190,
-0.000994634116068482,
-0.000998782459646463,
-0.00100294419098645,
-0.00100711931008846,
-0.00101130781695247,
-0.00101550959516317,
-0.00101972487755120,
-0.00102395366411656,
-0.00102819583844394,
-0.00103245174977928,
-0.00103672104887664,
-0.00104100408498198,
-0.00104530062526464,
-0.00104961078613997,
-0.00105393480043858,
-0.00105827255174518,
-0.00106262404005975,
-0.00106698926538229,
-0.00107136834412813,
-0.00107576127629727,
-0.00108016817830503,
-0.00108458893373609,
-0.00108902365900576,
-0.00109347247052938,
-0.00109793525189161,
-0.00110241223592311,
-0.00110690318979323,
-0.00111140834633261,
-0.00111592758912593,
-0.00112046103458852,
-0.00112500879913569,
-0.00112957076635212,
-0.00113414716906846,
-0.00113873777445406,
-0.00114334269892424,
-0.00114796217530966,
-0.00115259597077966,
-0.00115724431816489,
-0.00116190710105002,
-0.00116658443585038,
-0.00117127632256597,
-0.00117598287761211,
-0.00118070410098881,
-0.00118543987628073,
-0.00119019055273384,
-0.00119495589751750,
-0.00119973602704704,
-0.00120453094132245,
-0.00120934064034373,
-0.00121416524052620,
-0.00121900474186987,
-0.00122385926079005,
-0.00122872868087143,
-0.00123361323494464,
-0.00123851269017905,
-0.00124342727940530,
-0.00124835711903870,
-0.00125330197624862,
-0.00125826196745038,
-0.00126323732547462,
-0.00126822793390602,
-0.00127323379274458,
-0.00127825501840562,
-0.00128329149447382,
-0.00128834357019514,
-0.00129341089632362,
-0.00129849382210523,
-0.00130359211470932,
-0.00130870612338185,
-0.00131383549887687,
-0.00131898059044033,
-0.00132414139807224,
-0.00132931768894196,
-0.00133450981229544,
-0.00133971765171736,
-0.00134494132362306,
-0.00135018071159720,
-0.00135543593205512,
-0.00136070710141212,
-0.00136599410325289,
-0.00137129717040807,
-0.00137661618646234,
-0.00138195126783103,
-0.00138730229809880,
-0.00139266939368099,
-0.00139805278740823,
-0.00140345224644989,
-0.00140886788722128,
-0.00141429970972240,
-0.00141974783036858,
-0.00142521224915981,
-0.00143069308251143,
-0.00143619021400809,
-0.00144170387648046,
-0.00144723383709788,
-0.00145278021227568,
-0.00145834323484451,
-0.00146392278838903,
-0.00146951887290925,
-0.00147513160482049,
-0.00148076098412275,
-0.00148640701081604,
-0.00149206980131567,
-0.00149774935562164,
-0.00150344567373395,
-0.00150915887206793,
-0.00151488883420825,
-0.00152063579298556,
-0.00152639963198453,
-0.00153218046762049,
-0.00153797829989344,
-0.00154379312880337,
-0.00154962507076561,
-0.00155547412578017,
-0.00156134029384702,
-0.00156722369138151,
-0.00157312431838363,
-0.00157904217485338,
-0.00158497737720609,
-0.00159092980902642,
-0.00159689970314503,
-0.00160288705956191,
-0.00160889164544642,
-0.00161491381004453,
-0.00162095343694091,
-0.00162701064255089,
-0.00163308542687446,
-0.00163917778991163,
-0.00164528784807771,
-0.00165141548495740,
-0.00165756093338132,
-0.00166372419334948,
-0.00166990514844656,
-0.00167610391508788,
-0.00168232049327344,
-0.00168855499941856,
-0.00169480743352324,
-0.00170107791200280,
-0.00170736631844193,
-0.00171367276925594,
-0.00171999726444483,
-0.00172633992042393,
-0.00173270073719323,
-0.00173907959833741,
-0.00174547685310245,
-0.00175189226865768,
-0.00175832607783377,
-0.00176477816421539,
-0.00177124852780253,
-0.00177773728501052,
-0.00178424455225468,
-0.00179077021311969,
-0.00179731450043619,
-0.00180387718137354,
-0.00181045848876238,
-0.00181705853901804,
-0.00182367698289454,
-0.00183031428605318,
-0.00183697021566331,
-0.00184364500455558,
-0.00185033853631467,
-0.00185705081094056,
-0.00186378206126392,
-0.00187053205445409,
-0.00187730102334172,
-0.00188408896792680,
-0.00189089600462466,
-0.00189772190060467,
-0.00190456688869745,
-0.00191143108531833,
-0.00191831437405199,
-0.00192521675489843,
-0.00193213846068829,
-0.00193907937500626,
-0.00194603961426765,
-0.00195301906205714,
-0.00196001795120537,
-0.00196703616529703,
-0.00197407370433211,
-0.00198113080114126,
-0.00198820722289383,
-0.00199530320242047,
-0.00200241897255182,
-0.00200955406762660,
-0.00201670895330608,
-0.00202388339675963,
-0.00203107763081789,
-0.00203829142265022,
-0.00204552523791790,
-0.00205277861095965,
-0.00206005200743675,
-0.00206734519451857,
-0.00207465840503573,
-0.00208199140615761,
-0.00208934443071485,
-0.00209671747870743,
-0.00210411031730473,
-0.00211152341216803,
-0.00211895676329732,
-0.00212641037069261,
-0.00213388400152326,
-0.00214137788861990,
-0.00214889203198254,
-0.00215642643161118,
-0.00216398108750582,
-0.00217155623249710,
-0.00217915163375437,
-0.00218676752410829,
-0.00219440390355885,
-0.00220206077210605,
-0.00220973836258054,
-0.00221743620932102,
-0.00222515501081944,
-0.00223289430141449,
-0.00224065408110619,
-0.00224843504838645,
-0.00225623627193272,
-0.00226405868306756,
-0.00227190181612968,
-0.00227976590394974,
-0.00228765071369708,
-0.00229555647820234,
-0.00230348319746554,
-0.00231143110431731,
-0.00231939973309636,
-0.00232738954946399,
-0.00233540055342019,
-0.00234343274496496,
-0.00235148589126766,
-0.00235956045798957,
-0.00236765621230006,
-0.00237577338702977,
-0.00238391174934804,
-0.00239207153208554,
-0.00240025273524225,
-0.00240845535881817,
-0.00241667940281332,
-0.00242492510005832,
-0.00243319245055318,
-0.00244148122146726,
-0.00244979141280055,
-0.00245812349021435,
-0.00246647722087801,
-0.00247485283762217,
-0.00248325010761619,
-0.00249166926369071,
-0.00250011030584574,
-0.00250857300125062,
-0.00251705781556666,
-0.00252556428313255,
-0.00253409310244024,
-0.00254264404065907,
-0.00255121686495841,
-0.00255981180816889,
-0.00256842887029052,
-0.00257706805132329,
-0.00258572958409786,
-0.00259441323578358,
-0.00260311923921108,
-0.00261184759438038,
-0.00262059830129147,
-0.00262937135994434,
-0.00263816700316966,
-0.00264698499813676,
-0.00265582557767630,
-0.00266468874178827,
-0.00267357449047267,
-0.00268248282372952,
-0.00269141397438943,
-0.00270036770962179,
-0.00270934426225722,
-0.00271834363229573,
-0.00272736581973732,
-0.00273641059175134,
-0.00274547864682972,
-0.00275456951931119,
-0.00276368320919573,
-0.00277282018214464,
-0.00278198020532727,
-0.00279116327874362,
-0.00280036940239370,
-0.00280959880910814,
-0.00281885126605630,
-0.00282812700606883,
-0.00283742602914572,
-0.00284674856811762,
-0.00285609415732324,
-0.00286546349525452,
-0.00287485611625016,
-0.00288427225314081,
-0.00289371190592647,
-0.00290317507460713,
-0.00291266175918281,
-0.00292217219248414,
-0.00293170637451112,
-0.00294126407243311,
-0.00295084551908076,
-0.00296045118011534,
-0.00297008035704494,
-0.00297973328270018,
-0.00298941042274237,
-0.00299911107867956,
-0.00300883594900370,
-0.00301858480088413,
-0.00302835763432086,
-0.00303815491497517,
-0.00304797617718577,
-0.00305782165378332,
-0.00306769111193717,
-0.00307758478447795,
-0.00308750290423632,
-0.00309744523838162,
-0.00310741225257516,
-0.00311740348115563,
-0.00312741915695369,
-0.00313745927996933,
-0.00314752385020256,
-0.00315761310048401,
-0.00316772703081369,
-0.00317786540836096,
-0.00318802869878709,
-0.00319821643643081,
-0.00320842908695340,
-0.00321866665035486,
-0.00322892912663519,
-0.00323921628296375,
-0.00324952811934054,
-0.00325986510142684,
-0.00327022699639201,
-0.00328061403706670,
-0.00329102599062026,
-0.00330146308988333,
-0.00331192556768656,
-0.00332241319119930,
-0.00333292596042156,
-0.00334346410818398,
-0.00335402740165591,
-0.00336461607366800,
-0.00337522989138961,
-0.00338586932048202,
-0.00339653436094522,
-0.00340722477994859,
-0.00341794057749212,
-0.00342868221923709,
-0.00343944923952222,
-0.00345024233683944,
-0.00346106081269681,
-0.00347190513275564,
-0.00348277506418526,
-0.00349367107264698,
-0.00350459292531014,
-0.00351554062217474,
-0.00352651416324079,
-0.00353751378133893,
-0.00354853947646916,
-0.00355959124863148,
-0.00357066909782589,
-0.00358177302405238,
-0.00359290302731097,
-0.00360405957326293,
-0.00361524242907763,
-0.00362645136192441,
-0.00363768683746457,
-0.00364894862286747,
-0.00366023695096374,
-0.00367155158892274,
-0.00368289300240576,
-0.00369426072575152,
-0.00370565499179065,
-0.00371707603335381,
-0.00372852385044098,
-0.00373999844305217,
-0.00375149981118739,
-0.00376302795484662,
-0.00377458287402988,
-0.00378616480156779,
-0.00379777350462973,
-0.00380940944887698,
-0.00382107240147889,
-0.00383276212960482,
-0.00384447933174670,
-0.00385622354224324,
-0.00386799476109445,
-0.00387979345396161,
-0.00389161938801408,
-0.00390347279608250,
-0.00391535321250558,
-0.00392726156860590,
-0.00393919693306088,
-0.00395116023719311,
-0.00396315054968000,
-0.00397516880184412,
-0.00398721452802420,
-0.00399928772822022,
-0.00401138886809349,
-0.00402351794764400,
-0.00403567450121045,
-0.00404785899445415,
-0.00406007142737508,
-0.00407231179997325,
-0.00408458011224866,
-0.00409687636420131,
-0.00410920055583119,
-0.00412155315279961,
-0.00413393368944526,
-0.00414634216576815,
-0.00415877904742956,
-0.00417124433442950,
-0.00418373756110668,
-0.00419625965878367,
-0.00420880969613791,
-0.00422138860449195,
-0.00423399545252323,
-0.00424663117155433,
-0.00425929529592395,
-0.00427198782563210,
-0.00428470969200134,
-0.00429745996370912,
-0.00431023910641670,
-0.00432304665446281,
-0.00433588353917003,
-0.00434874882921577,
-0.00436164345592260,
-0.00437456695362926,
-0.00438751932233572,
-0.00440050102770329,
-0.00441351160407066,
-0.00442655105143786,
-0.00443962030112743,
-0.00445271842181683,
-0.00446584587916732,
-0.00447900267317891,
-0.00449218880385160,
-0.00450540427118540,
-0.00451864954084158,
-0.00453192414715886,
-0.00454522855579853,
-0.00455856230109930,
-0.00457192538306117,
-0.00458531873300672,
-0.00459874141961336,
-0.00461219390854240,
-0.00462567619979382,
-0.00463918875902891,
-0.00465273112058640,
-0.00466630328446627,
-0.00467990525066853,
-0.00469353748485446,
-0.00470719998702407,
-0.00472089275717735,
-0.00473461532965303,
-0.00474836863577366,
-0.00476215174421668,
-0.00477596512064338,
-0.00478980923071504,
-0.00480368360877037,
-0.00481758872047067,
-0.00483152410015464,
-0.00484549021348357,
-0.00485948706045747,
-0.00487351464107633,
-0.00488757248967886,
-0.00490166107192636,
-0.00491578085348010,
-0.00492993136867881,
-0.00494411215186119,
-0.00495832460001111,
-0.00497256778180599,
-0.00498684169724584,
-0.00500114727765322,
-0.00501548359170556,
-0.00502985157072544,
-0.00504425028339028,
-0.00505868019536138,
-0.00507314177230001,
-0.00508763454854488,
-0.00510215852409601,
-0.00511671416461468,
-0.00513130100443959,
-0.00514591950923204,
-0.00516056967899203,
-0.00517525104805827,
-0.00518996454775333,
-0.00520470924675465,
-0.00521948607638478,
-0.00523429503664374,
-0.00524913566187024,
-0.00526400795206428,
-0.00527891283854842,
-0.00529384892433882,
-0.00530881760641933,
-0.00532381841912866,
-0.00533885089680553,
-0.00535391550511122,
-0.00536901270970702,
-0.00538414204493165,
-0.00539930397644639,
-0.00541449803858995,
-0.00542972469702363,
-0.00544498395174742,
-0.00546027533710003,
-0.00547559978440404,
-0.00549095589667559,
-0.00550634553655982,
-0.00552176730707288,
-0.00553722213953733,
-0.00555271003395319,
-0.00556823052465916,
-0.00558378407731652,
-0.00559937022626400,
-0.00561498990282416,
-0.00563064217567444,
-0.00564632751047611,
-0.00566204637289047,
-0.00567779829725623,
-0.00569358328357339,
-0.00570940179750323,
-0.00572525383904576,
-0.00574113894253969,
-0.00575705757364631,
-0.00577300926670432,
-0.00578899495303631,
-0.00580501416698098,
-0.00582106690853834,
-0.00583715364336968,
-0.00585327344015241,
-0.00586942723020911,
-0.00588561501353979,
-0.00590183632448316,
-0.00591809162870050,
-0.00593438139185309,
-0.00595070514827967,
-0.00596706243231893,
-0.00598345417529345,
-0.00599987991154194,
-0.00601633964106441,
-0.00603283429518342,
-0.00604936294257641,
-0.00606592604890466,
-0.00608252361416817,
-0.00609915563836694,
-0.00611582165583968,
-0.00613252306357026,
-0.00614925846457481,
-0.00616602832451463,
-0.00618283357471228,
-0.00619967328384519,
-0.00621654745191336,
-0.00623345654457808,
-0.00625040056183934,
-0.00626737950369716,
-0.00628439383581281,
-0.00630144309252501,
-0.00631852727383375,
-0.00633564684540033,
-0.00635280134156346,
-0.00636999122798443,
-0.00638721650466323,
-0.00640447670593858,
-0.00642177276313305,
-0.00643910374492407,
-0.00645647058263421,
-0.00647387281060219,
-0.00649131089448929,
-0.00650878483429551,
-0.00652629369869828,
-0.00654383888468146,
-0.00656141946092248,
-0.00657903589308262,
-0.00659668818116188,
-0.00661437679082155,
-0.00663210125640035,
-0.00664986204355955,
-0.00666765822097659,
-0.00668549118563533,
-0.00670336000621319,
-0.00672126514837146,
-0.00673920661211014,
-0.00675718486309052,
-0.00677519850432873,
-0.00679324939846993,
-0.00681133614853025,
-0.00682946015149355,
-0.00684762001037598,
-0.00686581665650010,
-0.00688405055552721,
-0.00690232077613473,
-0.00692062778398395,
-0.00693897157907486,
-0.00695735262706876,
-0.00697577046230435,
-0.00699422508478165,
-0.00701271649450064,
-0.00703124515712261,
-0.00704981153830886,
-0.00706841470673680,
-0.00708705512806773,
-0.00710573326796293,
-0.00712444819509983,
-0.00714320084080100,
-0.00716199073940516,
-0.00718081789091229,
-0.00719968276098371,
-0.00721858534961939,
-0.00723752519115806,
-0.00725650321692228,
-0.00727551849558950,
-0.00729457195848227,
-0.00731366313993931,
-0.00733279203996062,
-0.00735195912420750,
-0.00737116392701864,
-0.00739040737971664,
-0.00740968855097890,
-0.00742900790646672,
-0.00744836544618011,
-0.00746776117011905,
-0.00748719507828355,
-0.00750666763633490,
-0.00752617837861180,
-0.00754572777077556,
-0.00756531534716487,
-0.00758494157344103,
-0.00760460644960403,
-0.00762431044131517,
-0.00764405261725187,
-0.00766383344307542,
-0.00768365291878581,
-0.00770351197570562,
-0.00772340921685100,
-0.00774334603920579,
-0.00776332151144743,
-0.00778333609923720,
-0.00780339026823640,
-0.00782348308712244,
-0.00784361548721790,
-0.00786378700286150,
-0.00788399763405323,
-0.00790424831211567,
-0.00792453717440367,
-0.00794486608356237,
-0.00796523503959179,
-0.00798564311116934,
-0.00800609029829502,
-0.00802657846361399,
-0.00804710481315851,
-0.00806767120957375,
-0.00808827858418226,
-0.00810892507433891,
-0.00812961161136627,
-0.00815033726394177,
-0.00817110389471054,
-0.00819191057235003,
-0.00821275729686022,
-0.00823364406824112,
-0.00825457181781530,
-0.00827553868293762,
-0.00829654652625322,
-0.00831759534776211,
-0.00833868328481913,
-0.00835981220006943,
-0.00838098209351301,
-0.00840219296514988,
-0.00842344388365746,
-0.00844473484903574,
-0.00846606679260731,
-0.00848743971437216,
-0.00850885454565287,
-0.00853030849248171,
-0.00855180434882641,
-0.00857334211468697,
-0.00859491899609566,
-0.00861653871834278,
-0.00863819848746061,
-0.00865990016609430,
-0.00868164375424385,
-0.00870342832058668,
-0.00872525386512280,
-0.00874712131917477,
-0.00876903068274260,
-0.00879098102450371,
-0.00881297234445810,
-0.00883500557392836,
-0.00885708071291447,
-0.00887919776141644,
-0.00890135578811169,
-0.00892355665564537,
-0.00894579850137234,
-0.00896808318793774,
-0.00899040885269642,
-0.00901277735829353,
-0.00903518777340651,
-0.00905764009803534,
-0.00908013526350260,
-0.00910267233848572,
-0.00912525225430727,
-0.00914787314832211,
-0.00917053688317537,
-0.00919324345886707,
-0.00921599194407463,
-0.00923878420144320,
-0.00926161929965019,
-0.00928449630737305,
-0.00930741615593433,
-0.00933037884533405,
-0.00935338437557221,
-0.00937643274664879,
-0.00939952395856381,
-0.00942265801131725,
-0.00944583490490913,
-0.00946905557066202,
-0.00949231907725334,
-0.00951562542468309,
-0.00953897554427385,
-0.00956236943602562,
-0.00958580709993839,
-0.00960928760468960,
-0.00963281095027924,
-0.00965637806802988,
-0.00967998802661896,
-0.00970364362001419,
-0.00972734205424786,
-0.00975108426064253,
-0.00977487023919821,
-0.00979869998991489,
-0.00982257351279259,
-0.00984649173915386,
-0.00987045280635357,
-0.00989445857703686,
-0.00991850811988115,
-0.00994260236620903,
-0.00996674038469791,
-0.00999092310667038,
-0.0100151496008039,
-0.0100394217297435,
-0.0100637366995215,
-0.0100880973041058,
-0.0101125016808510,
-0.0101369507610798,
-0.0101614454761148,
-0.0101859839633107,
-0.0102105671539903,
-0.0102351950481534,
-0.0102598695084453,
-0.0102845877408981,
-0.0103093506768346,
-0.0103341583162546,
-0.0103590125218034,
-0.0103839104995132,
-0.0104088550433517,
-0.0104338433593512,
-0.0104588782414794,
-0.0104839578270912,
-0.0105090830475092,
-0.0105342539027333,
-0.0105594703927636,
-0.0105847325176001,
-0.0106100402772427,
-0.0106353936716914,
-0.0106607936322689,
-0.0106862382963300,
-0.0107117295265198,
-0.0107372663915157,
-0.0107628488913178,
-0.0107884788885713,
-0.0108141535893083,
-0.0108398748561740,
-0.0108656426891685,
-0.0108914561569691,
-0.0109173161908984,
-0.0109432227909565,
-0.0109691759571433,
-0.0109951756894588,
-0.0110212210565805,
-0.0110473139211535,
-0.0110734533518553,
-0.0110996393486857,
-0.0111258728429675,
-0.0111521519720554,
-0.0111784795299172,
-0.0112048527225852,
-0.0112312734127045,
-0.0112577406689525,
-0.0112842554226518,
-0.0113108176738024,
-0.0113374264910817,
-0.0113640837371349,
-0.0113907875493169,
-0.0114175379276276,
-0.0114443367347121,
-0.0114711830392480,
-0.0114980768412352,
-0.0115250181406736,
-0.0115520078688860,
-0.0115790450945497,
-0.0116061298176646,
-0.0116332620382309,
-0.0116604417562485,
-0.0116876699030399,
-0.0117149464786053,
-0.0117422714829445,
-0.0117696439847350,
-0.0117970658466220,
-0.0118245342746377,
-0.0118520520627499,
-0.0118796182796359,
-0.0119072329252958,
-0.0119348959997296,
-0.0119626065716147,
-0.0119903665035963,
-0.0120181757956743,
-0.0120460325852036,
-0.0120739387348294,
-0.0121018942445517,
-0.0121298981830478,
-0.0121579514816403,
-0.0121860541403294,
-0.0122142052277923,
-0.0122424056753516,
-0.0122706545516849,
-0.0122989537194371,
-0.0123273013159633,
-0.0123556982725859,
-0.0123841445893049,
-0.0124126402661204,
-0.0124411853030324,
-0.0124697806313634,
-0.0124984234571457,
-0.0125271165743470,
-0.0125558590516448,
-0.0125846518203616,
-0.0126134939491749,
-0.0126423863694072,
-0.0126713290810585,
-0.0127003202214837,
-0.0127293625846505,
-0.0127584543079138,
-0.0127875963225961,
-0.0128167886286974,
-0.0128460321575403,
-0.0128753259778023,
-0.0129046700894833,
-0.0129340635612607,
-0.0129635091871023,
-0.0129930041730404,
-0.0130225503817201,
-0.0130521468818188,
-0.0130817946046591,
-0.0131114935502410,
-0.0131412427872419,
-0.0131710432469845,
-0.0132008939981461,
-0.0132307959720492,
-0.0132607501000166,
-0.0132907545194030,
-0.0133208101615310,
-0.0133509179577231,
-0.0133810760453343,
-0.0134112853556871,
-0.0134415468201041,
-0.0134718595072627,
-0.0135022243484855,
-0.0135326404124498,
-0.0135631086304784,
-0.0135936280712485,
-0.0136241996660829,
-0.0136548224836588,
-0.0136854983866215,
-0.0137162245810032,
-0.0137470038607717,
-0.0137778352946043,
-0.0138087188825011,
-0.0138396546244621,
-0.0138706415891647,
-0.0139016816392541,
-0.0139327738434076,
-0.0139639182016253,
-0.0139951156452298,
-0.0140263661742210,
-0.0140576688572764,
-0.0140890246257186,
-0.0141204325482249,
-0.0141518935561180,
-0.0141834067180753,
-0.0142149738967419,
-0.0142465941607952,
-0.0142782665789127,
-0.0143099920824170,
-0.0143417716026306,
-0.0143736042082310,
-0.0144054889678955,
-0.0144374277442694,
-0.0144694205373526,
-0.0145014664158225,
-0.0145335653796792,
-0.0145657183602452,
-0.0145979244261980,
-0.0146301835775375,
-0.0146624986082315,
-0.0146948657929897,
-0.0147272869944572,
-0.0147597631439567,
-0.0147922923788428,
-0.0148248756304383,
-0.0148575128987432,
-0.0148902051150799,
-0.0149229513481259,
-0.0149557515978813,
-0.0149886058643460,
-0.0150215150788426,
-0.0150544783100486,
-0.0150874964892864,
-0.0151205696165562,
-0.0151536967605352,
-0.0151868788525462,
-0.0152201158925891,
-0.0152534078806639,
-0.0152867548167706,
-0.0153201557695866,
-0.0153536135330796,
-0.0153871253132820,
-0.0154206920415163,
-0.0154543146491051,
-0.0154879922047257,
-0.0155217256397009,
-0.0155555130913854,
-0.0155893564224243,
-0.0156232556328177,
-0.0156572107225657,
-0.0156912207603455,
-0.0157252885401249,
-0.0157594103366137,
-0.0157935880124569,
-0.0158278215676546,
-0.0158621110022068,
-0.0158964563161135,
-0.0159308593720198,
-0.0159653164446354,
-0.0159998312592506,
-0.0160344019532204,
-0.0160690285265446,
-0.0161037128418684,
-0.0161384530365467,
-0.0161732491105795,
-0.0162081010639668,
-0.0162430107593536,
-0.0162779781967402,
-0.0163129996508360,
-0.0163480807095766,
-0.0163832176476717,
-0.0164184104651213,
-0.0164536610245705,
-0.0164889693260193,
-0.0165243353694677,
-0.0165597572922707,
-0.0165952369570732,
-0.0166307743638754,
-0.0166663695126772,
-0.0167020205408335,
-0.0167377311736345,
-0.0167734976857901,
-0.0168093219399452,
-0.0168452057987452,
-0.0168811455368996,
-0.0169171448796988,
-0.0169532001018524,
-0.0169893149286509,
-0.0170254856348038,
-0.0170617159456015,
-0.0170980039983988,
-0.0171343516558409,
-0.0171707551926374,
-0.0172072201967239,
-0.0172437410801649,
-0.0172803215682507,
-0.0173169597983360,
-0.0173536576330662,
-0.0173904150724411,
-0.0174272302538157,
-0.0174641031771898,
-0.0175010357052088,
-0.0175380259752274,
-0.0175750758498907,
-0.0176121853291988,
-0.0176493525505066,
-0.0176865831017494,
-0.0177238713949919,
-0.0177612174302340,
-0.0177986249327660,
-0.0178360901772976,
-0.0178736131638289,
-0.0179111994802952,
-0.0179488435387611,
-0.0179865472018719,
-0.0180243123322725,
-0.0180621352046728,
-0.0181000195443630,
-0.0181379634886980,
-0.0181759670376778,
-0.0182140301913023,
-0.0182521548122168,
-0.0182903390377760,
-0.0183285847306252,
-0.0183668900281191,
-0.0184052549302578,
-0.0184436831623316,
-0.0184821691364050,
-0.0185207165777683,
-0.0185593254864216,
-0.0185979958623648,
-0.0186367258429527,
-0.0186755154281855,
-0.0187143683433533,
-0.0187532808631659,
-0.0187922548502684,
-0.0188312903046608,
-0.0188703872263432,
-0.0189095456153154,
-0.0189487636089325,
-0.0189880449324846,
-0.0190273858606815,
-0.0190667901188135,
-0.0191062558442354,
-0.0191457830369473,
-0.0191853716969490,
-0.0192250218242407,
-0.0192647352814674,
-0.0193045102059841,
-0.0193443465977907,
-0.0193842463195324,
-0.0194242075085640,
-0.0194642320275307,
-0.0195043180137873,
-0.0195444673299789,
-0.0195846762508154,
-0.0196249503642321,
-0.0196652859449387,
-0.0197056848555803,
-0.0197461470961571,
-0.0197866708040237,
-0.0198272559791803,
-0.0198679063469172,
-0.0199086200445890,
-0.0199493970721960,
-0.0199902374297380,
-0.0200311392545700,
-0.0200721044093370,
-0.0201131328940392,
-0.0201542247086763,
-0.0201953817158937,
-0.0202366001904011,
-0.0202778838574886,
-0.0203192308545113,
-0.0203606411814690,
-0.0204021167010069,
-0.0204436555504799,
-0.0204852595925331,
-0.0205269251018763,
-0.0205686558037996,
-0.0206104516983032,
-0.0206523109227419,
-0.0206942353397608,
-0.0207362230867147,
-0.0207782760262489,
-0.0208203922957182,
-0.0208625756204128,
-0.0209048222750425,
-0.0209471341222525,
-0.0209895092993975,
-0.0210319496691227,
-0.0210744570940733,
-0.0211170278489590,
-0.0211596637964249,
-0.0212023649364710,
-0.0212451331317425,
-0.0212879665195942,
-0.0213308632373810,
-0.0213738251477480,
-0.0214168522506952,
-0.0214599464088678,
-0.0215031057596207,
-0.0215463321655989,
-0.0215896219015121,
-0.0216329786926508,
-0.0216764025390148,
-0.0217198915779591,
-0.0217634476721287,
-0.0218070689588785,
-0.0218507573008537,
-0.0218945108354092,
-0.0219383314251900,
-0.0219822190701962,
-0.0220261737704277,
-0.0220701936632395,
-0.0221142806112766,
-0.0221584346145391,
-0.0222026538103819,
-0.0222469419240952,
-0.0222912952303886,
-0.0223357174545527,
-0.0223802067339420,
-0.0224247612059116,
-0.0224693845957518,
-0.0225140750408173,
-0.0225588325411081,
-0.0226036570966244,
-0.0226485505700111,
-0.0226935110986233,
-0.0227385386824608,
-0.0227836351841688,
-0.0228288006037474,
-0.0228740330785513,
-0.0229193326085806,
-0.0229647010564804,
-0.0230101384222507,
-0.0230556428432465,
-0.0231012143194675,
-0.0231468547135592,
-0.0231925621628761,
-0.0232383403927088,
-0.0232841875404120,
-0.0233301017433405,
-0.0233760867267847,
-0.0234221387654543,
-0.0234682597219944,
-0.0235144495964050,
-0.0235607083886862,
-0.0236070360988379,
-0.0236534327268600,
-0.0236999001353979,
-0.0237464345991611,
-0.0237930398434401,
-0.0238397158682346,
-0.0238864589482546,
-0.0239332728087902,
-0.0239801555871964,
-0.0240271091461182,
-0.0240741316229105,
-0.0241212230175734,
-0.0241683851927519,
-0.0242156181484461,
-0.0242629200220108,
-0.0243102926760912,
-0.0243577361106873,
-0.0244052503257990,
-0.0244528297334909,
-0.0245004817843437,
-0.0245482027530670,
-0.0245959963649511,
-0.0246438588947058,
-0.0246917940676212,
-0.0247397981584072,
-0.0247878730297089,
-0.0248360205441713,
-0.0248842369765043,
-0.0249325260519981,
-0.0249808859080076,
-0.0250293184071779,
-0.0250778198242188,
-0.0251263957470655,
-0.0251750405877829,
-0.0252237562090158,
-0.0252725463360548,
-0.0253214072436094,
-0.0253703389316797,
-0.0254193432629108,
-0.0254684202373028,
-0.0255175679922104,
-0.0255667883902788,
-0.0256160795688629,
-0.0256654452532530,
-0.0257148817181587,
-0.0257643908262253,
-0.0258139725774527,
-0.0258636269718409,
-0.0259133540093899,
-0.0259631536900997,
-0.0260130260139704,
-0.0260629728436470,
-0.0261129904538393,
-0.0261630825698376,
-0.0262132454663515,
-0.0262634847313166,
-0.0263137947767973,
-0.0263641793280840,
-0.0264146365225315,
-0.0264651663601398,
-0.0265157725661993,
-0.0265664495527744,
-0.0266172029078007,
-0.0266680270433426,
-0.0267189256846905,
-0.0267699006944895,
-0.0268209464848042,
-0.0268720686435699,
-0.0269232634454966,
-0.0269745346158743,
-0.0270258784294128,
-0.0270772948861122,
-0.0271287877112627,
-0.0271803550422192,
-0.0272319968789816,
-0.0272837132215500,
-0.0273355040699244,
-0.0273873712867498,
-0.0274393111467361,
-0.0274913273751736,
-0.0275434181094170,
-0.0275955852121115,
-0.0276478268206120,
-0.0277001429349184,
-0.0277525372803211,
-0.0278050042688847,
-0.0278575476258993,
-0.0279101673513651,
-0.0279628615826368,
-0.0280156321823597,
-0.0280684791505337,
-0.0281214006245136,
-0.0281743984669447,
-0.0282274726778269,
-0.0282806251198053,
-0.0283338502049446,
-0.0283871535211802,
-0.0284405332058668,
-0.0284939892590046,
-0.0285475198179483,
-0.0286011286079884,
-0.0286548156291246,
-0.0287085771560669,
-0.0287624169141054,
-0.0288163330405951,
-0.0288703273981810,
-0.0289243962615728,
-0.0289785452187061,
-0.0290327686816454,
-0.0290870703756809,
-0.0291414503008127,
-0.0291959084570408,
-0.0292504429817200,
-0.0293050538748503,
-0.0293597448617220,
-0.0294145122170448,
-0.0294693578034639,
-0.0295242816209793,
-0.0295792818069458,
-0.0296343620866537,
-0.0296895205974579,
-0.0297447573393583,
-0.0298000723123550,
-0.0298554636538029,
-0.0299109350889921,
-0.0299664866179228,
-0.0300221163779497,
-0.0300778225064278,
-0.0301336087286472,
-0.0301894731819630,
-0.0302454177290201,
-0.0303014423698187,
-0.0303575433790684,
-0.0304137263447046,
-0.0304699875414372,
-0.0305263269692659,
-0.0305827464908361,
-0.0306392461061478,
-0.0306958239525557,
-0.0307524818927050,
-0.0308092199265957,
-0.0308660380542278,
-0.0309229362756014,
-0.0309799145907164,
-0.0310369729995728,
-0.0310941096395254,
-0.0311513282358646,
-0.0312086269259453,
-0.0312660038471222,
-0.0313234627246857,
-0.0313810035586357,
-0.0314386226236820,
-0.0314963236451149,
-0.0315541066229343,
-0.0316119715571404,
-0.0316699147224426,
-0.0317279398441315,
-0.0317860431969166,
-0.0318442322313786,
-0.0319024994969368,
-0.0319608524441719,
-0.0320192836225033,
-0.0320777967572212,
-0.0321363918483257,
-0.0321950688958168,
-0.0322538241744041,
-0.0323126651346684,
-0.0323715843260288,
-0.0324305891990662,
-0.0324896723031998,
-0.0325488410890102,
-0.0326080881059170,
-0.0326674208045006,
-0.0327268354594708,
-0.0327863283455372,
-0.0328459106385708,
-0.0329055711627007,
-0.0329653136432171,
-0.0330251418054104,
-0.0330850519239903,
-0.0331450439989567,
-0.0332051180303097,
-0.0332652777433395,
-0.0333255194127560,
-0.0333858430385590,
-0.0334462523460388,
-0.0335067436099052,
-0.0335673205554485,
-0.0336279757320881,
-0.0336887203156948,
-0.0337495431303978,
-0.0338104516267777,
-0.0338714458048344,
-0.0339325219392777,
-0.0339936800301075,
-0.0340549275279045,
-0.0341162569820881,
-0.0341776721179485,
-0.0342391692101955,
-0.0343007519841194,
-0.0343624167144299,
-0.0344241671264172,
-0.0344860032200813,
-0.0345479249954224,
-0.0346099287271500,
-0.0346720181405544,
-0.0347341969609261,
-0.0347964540123940,
-0.0348588004708290,
-0.0349212288856506,
-0.0349837467074394,
-0.0350463464856148,
-0.0351090356707573,
-0.0351718068122864,
-0.0352346636354923,
-0.0352976061403751,
-0.0353606343269348,
-0.0354237481951714,
-0.0354869477450848,
-0.0355502367019653,
-0.0356136076152325,
-0.0356770679354668,
-0.0357406102120876,
-0.0358042418956757,
-0.0358679592609406,
-0.0359317623078823,
-0.0359956510365009,
-0.0360596291720867,
-0.0361236967146397,
-0.0361878499388695,
-0.0362520851194859,
-0.0363164097070694,
-0.0363808162510395,
-0.0364453122019768,
-0.0365098938345909,
-0.0365745648741722,
-0.0366393178701401,
-0.0367041639983654,
-0.0367690958082676,
-0.0368341132998467,
-0.0368992201983929,
-0.0369644165039063,
-0.0370296984910965,
-0.0370950661599636,
-0.0371605232357979,
-0.0372260734438896,
-0.0372917056083679,
-0.0373574309051037,
-0.0374232418835163,
-0.0374891422688961,
-0.0375551283359528,
-0.0376212075352669,
-0.0376873724162579,
-0.0377536267042160,
-0.0378199666738510,
-0.0378863960504532,
-0.0379529185593128,
-0.0380195267498493,
-0.0380862243473530,
-0.0381530150771141,
-0.0382198914885521,
-0.0382868573069572,
-0.0383539125323296,
-0.0384210608899593,
-0.0384882912039757,
-0.0385556146502495,
-0.0386230312287807,
-0.0386905372142792,
-0.0387581326067448,
-0.0388258174061775,
-0.0388935916125774,
-0.0389614552259445,
-0.0390294082462788,
-0.0390974506735802,
-0.0391655862331390,
-0.0392338149249554,
-0.0393021292984486,
-0.0393705368041992,
-0.0394390337169170,
-0.0395076237618923,
-0.0395763032138348,
-0.0396450720727444,
-0.0397139340639114,
-0.0397828891873360,
-0.0398519337177277,
-0.0399210713803768,
-0.0399902984499931,
-0.0400596149265766,
-0.0401290245354176,
-0.0401985272765160,
-0.0402681231498718,
-0.0403378084301949,
-0.0404075905680656,
-0.0404774621129036,
-0.0405474230647087,
-0.0406174734234810,
-0.0406876243650913,
-0.0407578609883785,
-0.0408281944692135,
-0.0408986173570156,
-0.0409691333770752,
-0.0410397425293922,
-0.0411104448139668,
-0.0411812402307987,
-0.0412521287798882,
-0.0413231104612350,
-0.0413941815495491,
-0.0414653494954109,
-0.0415366142988205,
-0.0416079685091972,
-0.0416794158518314,
-0.0417509563267231,
-0.0418225899338722,
-0.0418943203985691,
-0.0419661402702332,
-0.0420380569994450,
-0.0421100705862045,
-0.0421821773052216,
-0.0422543734312058,
-0.0423266664147377,
-0.0423990525305271,
-0.0424715355038643,
-0.0425441153347492,
-0.0426167882978916,
-0.0426895506680012,
-0.0427624098956585,
-0.0428353659808636,
-0.0429084151983261,
-0.0429815612733364,
-0.0430548004806042,
-0.0431281365454197,
-0.0432015657424927,
-0.0432750955224037,
-0.0433487147092819,
-0.0434224307537079,
-0.0434962436556816,
-0.0435701496899128,
-0.0436441563069820,
-0.0437182597815990,
-0.0437924563884735,
-0.0438667498528957,
-0.0439411364495754,
-0.0440156199038029,
-0.0440902039408684,
-0.0441648811101913,
-0.0442396551370621,
-0.0443145260214806,
-0.0443894937634468,
-0.0444645583629608,
-0.0445397160947323,
-0.0446149781346321,
-0.0446903295814991,
-0.0447657853364944,
-0.0448413342237473,
-0.0449169799685478,
-0.0449927262961865,
-0.0450685657560825,
-0.0451445057988167,
-0.0452205389738083,
-0.0452966727316380,
-0.0453729070723057,
-0.0454492382705212,
-0.0455256700515747,
-0.0456021949648857,
-0.0456788204610348,
-0.0457555428147316,
-0.0458323620259762,
-0.0459092818200588,
-0.0459863021969795,
-0.0460634194314480,
-0.0461406335234642,
-0.0462179481983185,
-0.0462953634560108,
-0.0463728718459606,
-0.0464504845440388,
-0.0465281940996647,
-0.0466060042381287,
-0.0466839112341404,
-0.0467619225382805,
-0.0468400306999683,
-0.0469182394444943,
-0.0469965487718582,
-0.0470749586820602,
-0.0471534617245197,
-0.0472320690751076,
-0.0473107770085335,
-0.0473895855247974,
-0.0474684946238995,
-0.0475475005805492,
-0.0476266108453274,
-0.0477058179676533,
-0.0477851256728172,
-0.0478645339608192,
-0.0479440465569496,
-0.0480236560106278,
-0.0481033697724342,
-0.0481831803917885,
-0.0482630953192711,
-0.0483431033790112,
-0.0484232157468796,
-0.0485034249722958,
-0.0485837422311306,
-0.0486641563475132,
-0.0487446710467339,
-0.0488252900540829,
-0.0489060096442699,
-0.0489868335425854,
-0.0490677580237389,
-0.0491487868130207,
-0.0492299124598503,
-0.0493111461400986,
-0.0493924766778946,
-0.0494739152491093,
-0.0495554506778717,
-0.0496370941400528,
-0.0497188381850719,
-0.0498006828129292,
-0.0498826354742050,
-0.0499646887183189,
-0.0500468425452709,
-0.0501291006803513,
-0.0502114631235600,
-0.0502939336001873,
-0.0503765009343624,
-0.0504591725766659,
-0.0505419485270977,
-0.0506248287856579,
-0.0507078133523464,
-0.0507909059524536,
-0.0508740954101086,
-0.0509573891758919,
-0.0510407872498035,
-0.0511242933571339,
-0.0512079000473022,
-0.0512916110455990,
-0.0513754300773144,
-0.0514593496918678,
-0.0515433773398399,
-0.0516275130212307,
-0.0517117530107498,
-0.0517960935831070,
-0.0518805421888828,
-0.0519650951027870,
-0.0520497523248196,
-0.0521345175802708,
-0.0522193871438503,
-0.0523043610155582,
-0.0523894429206848,
-0.0524746328592300,
-0.0525599233806133,
-0.0526453219354153,
-0.0527308285236359,
-0.0528164431452751,
-0.0529021583497524,
-0.0529879815876484,
-0.0530739128589630,
-0.0531599521636963,
-0.0532460957765579,
-0.0533323474228382,
-0.0534187033772469,
-0.0535051710903645,
-0.0535917431116104,
-0.0536784194409847,
-0.0537652038037777,
-0.0538520999252796,
-0.0539391003549099,
-0.0540262088179588,
-0.0541134253144264,
-0.0542007498443127,
-0.0542881786823273,
-0.0543757192790508,
-0.0544633679091930,
-0.0545511245727539,
-0.0546389855444431,
-0.0547269545495510,
-0.0548150353133678,
-0.0549032241106033,
-0.0549915209412575,
-0.0550799295306206,
-0.0551684461534023,
-0.0552570670843124,
-0.0553457960486412,
-0.0554346367716789,
-0.0555235855281353,
-0.0556126423180103,
-0.0557018108665943,
-0.0557910911738873,
-0.0558804795145988,
-0.0559699796140194,
-0.0560595877468586,
-0.0561493039131165,
-0.0562391281127930,
-0.0563290640711784,
-0.0564191117882729,
-0.0565092712640762,
-0.0565995387732983,
-0.0566899143159390,
-0.0567804053425789,
-0.0568710044026375,
-0.0569617114961147,
-0.0570525340735912,
-0.0571434646844864,
-0.0572345070540905,
-0.0573256611824036,
-0.0574169233441353,
-0.0575083009898663,
-0.0575997866690159,
-0.0576913878321648,
-0.0577830970287323,
-0.0578749217092991,
-0.0579668544232845,
-0.0580588988959789,
-0.0581510551273823,
-0.0582433231174946,
-0.0583357065916061,
-0.0584281980991364,
-0.0585208050906658,
-0.0586135238409042,
-0.0587063506245613,
-0.0587992928922176,
-0.0588923506438732,
-0.0589855201542378,
-0.0590788051486015,
-0.0591721981763840,
-0.0592657029628754,
-0.0593593232333660,
-0.0594530589878559,
-0.0595469065010548,
-0.0596408694982529,
-0.0597349442541599,
-0.0598291344940662,
-0.0599234364926815,
-0.0600178539752960,
-0.0601123832166195,
-0.0602070279419422,
-0.0603017807006836,
-0.0603966489434242,
-0.0604916252195835,
-0.0605867207050324,
-0.0606819316744804,
-0.0607772581279278,
-0.0608726963400841,
-0.0609682500362396,
-0.0610639154911041,
-0.0611597001552582,
-0.0612556003034115,
-0.0613516122102737,
-0.0614477433264256,
-0.0615439899265766,
-0.0616403482854366,
-0.0617368258535862,
-0.0618334189057350,
-0.0619301274418831,
-0.0620269514620304,
-0.0621238909661770,
-0.0622209459543228,
-0.0623181201517582,
-0.0624154098331928,
-0.0625128149986267,
-0.0626103356480598,
-0.0627079755067825,
-0.0628057271242142,
-0.0629035979509354,
-0.0630015879869461,
-0.0630996972322464,
-0.0631979182362557,
-0.0632962584495544,
-0.0633947178721428,
-0.0634932965040207,
-0.0635919868946075,
-0.0636907964944840,
-0.0637897253036499,
-0.0638887733221054,
-0.0639879330992699,
-0.0640872195363045,
-0.0641866177320480,
-0.0642861351370812,
-0.0643857717514038,
-0.0644855350255966,
-0.0645854100584984,
-0.0646853968501091,
-0.0647855103015900,
-0.0648857429623604,
-0.0649860873818398,
-0.0650865584611893,
-0.0651871412992477,
-0.0652878507971764,
-0.0653886795043945,
-0.0654896274209023,
-0.0655906870961189,
-0.0656918734312058,
-0.0657931789755821,
-0.0658946037292481,
-0.0659961551427841,
-0.0660978183150291,
-0.0661996006965637,
-0.0663015097379684,
-0.0664035379886627,
-0.0665056854486466,
-0.0666079521179199,
-0.0667103379964829,
-0.0668128505349159,
-0.0669154822826386,
-0.0670182332396507,
-0.0671211034059525,
-0.0672240927815437,
-0.0673272088170052,
-0.0674304515123367,
-0.0675338059663773,
-0.0676372870802879,
-0.0677408874034882,
-0.0678446069359779,
-0.0679484531283379,
-0.0680524185299873,
-0.0681565105915070,
-0.0682607293128967,
-0.0683650597929955,
-0.0684695169329643,
-0.0685740932822228,
-0.0686787962913513,
-0.0687836185097694,
-0.0688885673880577,
-0.0689936354756355,
-0.0690988302230835,
-0.0692041516304016,
-0.0693095922470093,
-0.0694151520729065,
-0.0695208460092545,
-0.0696266517043114,
-0.0697325840592384,
-0.0698386430740356,
-0.0699448212981224,
-0.0700511261820793,
-0.0701575577259064,
-0.0702641159296036,
-0.0703708007931709,
-0.0704776048660278,
-0.0705845281481743,
-0.0706915780901909,
-0.0707987546920776,
-0.0709060579538345,
-0.0710134878754616,
-0.0711210444569588,
-0.0712287202477455,
-0.0713365152478218,
-0.0714444443583489,
-0.0715525001287460,
-0.0716606825590134,
-0.0717689916491509,
-0.0718774199485779,
-0.0719859749078751,
-0.0720946565270424,
-0.0722034648060799,
-0.0723123922944069,
-0.0724214389920235,
-0.0725306198000908,
-0.0726399272680283,
-0.0727493613958359,
-0.0728589221835136,
-0.0729686021804810,
-0.0730784237384796,
-0.0731883645057678,
-0.0732984319329262,
-0.0734086334705353,
-0.0735189542174339,
-0.0736294016242027,
-0.0737399756908417,
-0.0738506838679314,
-0.0739615187048912,
-0.0740724802017212,
-0.0741835609078407,
-0.0742947831749916,
-0.0744061246514320,
-0.0745176002383232,
-0.0746292024850845,
-0.0747409388422966,
-0.0748527944087982,
-0.0749647840857506,
-0.0750769004225731,
-0.0751891508698463,
-0.0753015279769898,
-0.0754140317440033,
-0.0755266696214676,
-0.0756394267082214,
-0.0757523253560066,
-0.0758653506636620,
-0.0759785026311874,
-0.0760917812585831,
-0.0762051939964294,
-0.0763187333941460,
-0.0764324069023132,
-0.0765462070703507,
-0.0766601413488388,
-0.0767742097377777,
-0.0768884047865868,
-0.0770027264952660,
-0.0771171823143959,
-0.0772317722439766,
-0.0773464962840080,
-0.0774613395333290,
-0.0775763168931007,
-0.0776914209127426,
-0.0778066664934158,
-0.0779220387339592,
-0.0780375450849533,
-0.0781531855463982,
-0.0782689601182938,
-0.0783848613500595,
-0.0785008966922760,
-0.0786170661449432,
-0.0787333697080612,
-0.0788498073816299,
-0.0789663717150688,
-0.0790830701589584,
-0.0791999027132988,
-0.0793168693780899,
-0.0794339627027512,
-0.0795511901378632,
-0.0796685516834259,
-0.0797860473394394,
-0.0799036771059036,
-0.0800214335322380,
-0.0801393315196037,
-0.0802573561668396,
-0.0803755149245262,
-0.0804938152432442,
-0.0806122422218323,
-0.0807308107614517,
-0.0808495059609413,
-0.0809683352708817,
-0.0810873061418533,
-0.0812064111232758,
-0.0813256502151489,
-0.0814450159668922,
-0.0815645232796669,
-0.0816841721534729,
-0.0818039476871491,
-0.0819238573312759,
-0.0820439085364342,
-0.0821640864014626,
-0.0822844058275223,
-0.0824048593640328,
-0.0825254544615746,
-0.0826461762189865,
-0.0827670395374298,
-0.0828880369663239,
-0.0830091685056686,
-0.0831304416060448,
-0.0832518413662911,
-0.0833733901381493,
-0.0834950655698776,
-0.0836168900132179,
-0.0837388411164284,
-0.0838609337806702,
-0.0839831605553627,
-0.0841055139899254,
-0.0842280089855194,
-0.0843506455421448,
-0.0844734087586403,
-0.0845963209867477,
-0.0847193673253059,
-0.0848425477743149,
-0.0849658623337746,
-0.0850893259048462,
-0.0852129161357880,
-0.0853366479277611,
-0.0854605212807655,
-0.0855845287442207,
-0.0857086777687073,
-0.0858329758048058,
-0.0859574005007744,
-0.0860819667577744,
-0.0862066745758057,
-0.0863315090537071,
-0.0864564925432205,
-0.0865816175937653,
-0.0867068842053413,
-0.0868322849273682,
-0.0869578272104263,
-0.0870835110545158,
-0.0872093364596367,
-0.0873352885246277,
-0.0874613896012306,
-0.0875876322388649,
-0.0877140164375305,
-0.0878405421972275,
-0.0879672095179558,
-0.0880940183997154,
-0.0882209613919258,
-0.0883480459451675,
-0.0884752720594406,
-0.0886026397347450,
-0.0887301489710808,
-0.0888577997684479,
-0.0889855921268463,
-0.0891135260462761,
-0.0892416015267372,
-0.0893698260188103,
-0.0894981846213341,
-0.0896266922354698,
-0.0897553339600563,
-0.0898841246962547,
-0.0900130495429039,
-0.0901421234011650,
-0.0902713388204575,
-0.0904006958007813,
-0.0905301943421364,
-0.0906598269939423,
-0.0907896235585213,
-0.0909195542335510,
-0.0910496264696121,
-0.0911798477172852,
-0.0913102030754089,
-0.0914407074451447,
-0.0915713533759117,
-0.0917021483182907,
-0.0918330848217011,
-0.0919641628861427,
-0.0920953899621964,
-0.0922267585992813,
-0.0923582687973976,
-0.0924899280071259,
-0.0926217362284660,
-0.0927536860108376,
-0.0928857773542404,
-0.0930180102586746,
-0.0931503921747208,
-0.0932829156517983,
-0.0934155955910683,
-0.0935484170913696,
-0.0936813801527023,
-0.0938144922256470,
-0.0939477458596230,
-0.0940811559557915,
-0.0942147001624107,
-0.0943483933806419,
-0.0944822356104851,
-0.0946162194013596,
-0.0947503596544266,
-0.0948846340179443,
-0.0950190648436546,
-0.0951536372303963,
-0.0952883586287499,
-0.0954232215881348,
-0.0955582410097122,
-0.0956934094429016,
-0.0958287194371223,
-0.0959641784429550,
-0.0960997715592384,
-0.0962355136871338,
-0.0963714122772217,
-0.0965074449777603,
-0.0966436341404915,
-0.0967799797654152,
-0.0969164595007896,
-0.0970530956983566,
-0.0971898809075356,
-0.0973268076777458,
-0.0974638909101486,
-0.0976011157035828,
-0.0977384969592094,
-0.0978760197758675,
-0.0980136990547180,
-0.0981515273451805,
-0.0982895046472549,
-0.0984276235103607,
-0.0985658988356590,
-0.0987043231725693,
-0.0988428965210915,
-0.0989816188812256,
-0.0991204977035523,
-0.0992595255374908,
-0.0993987023830414,
-0.0995380207896233,
-0.0996774956583977,
-0.0998171195387840,
-0.0999568998813629,
-0.100096829235554,
-0.100236907601357,
-0.100377142429352,
-0.100517526268959,
-0.100658059120178,
-0.100798740983009,
-0.100939579308033,
-0.101080574095249,
-0.101221710443497,
-0.101363003253937,
-0.101504445075989,
-0.101646043360233,
-0.101787798106670,
-0.101929709315300,
-0.102071762084961,
-0.102213971316814,
-0.102356337010860,
-0.102498851716518,
-0.102641515433788,
-0.102784343063831,
-0.102927319705486,
-0.103070445358753,
-0.103213727474213,
-0.103357158601284,
-0.103500753641129,
-0.103644497692585,
-0.103788390755653,
-0.103932447731495,
-0.104076661169529,
-0.104221016168594,
-0.104365535080433,
-0.104510210454464,
-0.104655034840107,
-0.104800015687943,
-0.104945152997971,
-0.105090446770191,
-0.105235889554024,
-0.105381488800049,
-0.105527251958847,
-0.105673164129257,
-0.105819232761860,
-0.105965457856655,
-0.106111831963062,
-0.106258369982243,
-0.106405064463615,
-0.106551915407181,
-0.106698915362358,
-0.106846079230309,
-0.106993392109871,
-0.107140868902206,
-0.107288502156734,
-0.107436291873455,
-0.107584245502949,
-0.107732340693474,
-0.107880607247353,
-0.108029015362263,
-0.108177579939365,
-0.108326300978661,
-0.108475185930729,
-0.108624227344990,
-0.108773425221443,
-0.108922779560089,
-0.109072290360928,
-0.109221957623959,
-0.109371796250343,
-0.109521783888340,
-0.109671927988529,
-0.109822236001492,
-0.109972700476646,
-0.110123328864574,
-0.110274121165276,
-0.110425062477589,
-0.110576160252094,
-0.110727421939373,
-0.110878847539425,
-0.111030429601669,
-0.111182175576687,
-0.111334078013897,
-0.111486144363880,
-0.111638374626637,
-0.111790753901005,
-0.111943297088146,
-0.112095996737480,
-0.112248860299587,
-0.112401887774467,
-0.112555071711540,
-0.112708419561386,
-0.112861931324005,
-0.113015606999397,
-0.113169446587563,
-0.113323442637920,
-0.113477602601051,
-0.113631926476955,
-0.113786406815052,
-0.113941051065922,
-0.114095859229565,
-0.114250823855400,
-0.114405952394009,
-0.114561252295971,
-0.114716708660126,
-0.114872328937054,
-0.115028113126755,
-0.115184053778648,
-0.115340165793896,
-0.115496441721916,
-0.115652874112129,
-0.115809470415115,
-0.115966238081455,
-0.116123162209988,
-0.116280250251293,
-0.116437509655952,
-0.116594932973385,
-0.116752512753010,
-0.116910263895988,
-0.117068178951740,
-0.117226250469685,
-0.117384500801563,
-0.117542907595634,
-0.117701478302479,
-0.117860220372677,
-0.118019118905067,
-0.118178188800812,
-0.118337415158749,
-0.118496820330620,
-0.118656381964684,
-0.118816114962101,
-0.118976011872292,
-0.119136072695255,
-0.119296297430992,
-0.119456693530083,
-0.119617260992527,
-0.119777992367744,
-0.119938880205154,
-0.120099924504757,
-0.120261140167713,
-0.120422534644604,
-0.120584078133106,
-0.120745800435543,
-0.120907694101334,
-0.121069744229317,
-0.121231965720654,
-0.121394358575344,
-0.121556915342808,
-0.121719636023045,
-0.121882535517216,
-0.122045598924160,
-0.122208826243877,
-0.122372224926949,
-0.122535794973373,
-0.122699536383152,
-0.122863441705704,
-0.123027525842190,
-0.123191766440868,
-0.123356178402901,
-0.123520761728287,
-0.123685516417027,
-0.123850435018539,
-0.124015532433987,
-0.124180801212788,
-0.124346233904362,
-0.124511837959290,
-0.124677620828152,
-0.124843567609787,
-0.125009685754776,
-0.125175967812538,
-0.125342428684235,
-0.125509068369865,
-0.125675857067108,
-0.125842839479446,
-0.126009970903397,
-0.126177296042442,
-0.126344770193100,
-0.126512423157692,
-0.126680254936218,
-0.126848250627518,
-0.127016425132751,
-0.127184763550758,
-0.127353280782700,
-0.127521976828575,
-0.127690836787224,
-0.127859860658646,
-0.128029078245163,
-0.128198459744453,
-0.128368005156517,
-0.128537729382515,
-0.128707632422447,
-0.128877699375153,
-0.129047945141792,
-0.129218369722366,
-0.129388973116875,
-0.129559725522995,
-0.129730671644211,
-0.129901796579361,
-0.130073085427284,
-0.130244553089142,
-0.130416184663773,
-0.130588009953499,
-0.130759999155998,
-0.130932152271271,
-0.131104499101639,
-0.131277009844780,
-0.131449699401855,
-0.131622567772865,
-0.131795600056648,
-0.131968796253204,
-0.132142186164856,
-0.132315739989281,
-0.132489457726479,
-0.132663369178772,
-0.132837459445000,
-0.133011713624001,
-0.133186146616936,
-0.133360758423805,
-0.133535549044609,
-0.133710518479347,
-0.133885666728020,
-0.134060993790627,
-0.134236484766006,
-0.134412154555321,
-0.134588018059731,
-0.134764045476913,
-0.134940251708031,
-0.135116636753082,
-0.135293215513229,
-0.135469958186150,
-0.135646879673004,
-0.135823979973793,
-0.136001259088516,
-0.136178717017174,
-0.136356353759766,
-0.136534169316292,
-0.136712163686752,
-0.136890336871147,
-0.137068688869476,
-0.137247219681740,
-0.137425929307938,
-0.137604817748070,
-0.137783885002136,
-0.137963145971298,
-0.138142570853233,
-0.138322189450264,
-0.138501986861229,
-0.138681963086128,
-0.138862118124962,
-0.139042451977730,
-0.139222964644432,
-0.139403656125069,
-0.139584526419640,
-0.139765590429306,
-0.139946833252907,
-0.140128254890442,
-0.140309855341911,
-0.140491649508476,
-0.140673607587814,
-0.140855759382248,
-0.141038089990616,
-0.141220614314079,
-0.141403302550316,
-0.141586184501648,
-0.141769260168076,
-0.141952499747276,
-0.142135933041573,
-0.142319545149803,
-0.142503336071968,
-0.142687305808067,
-0.142871469259262,
-0.143055826425552,
-0.143240347504616,
-0.143425062298775,
-0.143609955906868,
-0.143795013427734,
-0.143980279564857,
-0.144165709614754,
-0.144351333379745,
-0.144537121057510,
-0.144723117351532,
-0.144909292459488,
-0.145095661282539,
-0.145282194018364,
-0.145468935370445,
-0.145655855536461,
-0.145842954516411,
-0.146030232310295,
-0.146217703819275,
-0.146405369043350,
-0.146593213081360,
-0.146781221032143,
-0.146969452500343,
-0.147157847881317,
-0.147346422076225,
-0.147535204887390,
-0.147724166512489,
-0.147913306951523,
-0.148102641105652,
-0.148292168974876,
-0.148481875658035,
-0.148671776056290,
-0.148861855268478,
-0.149052128195763,
-0.149242594838142,
-0.149433240294456,
-0.149624079465866,
-0.149815097451210,
-0.150006324052811,
-0.150197714567184,
-0.150389298796654,
-0.150581091642380,
-0.150773048400879,
-0.150965213775635,
-0.151157557964325,
-0.151350095868111,
-0.151542812585831,
-0.151735737919807,
-0.151928842067719,
-0.152122139930725,
-0.152315616607666,
-0.152509301900864,
-0.152703166007996,
-0.152897223830223,
-0.153091475367546,
-0.153285920619965,
-0.153480529785156,
-0.153675362467766,
-0.153870359063149,
-0.154065564274788,
-0.154260948300362,
-0.154456526041031,
-0.154652312397957,
-0.154848277568817,
-0.155044436454773,
-0.155240789055824,
-0.155437320470810,
-0.155634060502052,
-0.155830979347229,
-0.156028077006340,
-0.156225368380547,
-0.156422853469849,
-0.156620547175407,
-0.156818404793739,
-0.157016471028328,
-0.157214745879173,
-0.157413184642792,
-0.157611832022667,
-0.157810673117638,
-0.158009707927704,
-0.158208936452866,
-0.158408358693123,
-0.158607974648476,
-0.158807784318924,
-0.159007787704468,
-0.159207999706268,
-0.159408390522003,
-0.159608975052834,
-0.159809753298759,
-0.160010740160942,
-0.160211905837059,
-0.160413265228271,
-0.160614833235741,
-0.160816594958305,
-0.161018565297127,
-0.161220714449883,
-0.161423057317734,
-0.161625593900681,
-0.161828339099884,
-0.162031292915344,
-0.162234410643578,
-0.162437736988068,
-0.162641257047653,
-0.162844985723495,
-0.163048908114433,
-0.163253039121628,
-0.163457348942757,
-0.163661852478981,
-0.163866564631462,
-0.164071470499039,
-0.164276570081711,
-0.164481878280640,
-0.164687380194664,
-0.164893075823784,
-0.165098980069160,
-0.165305078029633,
-0.165511384606361,
-0.165717884898186,
-0.165924564003944,
-0.166131451725960,
-0.166338533163071,
-0.166545823216438,
-0.166753306984901,
-0.166960984468460,
-0.167168870568275,
-0.167376950383186,
-0.167585223913193,
-0.167793691158295,
-0.168002352118492,
-0.168211221694946,
-0.168420284986496,
-0.168629541993141,
-0.168839022517204,
-0.169048711657524,
-0.169258594512939,
-0.169468671083450,
-0.169678956270218,
-0.169889435172081,
-0.170100107789040,
-0.170310989022255,
-0.170522078871727,
-0.170733347535133,
-0.170944839715958,
-0.171156510710716,
-0.171368420124054,
-0.171580508351326,
-0.171792805194855,
-0.172005310654640,
-0.172218009829521,
-0.172430902719498,
-0.172644004225731,
-0.172857329249382,
-0.173070847988129,
-0.173284560441971,
-0.173498481512070,
-0.173712596297264,
-0.173926934599876,
-0.174141466617584,
-0.174356207251549,
-0.174571141600609,
-0.174786299467087,
-0.175001651048660,
-0.175217196345329,
-0.175432950258255,
-0.175648927688599,
-0.175865098834038,
-0.176081478595734,
-0.176298052072525,
-0.176514849066734,
-0.176731839776039,
-0.176949024200439,
-0.177166447043419,
-0.177384048700333,
-0.177601873874664,
-0.177819892764092,
-0.178038135170937,
-0.178256556391716,
-0.178475216031075,
-0.178694054484367,
-0.178913116455078,
-0.179132387042046,
-0.179351851344109,
-0.179571494460106,
-0.179791375994682,
-0.180011436343193,
-0.180231735110283,
-0.180452212691307,
-0.180672913789749,
-0.180893823504448,
-0.181114926934242,
-0.181336253881454,
-0.181557789444923,
-0.181779533624649,
-0.182001471519470,
-0.182223647832870,
-0.182446002960205,
-0.182668581604958,
-0.182891353964806,
-0.183114349842072,
-0.183337554335594,
-0.183560952544212,
-0.183784574270248,
-0.184008419513702,
-0.184232473373413,
-0.184456735849381,
-0.184681192040443,
-0.184905871748924,
-0.185130760073662,
-0.185355857014656,
-0.185581162571907,
-0.185806676745415,
-0.186032414436340,
-0.186258360743523,
-0.186484515666962,
-0.186710879206657,
-0.186937451362610,
-0.187164247035980,
-0.187391251325607,
-0.187618464231491,
-0.187845885753632,
-0.188073530793190,
-0.188301384449005,
-0.188529446721077,
-0.188757717609406,
-0.188986212015152,
-0.189214900135994,
-0.189443826675415,
-0.189672961831093,
-0.189902290701866,
-0.190131843090057,
-0.190361618995667,
-0.190591603517532,
-0.190821796655655,
-0.191052213311195,
-0.191282853484154,
-0.191513672471046,
-0.191744714975357,
-0.191975966095924,
-0.192207425832748,
-0.192439123988152,
-0.192671015858650,
-0.192903116345406,
-0.193135440349579,
-0.193367987871170,
-0.193600758910179,
-0.193833723664284,
-0.194066911935806,
-0.194300323724747,
-0.194533944129944,
-0.194767788052559,
-0.195001855492592,
-0.195236116647720,
-0.195470601320267,
-0.195705309510231,
-0.195940226316452,
-0.196175381541252,
-0.196410730481148,
-0.196646317839623,
-0.196882113814354,
-0.197118133306503,
-0.197354361414909,
-0.197590798139572,
-0.197827458381653,
-0.198064342141151,
-0.198301434516907,
-0.198538750410080,
-0.198776289820671,
-0.199014052748680,
-0.199252024292946,
-0.199490219354630,
-0.199728637933731,
-0.199967280030251,
-0.200206130743027,
-0.200445204973221,
-0.200684502720833,
-0.200924009084702,
-0.201163753867149,
-0.201403707265854,
-0.201643869280815,
-0.201884269714355,
-0.202124878764153,
-0.202365711331368,
-0.202606767416000,
-0.202848047018051,
-0.203089565038681,
-0.203331291675568,
-0.203573212027550,
-0.203815355896950,
-0.204057723283768,
-0.204300314188004,
-0.204543113708496,
-0.204786151647568,
-0.205029413104057,
-0.205272898077965,
-0.205516591668129,
-0.205760523676872,
-0.206004664301872,
-0.206249028444290,
-0.206493616104126,
-0.206738442182541,
-0.206983476877213,
-0.207228735089302,
-0.207474216818810,
-0.207719936966896,
-0.207965880632401,
-0.208212032914162,
-0.208458408713341,
-0.208705022931099,
-0.208951860666275,
-0.209198921918869,
-0.209446191787720,
-0.209693714976311,
-0.209941446781158,
-0.210189402103424,
-0.210437580943108,
-0.210685998201370,
-0.210934624075890,
-0.211183488368988,
-0.211432576179504,
-0.211681887507439,
-0.211931407451630,
-0.212181180715561,
-0.212431177496910,
-0.212681397795677,
-0.212931841611862,
-0.213182508945465,
-0.213433414697647,
-0.213684543967247,
-0.213935896754265,
-0.214187473058701,
-0.214439287781715,
-0.214691326022148,
-0.214943587779999,
-0.215196087956429,
-0.215448796749115,
-0.215701714158058,
-0.215954869985580,
-0.216208249330521,
-0.216461867094040,
-0.216715708374977,
-0.216969773173332,
-0.217224076390266,
-0.217478603124619,
-0.217733368277550,
-0.217988356947899,
-0.218243569135666,
-0.218499019742012,
-0.218754693865776,
-0.219010606408119,
-0.219266757369041,
-0.219523131847382,
-0.219779744744301,
-0.220036566257477,
-0.220293641090393,
-0.220550924539566,
-0.220808461308479,
-0.221066221594810,
-0.221324205398560,
-0.221582427620888,
-0.221840873360634,
-0.222099557518959,
-0.222358494997025,
-0.222617626190186,
-0.222877010703087,
-0.223136633634567,
-0.223396480083466,
-0.223656564950943,
-0.223916873335838,
-0.224177420139313,
-0.224438205361366,
-0.224699214100838,
-0.224960461258888,
-0.225221931934357,
-0.225483655929565,
-0.225745603442192,
-0.226007789373398,
-0.226270198822021,
-0.226532861590385,
-0.226795747876167,
-0.227058857679367,
-0.227322190999985,
-0.227585762739182,
-0.227849572896957,
-0.228113621473312,
-0.228377878665924,
-0.228642389178276,
-0.228907138109207,
-0.229172125458717,
-0.229437351226807,
-0.229702800512314,
-0.229968488216400,
-0.230234414339066,
-0.230500578880310,
-0.230766981840134,
-0.231033623218536,
-0.231300503015518,
-0.231567621231079,
-0.231834977865219,
-0.232102558016777,
-0.232370376586914,
-0.232638433575630,
-0.232906728982925,
-0.233175262808800,
-0.233444035053253,
-0.233713045716286,
-0.233982294797897,
-0.234251797199249,
-0.234521523118019,
-0.234791502356529,
-0.235061705112457,
-0.235332161188126,
-0.235602855682373,
-0.235873773694038,
-0.236144945025444,
-0.236416354775429,
-0.236688002943993,
-0.236959889531136,
-0.237232014536858,
-0.237504377961159,
-0.237776979804039,
-0.238049834966660,
-0.238322913646698,
-0.238596245646477,
-0.238869816064835,
-0.239143639802933,
-0.239417672157288,
-0.239691957831383,
-0.239966467022896,
-0.240241214632988,
-0.240516215562820,
-0.240791454911232,
-0.241066932678223,
-0.241342663764954,
-0.241618633270264,
-0.241894856095314,
-0.242171302437782,
-0.242447987198830,
-0.242724940180779,
-0.243002131581306,
-0.243279546499252,
-0.243557214736938,
-0.243835121393204,
-0.244113296270370,
-0.244391694664955,
-0.244670331478119,
-0.244949221611023,
-0.245228365063667,
-0.245507746934891,
-0.245787367224693,
-0.246067240834236,
-0.246347367763519,
-0.246627718210220,
-0.246908321976662,
-0.247189179062843,
-0.247470274567604,
-0.247751608490944,
-0.248033210635185,
-0.248315036296844,
-0.248597130179405,
-0.248879462480545,
-0.249162048101425,
-0.249444872140884,
-0.249727949500084,
-0.250011265277863,
-0.250294834375381,
-0.250578641891480,
-0.250862717628479,
-0.251147001981735,
-0.251431554555893,
-0.251716345548630,
-0.252001345157623,
-0.252286642789841,
-0.252572149038315,
-0.252857923507690,
-0.253143936395645,
-0.253430217504501,
-0.253716737031937,
-0.254003524780273,
-0.254290521144867,
-0.254577785730362,
-0.254865318536758,
-0.255153089761734,
-0.255441099405289,
-0.255729377269745,
-0.256017893552780,
-0.256306648254395,
-0.256595671176910,
-0.256884932518005,
-0.257174462080002,
-0.257464230060577,
-0.257754266262054,
-0.258044540882111,
-0.258335083723068,
-0.258625864982605,
-0.258916884660721,
-0.259208172559738,
-0.259499698877335,
-0.259791493415833,
-0.260083526372910,
-0.260375827550888,
-0.260668367147446,
-0.260961174964905,
-0.261254221200943,
-0.261547505855560,
-0.261841058731079,
-0.262134879827499,
-0.262428969144821,
-0.262723267078400,
-0.263017863035202,
-0.263312667608261,
-0.263607710599899,
-0.263903021812439,
-0.264198571443558,
-0.264494419097900,
-0.264790475368500,
-0.265086799860001,
-0.265383392572403,
-0.265680223703384,
-0.265977323055267,
-0.266274690628052,
-0.266572296619415,
-0.266870141029358,
-0.267168253660202,
-0.267466634511948,
-0.267765253782272,
-0.268064171075821,
-0.268363326787949,
-0.268662720918655,
-0.268962353467941,
-0.269262284040451,
-0.269562453031540,
-0.269862860441208,
-0.270163565874100,
-0.270464509725571,
-0.270765721797943,
-0.271067172288895,
-0.271368920803070,
-0.271670877933502,
-0.271973133087158,
-0.272275626659393,
-0.272578388452530,
-0.272881418466568,
-0.273184686899185,
-0.273488253355026,
-0.273792028427124,
-0.274096101522446,
-0.274400413036346,
-0.274704992771149,
-0.275009840726852,
-0.275314897298813,
-0.275620222091675,
-0.275925815105438,
-0.276231646537781,
-0.276537775993347,
-0.276844143867493,
-0.277150750160217,
-0.277457654476166,
-0.277764797210693,
-0.278072208166122,
-0.278379917144775,
-0.278687834739685,
-0.278996050357819,
-0.279304504394531,
-0.279613226652145,
-0.279922217130661,
-0.280231475830078,
-0.280541002750397,
-0.280850768089294,
-0.281160801649094,
-0.281471103429794,
-0.281781673431397,
-0.282092511653900,
-0.282403618097305,
-0.282714962959290,
-0.283026605844498,
-0.283338487148285,
-0.283650636672974,
-0.283963084220886,
-0.284275770187378,
-0.284588694572449,
-0.284901916980743,
-0.285215407609940,
-0.285529136657715,
-0.285843133926392,
-0.286157429218292,
-0.286471962928772,
-0.286786764860153,
-0.287101835012436,
-0.287417143583298,
-0.287732690572739,
-0.288048565387726,
-0.288364678621292,
-0.288681060075760,
-0.288997709751129,
-0.289314627647400,
-0.289631813764572,
-0.289949268102646,
-0.290266960859299,
-0.290584981441498,
-0.290903240442276,
-0.291221737861633,
-0.291540533304215,
-0.291859567165375,
-0.292178899049759,
-0.292498499155045,
-0.292818367481232,
-0.293138474225998,
-0.293458908796310,
-0.293779581785202,
-0.294100522994995,
-0.294421732425690,
-0.294743239879608,
-0.295064985752106,
-0.295386999845505,
-0.295709311962128,
-0.296031892299652,
-0.296354711055756,
-0.296677827835083,
-0.297001212835312,
-0.297324866056442,
-0.297648787498474,
-0.297972977161407,
-0.298297464847565,
-0.298622190952301,
-0.298947155475616,
-0.299272418022156,
-0.299597948789597,
-0.299923747777939,
-0.300249814987183,
-0.300576150417328,
-0.300902783870697,
-0.301229655742645,
-0.301556795835495,
-0.301884263753891,
-0.302211970090866,
-0.302539974451065,
-0.302868217229843,
-0.303196758031845,
-0.303525567054749,
-0.303854644298553,
-0.304183989763260,
-0.304513633251190,
-0.304843544960022,
-0.305173724889755,
-0.305504202842712,
-0.305834919214249,
-0.306165933609009,
-0.306497216224670,
-0.306828767061234,
-0.307160615921021,
-0.307492733001709,
-0.307825148105621,
-0.308157801628113,
-0.308490753173828,
-0.308823943138123,
-0.309157460927963,
-0.309491217136383,
-0.309825301170349,
-0.310159623622894,
-0.310494244098663,
-0.310829102993012,
-0.311164230108261,
-0.311499625444412,
-0.311835318803787,
-0.312171280384064,
-0.312507510185242,
-0.312844038009644,
-0.313180834054947,
-0.313517928123474,
-0.313855260610580,
-0.314192920923233,
-0.314530819654465,
-0.314869046211243,
-0.315207511186600,
-0.315546274185181,
-0.315885335206986,
-0.316224634647369,
-0.316564261913300,
-0.316904157400131,
-0.317244321107864,
-0.317584782838821,
-0.317925512790680,
-0.318266510963440,
-0.318607807159424,
-0.318949371576309,
-0.319291234016418,
-0.319633364677429,
-0.319975793361664,
-0.320318490266800,
-0.320661485195160,
-0.321004748344421,
-0.321348309516907,
-0.321692138910294,
-0.322036296129227,
-0.322380661964417,
-0.322725355625153,
-0.323070317506790,
-0.323415547609329,
-0.323761045932770,
-0.324106812477112,
-0.324452906847000,
-0.324799269437790,
-0.325145900249481,
-0.325492829084396,
-0.325840055942535,
-0.326187551021576,
-0.326535344123840,
-0.326883405447006,
-0.327231764793396,
-0.327580422163010,
-0.327929347753525,
-0.328278571367264,
-0.328628063201904,
-0.328977853059769,
-0.329327940940857,
-0.329678297042847,
-0.330028951168060,
-0.330379873514175,
-0.330731093883514,
-0.331082612276077,
-0.331434398889542,
-0.331786483526230,
-0.332138866186142,
-0.332491517066956,
-0.332844465970993,
-0.333197712898254,
-0.333551228046417,
-0.333905071020126,
-0.334259152412415,
-0.334613561630249,
-0.334968209266663,
-0.335323154926300,
-0.335678398609161,
-0.336033910512924,
-0.336389720439911,
-0.336745828390121,
-0.337102204561234,
-0.337458878755569,
-0.337815850973129,
-0.338173121213913,
-0.338530689477921,
-0.338888525962830,
-0.339246660470963,
-0.339605093002319,
-0.339963793754578,
-0.340322822332382,
-0.340682119131088,
-0.341041713953018,
-0.341401606798172,
-0.341761767864227,
-0.342122256755829,
-0.342483043670654,
-0.342844098806381,
-0.343205422163010,
-0.343567073345184,
-0.343929022550583,
-0.344291239976883,
-0.344653785228729,
-0.345016598701477,
-0.345379680395126,
-0.345743089914322,
-0.346106797456741,
-0.346470773220062,
-0.346835047006607,
-0.347199618816376,
-0.347564458847046,
-0.347929626703262,
-0.348295032978058,
-0.348660767078400,
-0.349026769399643,
-0.349393099546433,
-0.349759697914124,
-0.350126624107361,
-0.350493848323822,
-0.350861340761185,
-0.351229161024094,
-0.351597279310226,
-0.351965695619583,
-0.352334380149841,
-0.352703392505646,
-0.353072702884674,
-0.353442311286926,
-0.353812187910080,
-0.354182362556458,
-0.354552835226059,
-0.354923605918884,
-0.355294674634933,
-0.355666041374207,
-0.356037706136704,
-0.356409668922424,
-0.356781929731369,
-0.357154488563538,
-0.357527375221252,
-0.357900530099869,
-0.358273983001709,
-0.358647704124451,
-0.359021753072739,
-0.359396070241928,
-0.359770685434341,
-0.360145658254623,
-0.360520899295807,
-0.360896468162537,
-0.361272335052490,
-0.361648470163345,
-0.362024933099747,
-0.362401694059372,
-0.362778753042221,
-0.363156110048294,
-0.363533765077591,
-0.363911718130112,
-0.364289969205856,
-0.364668548107147,
-0.365047395229340,
-0.365426540374756,
-0.365806043148041,
-0.366185814142227,
-0.366565912961960,
-0.366946309804916,
-0.367327004671097,
-0.367707997560501,
-0.368089288473129,
-0.368470877408981,
-0.368852794170380,
-0.369235008955002,
-0.369617551565170,
-0.370000362396240,
-0.370383501052856,
-0.370766878128052,
-0.371150583028793,
-0.371534615755081,
-0.371918916702271,
-0.372303545475006,
-0.372688472270966,
-0.373073697090149,
-0.373459219932556,
-0.373845100402832,
-0.374231249094009,
-0.374617725610733,
-0.375004470348358,
-0.375391542911530,
-0.375778943300247,
-0.376166641712189,
-0.376554638147354,
-0.376942932605743,
-0.377331554889679,
-0.377720504999161,
-0.378109753131866,
-0.378499269485474,
-0.378889113664627,
-0.379279285669327,
-0.379669755697250,
-0.380060553550720,
-0.380451619625092,
-0.380843043327332,
-0.381234735250473,
-0.381626754999161,
-0.382019102573395,
-0.382411718368530,
-0.382804632186890,
-0.383197844028473,
-0.383591383695602,
-0.383985251188278,
-0.384379386901855,
-0.384773880243301,
-0.385168671607971,
-0.385563760995865,
-0.385959178209305,
-0.386354893445969,
-0.386750936508179,
-0.387147307395935,
-0.387543946504593,
-0.387940913438797,
-0.388338238000870,
-0.388735830783844,
-0.389133721590042,
-0.389531970024109,
-0.389930516481400,
-0.390329360961914,
-0.390728533267975,
-0.391128033399582,
-0.391527831554413,
-0.391927957534790,
-0.392328381538391,
-0.392729133367538,
-0.393130183219910,
-0.393531560897827,
-0.393933266401291,
-0.394335210323334,
-0.394737511873245,
-0.395140111446381,
-0.395543038845062,
-0.395946264266968,
-0.396349817514420,
-0.396753668785095,
-0.397157847881317,
-0.397562354803085,
-0.397967189550400,
-0.398372322320938,
-0.398777782917023,
-0.399183571338654,
-0.399589657783508,
-0.399996101856232,
-0.400402814149857,
-0.400809854269028,
-0.401217222213745,
-0.401624888181686,
-0.402032881975174,
-0.402441203594208,
-0.402849853038788,
-0.403258800506592,
-0.403668075799942,
-0.404077678918839,
-0.404487609863281,
-0.404897868633270,
-0.405308425426483,
-0.405719310045242,
-0.406130522489548,
-0.406542032957077,
-0.406953841447830,
-0.407365977764130,
-0.407778412103653,
-0.408191174268723,
-0.408604264259338,
-0.409017682075501,
-0.409431457519531,
-0.409845501184464,
-0.410259902477264,
-0.410674601793289,
-0.411089628934860,
-0.411504983901978,
-0.411920636892319,
-0.412336647510529,
-0.412752985954285,
-0.413169622421265,
-0.413586586713791,
-0.414003878831863,
-0.414421498775482,
-0.414839446544647,
-0.415257722139359,
-0.415676325559616,
-0.416095256805420,
-0.416514486074448,
-0.416934072971344,
-0.417353987693787,
-0.417774200439453,
-0.418194741010666,
-0.418615549802780,
-0.419036716222763,
-0.419458240270615,
-0.419880032539368,
-0.420302182435989,
-0.420724660158157,
-0.421147435903549,
-0.421570569276810,
-0.421994030475616,
-0.422417789697647,
-0.422841906547546,
-0.423266351222992,
-0.423691093921661,
-0.424116164445877,
-0.424541592597961,
-0.424967348575592,
-0.425393432378769,
-0.425819814205170,
-0.426246553659439,
-0.426673650741577,
-0.427101016044617,
-0.427528738975525,
-0.427956789731979,
-0.428385198116303,
-0.428813904523850,
-0.429242938756943,
-0.429672330617905,
-0.430102020502090,
-0.430532008409500,
-0.430962324142456,
-0.431392967700958,
-0.431823968887329,
-0.432255297899246,
-0.432686924934387,
-0.433118909597397,
-0.433551222085953,
-0.433983862400055,
-0.434416860342026,
-0.434850156307220,
-0.435283780097961,
-0.435717761516571,
-0.436152070760727,
-0.436586737632751,
-0.437021702528000,
-0.437456995248795,
-0.437892645597458,
-0.438328623771668,
-0.438764929771423,
-0.439201563596725,
-0.439638555049896,
-0.440075874328613,
-0.440513521432877,
-0.440951496362686,
-0.441389799118042,
-0.441828459501267,
-0.442267388105392,
-0.442706674337387,
-0.443146288394928,
-0.443586260080338,
-0.444026559591293,
-0.444467157125473,
-0.444908112287521,
-0.445349395275116,
-0.445791006088257,
-0.446232974529266,
-0.446675270795822,
-0.447117924690247,
-0.447560906410217,
-0.448004215955734,
-0.448447883129120,
-0.448891878128052,
-0.449336230754852,
-0.449780911207199,
-0.450225919485092,
-0.450671285390854,
-0.451116979122162,
-0.451563030481339,
-0.452009379863739,
-0.452456057071686,
-0.452903091907501,
-0.453350454568863,
-0.453798145055771,
-0.454246133565903,
-0.454694479703903,
-0.455143153667450,
-0.455592185258865,
-0.456041544675827,
-0.456491231918335,
-0.456941276788712,
-0.457391649484634,
-0.457842350006104,
-0.458293437957764,
-0.458744883537293,
-0.459196656942368,
-0.459648758172989,
-0.460101217031479,
-0.460554033517838,
-0.461007148027420,
-0.461460620164871,
-0.461914449930191,
-0.462368607521057,
-0.462823092937470,
-0.463277935981751,
-0.463733106851578,
-0.464188635349274,
-0.464644491672516,
-0.465100675821304,
-0.465557217597961,
-0.466014087200165,
-0.466471284627914,
-0.466928839683533,
-0.467386722564697,
-0.467844963073730,
-0.468303531408310,
-0.468762427568436,
-0.469221681356430,
-0.469681292772293,
-0.470141261816025,
-0.470601558685303,
-0.471062213182449,
-0.471523195505142,
-0.471984535455704,
-0.472446203231812,
-0.472908228635788,
-0.473370611667633,
-0.473833352327347,
-0.474296420812607,
-0.474759817123413,
-0.475223571062088,
-0.475687682628632,
-0.476152122020721,
-0.476616919040680,
-0.477082073688507,
-0.477547556161881,
-0.478013366460800,
-0.478479474782944,
-0.478946000337601,
-0.479412823915482,
-0.479880034923553,
-0.480347543954849,
-0.480815410614014,
-0.481283664703369,
-0.481752246618271,
-0.482221186161041,
-0.482690453529358,
-0.483160108327866,
-0.483630090951920,
-0.484100431203842,
-0.484571099281311,
-0.485042095184326,
-0.485513508319855,
-0.485985219478607,
-0.486457288265228,
-0.486929714679718,
-0.487402498722076,
-0.487875640392303,
-0.488349109888077,
-0.488822966814041,
-0.489297151565552,
-0.489771664142609,
-0.490246474742889,
-0.490721672773361,
-0.491197228431702,
-0.491673111915588,
-0.492149382829666,
-0.492625981569290,
-0.493102937936783,
-0.493580251932144,
-0.494057893753052,
-0.494535923004150,
-0.495014280080795,
-0.495492994785309,
-0.495972067117691,
-0.496451497077942,
-0.496931284666061,
-0.497411429882050,
-0.497891902923584,
-0.498372733592987,
-0.498853951692581,
-0.499335467815399,
-0.499817401170731,
-0.500299632549286,
-0.500782251358032,
-0.501265227794647,
-0.501748502254486,
-0.502232134342194,
-0.502716124057770,
-0.503200471401215,
-0.503685176372528,
-0.504170238971710,
-0.504655659198761,
-0.505141437053680,
-0.505627572536469,
-0.506114065647125,
-0.506600916385651,
-0.507088124752045,
-0.507575631141663,
-0.508063554763794,
-0.508551836013794,
-0.509040474891663,
-0.509529471397400,
-0.510018765926361,
-0.510508477687836,
-0.510998547077179,
-0.511488974094391,
-0.511979758739471,
-0.512470841407776,
-0.512962341308594,
-0.513454198837280,
-0.513946354389191,
-0.514438927173615,
-0.514931797981262,
-0.515425026416779,
-0.515918612480164,
-0.516412556171417,
-0.516906857490540,
-0.517401576042175,
-0.517896592617035,
-0.518391966819763,
-0.518887698650360,
-0.519383847713471,
-0.519880294799805,
-0.520377159118652,
-0.520874381065369,
-0.521371901035309,
-0.521869838237763,
-0.522368133068085,
-0.522866785526276,
-0.523365795612335,
-0.523865103721619,
-0.524364888668060,
-0.524864971637726,
-0.525365412235260,
-0.525866210460663,
-0.526367366313934,
-0.526868820190430,
-0.527370691299439,
-0.527872920036316,
-0.528375506401062,
-0.528878450393677,
-0.529381752014160,
-0.529885411262512,
-0.530389487743378,
-0.530893862247467,
-0.531398653984070,
-0.531903743743897,
-0.532409250736237,
-0.532915115356445,
-0.533421337604523,
-0.533927977085114,
-0.534434914588928,
-0.534942209720612,
-0.535449922084808,
-0.535957992076874,
-0.536466419696808,
-0.536975145339966,
-0.537484288215637,
-0.537993729114533,
-0.538503587245941,
-0.539013743400574,
-0.539524316787720,
-0.540035247802734,
-0.540546596050263,
-0.541058242321014,
-0.541570246219635,
-0.542082667350769,
-0.542595386505127,
-0.543108522891998,
-0.543622016906738,
-0.544135868549347,
-0.544650137424469,
-0.545164763927460,
-0.545679688453674,
-0.546195030212402,
-0.546710729598999,
-0.547226786613464,
-0.547743260860443,
-0.548260092735291,
-0.548777282238007,
-0.549294829368591,
-0.549812674522400,
-0.550330936908722,
-0.550849556922913,
-0.551368534564972,
-0.551887869834900,
-0.552407622337341,
-0.552927732467651,
-0.553448140621185,
-0.553969025611877,
-0.554490208625794,
-0.555011749267578,
-0.555533707141876,
-0.556056022644043,
-0.556578695774078,
-0.557101786136627,
-0.557625174522400,
-0.558149039745331,
-0.558673202991486,
-0.559197723865509,
-0.559722661972046,
-0.560247957706451,
-0.560773611068726,
-0.561299622058868,
-0.561825990676880,
-0.562352716922760,
-0.562879860401154,
-0.563407301902771,
-0.563935160636902,
-0.564463376998901,
-0.564992010593414,
-0.565520942211151,
-0.566050350666046,
-0.566580057144165,
-0.567110121250153,
-0.567640602588654,
-0.568171441555023,
-0.568702638149262,
-0.569234251976013,
-0.569766223430634,
-0.570298552513123,
-0.570831239223480,
-0.571364343166351,
-0.571897864341736,
-0.572431683540344,
-0.572965919971466,
-0.573500454425812,
-0.574035346508026,
-0.574570655822754,
-0.575106322765350,
-0.575642347335815,
-0.576178789138794,
-0.576715588569641,
-0.577252745628357,
-0.577790319919586,
-0.578328251838684,
-0.578866541385651,
-0.579405248165131,
-0.579944312572479,
-0.580483734607697,
-0.581023573875427,
-0.581563770771027,
-0.582104384899139,
-0.582645297050476,
-0.583186626434326,
-0.583728313446045,
-0.584270417690277,
-0.584812879562378,
-0.585355699062347,
-0.585898876190186,
-0.586442410945892,
-0.586986362934113,
-0.587530672550201,
-0.588075399398804,
-0.588620483875275,
-0.589165925979614,
-0.589711785316467,
-0.590257942676544,
-0.590804517269135,
-0.591351509094238,
-0.591898858547211,
-0.592446565628052,
-0.592994630336762,
-0.593543171882629,
-0.594092011451721,
-0.594641268253326,
-0.595190882682800,
-0.595740914344788,
-0.596291303634644,
-0.596842110157013,
-0.597393155097961,
-0.597944676876068,
-0.598496556282044,
-0.599048793315888,
-0.599601387977600,
-0.600154399871826,
-0.600707828998566,
-0.601261615753174,
-0.601815760135651,
-0.602370262145996,
-0.602925240993500,
-0.603480517864227,
-0.604036211967468,
-0.604592263698578,
-0.605148732662201,
-0.605705559253693,
-0.606262803077698,
-0.606820464134216,
-0.607378542423248,
-0.607936978340149,
-0.608495771884918,
-0.609054982662201,
-0.609614491462708,
-0.610174417495728,
-0.610734701156616,
-0.611295402050018,
-0.611856460571289,
-0.612417876720429,
-0.612979710102081,
-0.613541901111603,
-0.614104509353638,
-0.614667475223541,
-0.615230798721314,
-0.615794539451599,
-0.616358637809753,
-0.616923153400421,
-0.617488026618958,
-0.618053376674652,
-0.618619143962860,
-0.619185209274292,
-0.619751691818237,
-0.620318591594696,
-0.620885848999023,
-0.621453404426575,
-0.622021377086639,
-0.622589707374573,
-0.623158454895020,
-0.623727560043335,
-0.624297082424164,
-0.624866962432861,
-0.625437200069428,
-0.626007914543152,
-0.626578986644745,
-0.627150475978851,
-0.627722382545471,
-0.628294587135315,
-0.628867208957672,
-0.629440248012543,
-0.630013644695282,
-0.630587458610535,
-0.631161630153656,
-0.631736218929291,
-0.632311224937439,
-0.632886648178101,
-0.633462309837341,
-0.634038448333740,
-0.634614884853363,
-0.635191738605499,
-0.635769009590149,
-0.636346638202667,
-0.636924743652344,
-0.637503206729889,
-0.638082027435303,
-0.638661265373230,
-0.639240920543671,
-0.639820933341980,
-0.640401303768158,
-0.640982091426849,
-0.641563296318054,
-0.642144918441773,
-0.642726898193359,
-0.643309295177460,
-0.643892049789429,
-0.644475162029266,
-0.645058631896973,
-0.645642578601837,
-0.646226882934570,
-0.646811604499817,
-0.647396683692932,
-0.647982120513916,
-0.648567974567413,
-0.649154186248779,
-0.649740874767304,
-0.650327920913696,
-0.650915384292603,
-0.651503264904022,
-0.652091443538666,
-0.652680039405823,
-0.653269112110138,
-0.653858602046967,
-0.654448390007019,
-0.655038654804230,
-0.655629217624664,
-0.656220197677612,
-0.656811594963074,
-0.657403349876404,
-0.657995522022247,
-0.658588051795960,
-0.659180939197540,
-0.659774243831635,
-0.660368025302887,
-0.660962164402008,
-0.661556661128998,
-0.662151575088501,
-0.662746846675873,
-0.663342654705048,
-0.663938760757446,
-0.664535284042358,
-0.665132224559784,
-0.665729463100433,
-0.666327238082886,
-0.666925370693207,
-0.667523860931397,
-0.668122768402100,
-0.668722033500671,
-0.669321715831757,
-0.669921755790710,
-0.670522212982178,
-0.671123027801514,
-0.671724259853363,
-0.672325909137726,
-0.672927975654602,
-0.673530459403992,
-0.674133300781250,
-0.674736559391022,
-0.675340235233307,
-0.675944328308106,
-0.676548779010773,
-0.677153587341309,
-0.677758872509003,
-0.678364515304565,
-0.678970575332642,
-0.679577052593231,
-0.680183947086334,
-0.680791139602661,
-0.681398749351502,
-0.682006776332855,
-0.682615220546722,
-0.683224022388458,
-0.683833241462708,
-0.684442877769470,
-0.685052871704102,
-0.685663282871246,
-0.686274111270905,
-0.686885356903076,
-0.687496960163117,
-0.688109040260315,
-0.688721477985382,
-0.689334332942963,
-0.689947605133057,
-0.690561294555664,
-0.691175341606140,
-0.691789805889130,
-0.692404687404633,
-0.693019926548004,
-0.693635523319244,
-0.694251537322998,
-0.694867968559265,
-0.695484817028046,
-0.696102082729340,
-0.696719646453857,
-0.697337746620178,
-0.697956204414368,
-0.698575019836426,
-0.699194371700287,
-0.699814021587372,
-0.700434088706970,
-0.701054573059082,
-0.701675474643707,
-0.702296793460846,
-0.702918469905853,
-0.703540623188019,
-0.704163193702698,
-0.704786002635956,
-0.705409228801727,
-0.706032931804657,
-0.706657052040100,
-0.707281529903412,
-0.707906424999237,
-0.708531737327576,
-0.709157466888428,
-0.709783613681793,
-0.710410177707672,
-0.711037099361420,
-0.711664497852325,
-0.712292253971100,
-0.712920427322388,
-0.713548958301544,
-0.714177966117859,
-0.714807391166687,
-0.715437173843384,
-0.716067433357239,
-0.716697990894318,
-0.717328906059265,
-0.717960298061371,
-0.718592107295990,
-0.719224274158478,
-0.719856917858124,
-0.720489919185638,
-0.721123337745667,
-0.721757233142853,
-0.722391486167908,
-0.723026096820831,
-0.723661243915558,
-0.724296689033508,
-0.724932551383972,
-0.725568890571594,
-0.726205646991730,
-0.726842761039734,
-0.727480292320252,
-0.728118300437927,
-0.728756546974182,
-0.729395270347595,
-0.730034410953522,
-0.730673968791962,
-0.731313943862915,
-0.731954276561737,
-0.732595086097717,
-0.733236312866211,
-0.733877897262573,
-0.734519898891449,
-0.735162377357483,
-0.735805153846741,
-0.736448466777802,
-0.737092137336731,
-0.737736225128174,
-0.738380730152130,
-0.739025652408600,
-0.739671051502228,
-0.740316689014435,
-0.740962743759155,
-0.741609275341034,
-0.742256164550781,
-0.742903590202332,
-0.743551313877106,
-0.744199454784393,
-0.744848072528839,
-0.745497047901154,
-0.746146500110626,
-0.746796369552612,
-0.747446596622467,
-0.748097300529480,
-0.748748362064362,
-0.749399900436401,
-0.750051796436310,
-0.750704109668732,
-0.751356899738312,
-0.752010047435761,
-0.752663612365723,
-0.753317534923554,
-0.753971874713898,
-0.754626631736755,
-0.755281805992127,
-0.755937457084656,
-0.756593465805054,
-0.757249891757965,
-0.757906734943390,
-0.758563995361328,
-0.759221732616425,
-0.759879827499390,
-0.760538399219513,
-0.761197328567505,
-0.761856675148010,
-0.762516498565674,
-0.763176679611206,
-0.763837337493897,
-0.764498293399811,
-0.765159726142883,
-0.765821516513825,
-0.766483724117279,
-0.767146348953247,
-0.767809391021729,
-0.768472909927368,
-0.769136846065521,
-0.769801199436188,
-0.770465910434723,
-0.771131098270416,
-0.771796643733978,
-0.772462666034699,
-0.773129105567932,
-0.773795962333679,
-0.774463236331940,
-0.775130927562714,
-0.775799095630646,
-0.776467502117157,
-0.777136445045471,
-0.777805745601654,
-0.778475463390350,
-0.779145598411560,
-0.779816150665283,
-0.780487179756165,
-0.781158566474915,
-0.781830430030823,
-0.782502651214600,
-0.783175408840179,
-0.783848464488983,
-0.784522056579590,
-0.785196006298065,
-0.785870373249054,
-0.786545217037201,
-0.787220478057861,
-0.787896096706390,
-0.788572132587433,
-0.789248526096344,
-0.789925456047058,
-0.790602684020996,
-0.791280388832092,
-0.791958510875702,
-0.792636990547180,
-0.793316006660461,
-0.793995320796967,
-0.794675171375275,
-0.795355379581451,
-0.796036064624786,
-0.796717107295990,
-0.797398626804352,
-0.798080563545227,
-0.798762917518616,
-0.799445688724518,
-0.800128877162933,
-0.800812423229218,
-0.801496386528015,
-0.802180826663971,
-0.802865624427795,
-0.803550899028778,
-0.804236590862274,
-0.804922699928284,
-0.805609226226807,
-0.806296288967133,
-0.806983649730682,
-0.807671546936035,
-0.808359801769257,
-0.809048533439636,
-0.809737622737885,
-0.810427188873291,
-0.811117172241211,
-0.811807572841644,
-0.812498331069946,
-0.813189506530762,
-0.813881099224091,
-0.814573168754578,
-0.815265595912933,
-0.815958499908447,
-0.816651821136475,
-0.817345559597015,
-0.818039715290070,
-0.818734288215637,
-0.819429397583008,
-0.820124864578247,
-0.820820748806000,
-0.821517050266266,
-0.822213828563690,
-0.822911024093628,
-0.823608636856079,
-0.824306607246399,
-0.825004994869232,
-0.825703799724579,
-0.826403021812439,
-0.827102720737457,
-0.827802836894989,
-0.828503429889679,
-0.829204380512238,
-0.829905807971954,
-0.830607593059540,
-0.831309854984283,
-0.832012534141541,
-0.832715690135956,
-0.833419263362885,
-0.834123253822327,
-0.834827661514282,
-0.835532546043396,
-0.836237728595734,
-0.836943328380585,
-0.837649405002594,
-0.838355958461762,
-0.839062869548798,
-0.839770257472992,
-0.840478003025055,
-0.841186285018921,
-0.841894924640656,
-0.842603981494904,
-0.843313574790955,
-0.844023466110230,
-0.844733893871307,
-0.845444679260254,
-0.846156001091003,
-0.846867620944977,
-0.847579777240753,
-0.848292231559753,
-0.849005162715912,
-0.849718511104584,
-0.850432217121124,
-0.851146459579468,
-0.851861119270325,
-0.852576196193695,
-0.853291690349579,
-0.854007601737976,
-0.854723989963532,
-0.855440855026245,
-0.856158077716827,
-0.856875777244568,
-0.857593894004822,
-0.858312427997589,
-0.859031438827515,
-0.859750747680664,
-0.860470533370972,
-0.861190736293793,
-0.861911356449127,
-0.862632453441620,
-0.863353967666626,
-0.864075958728790,
-0.864798307418823,
-0.865521132946014,
-0.866244375705719,
-0.866968035697937,
-0.867692172527313,
-0.868416726589203,
-0.869141697883606,
-0.869867205619812,
-0.870593011379242,
-0.871319353580475,
-0.872046053409576,
-0.872773110866547,
-0.873500645160675,
-0.874228596687317,
-0.874957025051117,
-0.875685870647430,
-0.876415133476257,
-0.877144873142242,
-0.877875030040741,
-0.878605604171753,
-0.879336655139923,
-0.880068063735962,
-0.880800008773804,
-0.881532371044159,
-0.882265090942383,
-0.882998347282410,
-0.883731901645660,
-0.884465932846069,
-0.885200381278992,
-0.885935306549072,
-0.886670589447022,
-0.887406349182129,
-0.888142585754395,
-0.888879239559174,
-0.889616310596466,
-0.890353798866272,
-0.891091763973236,
-0.891830205917358,
-0.892569005489349,
-0.893308281898499,
-0.894048035144806,
-0.894788146018982,
-0.895528674125671,
-0.896269619464874,
-0.897010982036591,
-0.897752821445465,
-0.898495137691498,
-0.899237811565399,
-0.899980962276459,
-0.900724589824677,
-0.901468575000763,
-0.902213037014008,
-0.902957975864410,
-0.903703331947327,
-0.904449105262756,
-0.905195355415344,
-0.905942022800446,
-0.906689167022705,
-0.907436668872833,
-0.908184528350830,
-0.908932864665985,
-0.909681677818298,
-0.910430908203125,
-0.911180615425110,
-0.911930739879608,
-0.912681281566620,
-0.913432240486145,
-0.914183735847473,
-0.914935588836670,
-0.915687918663025,
-0.916440725326538,
-0.917193889617920,
-0.917947530746460,
-0.918701648712158,
-0.919456064701080,
-0.920210957527161,
-0.920966267585754,
-0.921722054481506,
-0.922478258609772,
-0.923234879970551,
-0.923991978168488,
-0.924749493598938,
-0.925507485866547,
-0.926265895366669,
-0.927024722099304,
-0.927784025669098,
-0.928543746471405,
-0.929303944110870,
-0.930064558982849,
-0.930825710296631,
-0.931587100028992,
-0.932348966598511,
-0.933111310005188,
-0.933874070644379,
-0.934637248516083,
-0.935400903224945,
-0.936164975166321,
-0.936929523944855,
-0.937694489955902,
-0.938459992408752,
-0.939225792884827,
-0.939992129802704,
-0.940758943557739,
-0.941526114940643,
-0.942293763160706,
-0.943061769008637,
-0.943830192089081,
-0.944599032402039,
-0.945368409156799,
-0.946138203144074,
-0.946908414363861,
-0.947679102420807,
-0.948450207710266,
-0.949221730232239,
-0.949993729591370,
-0.950766205787659,
-0.951539158821106,
-0.952312469482422,
-0.953086256980896,
-0.953860521316528,
-0.954635143280029,
-0.955410182476044,
-0.956185638904572,
-0.956961631774902,
-0.957737982273102,
-0.958514809608460,
-0.959292054176331,
-0.960069715976715,
-0.960847914218903,
-0.961626470088959,
-0.962405562400818,
-0.963185071945190,
-0.963964998722076,
-0.964745402336121,
-0.965526163578033,
-0.966307461261749,
-0.967089056968689,
-0.967871189117432,
-0.968653678894043,
-0.969436645507813,
-0.970220088958740,
-0.971003949642181,
-0.971788287162781,
-0.972573041915894,
-0.973358273506165,
-0.974143862724304,
-0.974929988384247,
-0.975716531276703,
-0.976503551006317,
-0.977290928363800,
-0.978078842163086,
-0.978867113590241,
-0.979655802249908,
-0.980444908142090,
-0.981234490871429,
-0.982024550437927,
-0.982815086841583,
-0.983605980873108,
-0.984397351741791,
-0.985189199447632,
-0.985981523990631,
-0.986774206161499,
-0.987567424774170,
-0.988361060619354,
-0.989155113697052,
-0.989949584007263,
-0.990744590759277,
-0.991539895534515,
-0.992335617542267,
-0.993131875991821,
-0.993928492069244,
-0.994725644588471,
-0.995523214340210,
-0.996321201324463,
-0.997119665145874,
-0.997918605804443,
-0.998717904090881,
-0.999517738819122,
-1.00031805038452,
-1.00111877918243,
-1.00191986560822,
-1.00272130966187,
-1.00352334976196,
-1.00432574748993,
-1.00512862205505,
-1.00593185424805,
-1.00673568248749,
-1.00753986835480,
-1.00834453105927,
-1.00914967060089,
-1.00995528697968,
-1.01076126098633,
-1.01156783103943,
-1.01237463951111,
-1.01318204402924,
-1.01398980617523,
-1.01479804515839,
-1.01560664176941,
-1.01641571521759,
-1.01722526550293,
-1.01803529262543,
-1.01884567737579,
-1.01965653896332,
-1.02046787738800,
-1.02127957344055,
-1.02209186553955,
-1.02290451526642,
-1.02371764183044,
-1.02453124523163,
-1.02534532546997,
-1.02615976333618,
-1.02697467803955,
-1.02778995037079,
-1.02860569953918,
-1.02942192554474,
-1.03023850917816,
-1.03105556964874,
-1.03187322616577,
-1.03269124031067,
-1.03350961208344,
-1.03432857990265,
-1.03514790534973,
-1.03596770763397,
-1.03678798675537,
-1.03760874271393,
-1.03842985630035,
-1.03925144672394,
-1.04007339477539,
-1.04089581966400,
-1.04171872138977,
-1.04254209995270,
-1.04336583614349,
-1.04419016838074,
-1.04501485824585,
-1.04583990573883,
-1.04666554927826,
-1.04749166965485,
-1.04831814765930,
-1.04914510250092,
-1.04997253417969,
-1.05080032348633,
-1.05162858963013,
-1.05245721340179,
-1.05328631401062,
-1.05411589145660,
-1.05494594573975,
-1.05577647686005,
-1.05660736560822,
-1.05743873119354,
-1.05827057361603,
-1.05910289287567,
-1.05993568897247,
-1.06076896190643,
-1.06160259246826,
-1.06243658065796,
-1.06327104568481,
-1.06410598754883,
-1.06494140625000,
-1.06577718257904,
-1.06661355495453,
-1.06745028495789,
-1.06828749179840,
-1.06912517547607,
-1.06996321678162,
-1.07080173492432,
-1.07164084911346,
-1.07248032093048,
-1.07332026958466,
-1.07416069507599,
-1.07500135898590,
-1.07584261894226,
-1.07668423652649,
-1.07752645015717,
-1.07836902141571,
-1.07921195030212,
-1.08005547523499,
-1.08089935779572,
-1.08174383640289,
-1.08258867263794,
-1.08343398571014,
-1.08427977561951,
-1.08512592315674,
-1.08597266674042,
-1.08681976795197,
-1.08766722679138,
-1.08851516246796,
-1.08936345577240,
-1.09021234512329,
-1.09106171131134,
-1.09191143512726,
-1.09276163578033,
-1.09361231327057,
-1.09446346759796,
-1.09531509876251,
-1.09616720676422,
-1.09701979160309,
-1.09787273406982,
-1.09872603416443,
-1.09957981109619,
-1.10043406486511,
-1.10128867626190,
-1.10214388370514,
-1.10299944877625,
-1.10385560989380,
-1.10471212863922,
-1.10556912422180,
-1.10642647743225,
-1.10728442668915,
-1.10814285278320,
-1.10900163650513,
-1.10986089706421,
-1.11072051525116,
-1.11158061027527,
-1.11244118213654,
-1.11330211162567,
-1.11416363716125,
-1.11502552032471,
-1.11588788032532,
-1.11675071716309,
-1.11761403083801,
-1.11847782135010,
-1.11934208869934,
-1.12020671367645,
-1.12107181549072,
-1.12193739414215,
-1.12280344963074,
-1.12366986274719,
-1.12453675270081,
-1.12540400028229,
-1.12627184391022,
-1.12714004516602,
-1.12800872325897,
-1.12887787818909,
-1.12974762916565,
-1.13061773777008,
-1.13148820400238,
-1.13235926628113,
-1.13323068618774,
-1.13410246372223,
-1.13497483730316,
-1.13584756851196,
-1.13672077655792,
-1.13759446144104,
-1.13846850395203,
-1.13934314250946,
-1.14021813869476,
-1.14109361171722,
-1.14196968078613,
-1.14284610748291,
-1.14372289180756,
-1.14460027217865,
-1.14547801017761,
-1.14635622501373,
-1.14723479747772,
-1.14811396598816,
-1.14899349212646,
-1.14987349510193,
-1.15075397491455,
-1.15163493156433,
-1.15251624584198,
-1.15339815616608,
-1.15428042411804,
-1.15516316890717,
-1.15604650974274,
-1.15693020820618,
-1.15781426429749,
-1.15869867801666,
-1.15958368778229,
-1.16046905517578,
-1.16135501861572,
-1.16224133968353,
-1.16312825679779,
-1.16401553153992,
-1.16490328311920,
-1.16579139232636,
-1.16668009757996,
-1.16756916046143,
-1.16845881938934,
-1.16934883594513,
-1.17023932933807,
-1.17113018035889,
-1.17202150821686,
-1.17291331291199,
-1.17380559444428,
-1.17469823360443,
-1.17559146881104,
-1.17648506164551,
-1.17737925052643,
-1.17827379703522,
-1.17916893959045,
-1.18006443977356,
-1.18096041679382,
-1.18185663223267,
-1.18275344371796,
-1.18365061283112,
-1.18454837799072,
-1.18544650077820,
-1.18634521961212,
-1.18724429607391,
-1.18814396858215,
-1.18904387950897,
-1.18994438648224,
-1.19084537029266,
-1.19174671173096,
-1.19264864921570,
-1.19355082511902,
-1.19445359706879,
-1.19535672664642,
-1.19626033306122,
-1.19716453552246,
-1.19806909561157,
-1.19897413253784,
-1.19987952709198,
-1.20078551769257,
-1.20169186592102,
-1.20259881019592,
-1.20350611209869,
-1.20441389083862,
-1.20532226562500,
-1.20623087882996,
-1.20713996887207,
-1.20804953575134,
-1.20895969867706,
-1.20987021923065,
-1.21078121662140,
-1.21169269084930,
-1.21260464191437,
-1.21351695060730,
-1.21442961692810,
-1.21534287929535,
-1.21625661849976,
-1.21717071533203,
-1.21808528900146,
-1.21900022029877,
-1.21991574764252,
-1.22083163261414,
-1.22174811363220,
-1.22266495227814,
-1.22358226776123,
-1.22450017929077,
-1.22541844844818,
-1.22633719444275,
-1.22725641727448,
-1.22817611694336,
-1.22909641265869,
-1.23001694679260,
-1.23093795776367,
-1.23185944557190,
-1.23278129100800,
-1.23370373249054,
-1.23462665081024,
-1.23555004596710,
-1.23647379875183,
-1.23739790916443,
-1.23832261562347,
-1.23924767971039,
-1.24017333984375,
-1.24109935760498,
-1.24202573299408,
-1.24295270442963,
-1.24388003349304,
-1.24480783939362,
-1.24573612213135,
-1.24666488170624,
-1.24759411811829,
-1.24852395057678,
-1.24945414066315,
-1.25038480758667,
-1.25131595134735,
-1.25224745273590,
-1.25317943096161,
-1.25411188602448,
-1.25504481792450,
-1.25597822666168,
-1.25691199302673,
-1.25784635543823,
-1.25878119468689,
-1.25971639156342,
-1.26065218448639,
-1.26158845424652,
-1.26252508163452,
-1.26346230506897,
-1.26439988613129,
-1.26533770561218,
-1.26627600193024,
-1.26721489429474,
-1.26815414428711,
-1.26909387111664,
-1.27003407478333,
-1.27097475528717,
-1.27191591262817,
-1.27285754680634,
-1.27379953861237,
-1.27474212646484,
-1.27568519115448,
-1.27662873268127,
-1.27757263183594,
-1.27851688861847,
-1.27946174144745,
-1.28040707111359,
-1.28135275840759,
-1.28229904174805,
-1.28324568271637,
-1.28419291973114,
-1.28514051437378,
-1.28608870506287,
-1.28703725337982,
-1.28798627853394,
-1.28893589973450,
-1.28988575935364,
-1.29083609580994,
-1.29178690910339,
-1.29273831844330,
-1.29369008541107,
-1.29464232921600,
-1.29559504985809,
-1.29654824733734,
-1.29750192165375,
-1.29845607280731,
-1.29941070079803,
-1.30036580562592,
-1.30132126808167,
-1.30227708816528,
-1.30323338508606,
-1.30419003963470,
-1.30514729022980,
-1.30610489845276,
-1.30706310272217,
-1.30802166461945,
-1.30898082256317,
-1.30994033813477,
-1.31090033054352,
-1.31186091899872,
-1.31282174587250,
-1.31378304958344,
-1.31474483013153,
-1.31570708751678,
-1.31666994094849,
-1.31763315200806,
-1.31859683990479,
-1.31956100463867,
-1.32052564620972,
-1.32149076461792,
-1.32245635986328,
-1.32342243194580,
-1.32438886165619,
-1.32535576820374,
-1.32632315158844,
-1.32729101181030,
-1.32825922966003,
-1.32922804355621,
-1.33019733428955,
-1.33116698265076,
-1.33213722705841,
-1.33310794830322,
-1.33407902717590,
-1.33505070209503,
-1.33602273464203,
-1.33699512481689,
-1.33796811103821,
-1.33894145488739,
-1.33991527557373,
-1.34088969230652,
-1.34186446666718,
-1.34283971786499,
-1.34381544589996,
-1.34479176998138,
-1.34576845169067,
-1.34674561023712,
-1.34772324562073,
-1.34870123863220,
-1.34967970848084,
-1.35065865516663,
-1.35163807868958,
-1.35261797904968,
-1.35359835624695,
-1.35457921028137,
-1.35556042194366,
-1.35654222965240,
-1.35752451419830,
-1.35850727558136,
-1.35949027538300,
-1.36047387123108,
-1.36145770549774,
-1.36244201660156,
-1.36342692375183,
-1.36441218852997,
-1.36539793014526,
-1.36638426780701,
-1.36737096309662,
-1.36835813522339,
-1.36934578418732,
-1.37033402919769,
-1.37132263183594,
-1.37231171131134,
-1.37330114841461,
-1.37429106235504,
-1.37528145313263,
-1.37627232074738,
-1.37726366519928,
-1.37825548648834,
-1.37924766540527,
-1.38024044036865,
-1.38123369216919,
-1.38222742080688,
-1.38322162628174,
-1.38421618938446,
-1.38521122932434,
-1.38620674610138,
-1.38720262050629,
-1.38819909095764,
-1.38919591903687,
-1.39019334316254,
-1.39119112491608,
-1.39218950271606,
-1.39318823814392,
-1.39418756961823,
-1.39518725872040,
-1.39618754386902,
-1.39718806743622,
-1.39818906784058,
-1.39919054508209,
-1.40019261837006,
-1.40119504928589,
-1.40219795703888,
-1.40320134162903,
-1.40420520305634,
-1.40520954132080,
-1.40621447563171,
-1.40721976757050,
-1.40822541713715,
-1.40923142433167,
-1.41023802757263,
-1.41124510765076,
-1.41225266456604,
-1.41326069831848,
-1.41426920890808,
-1.41527807712555,
-1.41628754138947,
-1.41729748249054,
-1.41830790042877,
-1.41931867599487,
-1.42032992839813,
-1.42134165763855,
-1.42235374450684,
-1.42336642742157,
-1.42437946796417,
-1.42539310455322,
-1.42640709877014,
-1.42742156982422,
-1.42843663692474,
-1.42945206165314,
-1.43046808242798,
-1.43148446083069,
-1.43250119686127,
-1.43351840972900,
-1.43453621864319,
-1.43555438518524,
-1.43657302856445,
-1.43759214878082,
-1.43861174583435,
-1.43963181972504,
-1.44065237045288,
-1.44167339801788,
-1.44269490242004,
-1.44371688365936,
-1.44473922252655,
-1.44576203823090,
-1.44678533077240,
-1.44780910015106,
-1.44883334636688,
-1.44985795021057,
-1.45088315010071,
-1.45190882682800,
-1.45293498039246,
-1.45396149158478,
-1.45498859882355,
-1.45601606369019,
-1.45704388618469,
-1.45807230472565,
-1.45910108089447,
-1.46013033390045,
-1.46116018295288,
-1.46219038963318,
-1.46322119235992,
-1.46425235271454,
-1.46528410911560,
-1.46631622314453,
-1.46734881401062,
-1.46838176250458,
-1.46941530704498,
-1.47044920921326,
-1.47148358821869,
-1.47251844406128,
-1.47355377674103,
-1.47458958625793,
-1.47562587261200,
-1.47666263580322,
-1.47769987583160,
-1.47873771190643,
-1.47977566719055,
-1.48081421852112,
-1.48185324668884,
-1.48289275169373,
-1.48393273353577,
-1.48497307300568,
-1.48601400852203,
-1.48705542087555,
-1.48809731006622,
-1.48913955688477,
-1.49018239974976,
-1.49122571945190,
-1.49226927757263,
-1.49331343173981,
-1.49435794353485,
-1.49540305137634,
-1.49644851684570,
-1.49749457836151,
-1.49854099750519,
-1.49958789348602,
-1.50063538551331,
-1.50168323516846,
-1.50273168087006,
-1.50378036499023,
-1.50482952594757,
-1.50587904453278,
-1.50692903995514,
-1.50797951221466,
-1.50903046131134,
-1.51008176803589,
-1.51113367080688,
-1.51218605041504,
-1.51323890686035,
-1.51429224014282,
-1.51534605026245,
-1.51640009880066,
-1.51745474338532,
-1.51850986480713,
-1.51956534385681,
-1.52062141895294,
-1.52167785167694,
-1.52273488044739,
-1.52379226684570,
-1.52485024929047,
-1.52590858936310,
-1.52696752548218,
-1.52802670001984,
-1.52908647060394,
-1.53014659881592,
-1.53120720386505,
-1.53226828575134,
-1.53332984447479,
-1.53439199924469,
-1.53545451164246,
-1.53651750087738,
-1.53758096694946,
-1.53864502906799,
-1.53970932960510,
-1.54077398777008,
-1.54183924198151,
-1.54290497303009,
-1.54397118091583,
-1.54503786563873,
-1.54610502719879,
-1.54717266559601,
-1.54824078083038,
-1.54930937290192,
-1.55037844181061,
-1.55144774913788,
-1.55251765251160,
-1.55358791351318,
-1.55465877056122,
-1.55572998523712,
-1.55680179595947,
-1.55787408351898,
-1.55894672870636,
-1.56001996994019,
-1.56109356880188,
-1.56216776371002,
-1.56324231624603,
-1.56431734561920,
-1.56539273262024,
-1.56646859645844,
-1.56754493713379,
-1.56862187385559,
-1.56969916820526,
-1.57077693939209,
-1.57185518741608,
-1.57293403148651,
-1.57401323318481,
-1.57509291172028,
-1.57617294788361,
-1.57725346088409,
-1.57833445072174,
-1.57941591739655,
-1.58049786090851,
-1.58158028125763,
-1.58266305923462,
-1.58374643325806,
-1.58483028411865,
-1.58591461181641,
-1.58699941635132,
-1.58808457851410,
-1.58917009830475,
-1.59025621414185,
-1.59134268760681,
-1.59242975711823,
-1.59351718425751,
-1.59460520744324,
-1.59569370746613,
-1.59678256511688,
-1.59787201881409,
-1.59896183013916,
-1.60005211830139,
-1.60114276409149,
-1.60223388671875,
-1.60332548618317,
-1.60441756248474,
-1.60551023483276,
-1.60660326480865,
-1.60769677162170,
-1.60879075527191,
-1.60988533496857,
-1.61098015308380,
-1.61207532882690,
-1.61317110061646,
-1.61426734924316,
-1.61536407470703,
-1.61646127700806,
-1.61755895614624,
-1.61865711212158,
-1.61975574493408,
-1.62085485458374,
-1.62195432186127,
-1.62305426597595,
-1.62415468692780,
-1.62525546550751,
-1.62635684013367,
-1.62745857238770,
-1.62856090068817,
-1.62966358661652,
-1.63076686859131,
-1.63187050819397,
-1.63297474384308,
-1.63407933712006,
-1.63518440723419,
-1.63628983497620,
-1.63739573955536,
-1.63850212097168,
-1.63960909843445,
-1.64071643352509,
-1.64182424545288,
-1.64293253421783,
-1.64404129981995,
-1.64515066146851,
-1.64626038074493,
-1.64737045764923,
-1.64848089218140,
-1.64959192276001,
-1.65070343017578,
-1.65181541442871,
-1.65292787551880,
-1.65404081344605,
-1.65515410900116,
-1.65626800060272,
-1.65738236904144,
-1.65849721431732,
-1.65961241722107,
-1.66072797775269,
-1.66184413433075,
-1.66296064853668,
-1.66407775878906,
-1.66519522666931,
-1.66631317138672,
-1.66743171215057,
-1.66855061054230,
-1.66967010498047,
-1.67078983783722,
-1.67191004753113,
-1.67303073406219,
-1.67415201663971,
-1.67527365684509,
-1.67639577388763,
-1.67751836776733,
-1.67864143848419,
-1.67976498603821,
-1.68088901042938,
-1.68201351165771,
-1.68313837051392,
-1.68426370620728,
-1.68538951873779,
-1.68651580810547,
-1.68764245510101,
-1.68876969814301,
-1.68989741802216,
-1.69102561473846,
-1.69215416908264,
-1.69328331947327,
-1.69441294670105,
-1.69554281234741,
-1.69667327404022,
-1.69780409336090,
-1.69893538951874,
-1.70006728172302,
-1.70119953155518,
-1.70233237743378,
-1.70346558094025,
-1.70459926128387,
-1.70573353767395,
-1.70686805248261,
-1.70800304412842,
-1.70913851261139,
-1.71027445793152,
-1.71141088008881,
-1.71254777908325,
-1.71368515491486,
-1.71482300758362,
-1.71596133708954,
-1.71710014343262,
-1.71823942661285,
-1.71937906742096,
-1.72051906585693,
-1.72165966033936,
-1.72280073165894,
-1.72394216060638,
-1.72508418560028,
-1.72622668743134,
-1.72736954689026,
-1.72851300239563,
-1.72965693473816,
-1.73080110549927,
-1.73194575309753,
-1.73309087753296,
-1.73423647880554,
-1.73538267612457,
-1.73652923107147,
-1.73767626285553,
-1.73882377147675,
-1.73997187614441,
-1.74112033843994,
-1.74226915836334,
-1.74341845512390,
-1.74456822872162,
-1.74571835994720,
-1.74686908721924,
-1.74802029132843,
-1.74917197227478,
-1.75032413005829,
-1.75147676467896,
-1.75262987613678,
-1.75378334522247,
-1.75493729114532,
-1.75609159469605,
-1.75724649429321,
-1.75840175151825,
-1.75955760478973,
-1.76071381568909,
-1.76187062263489,
-1.76302778720856,
-1.76418542861938,
-1.76534366607666,
-1.76650214195251,
-1.76766109466553,
-1.76882052421570,
-1.76998043060303,
-1.77114081382751,
-1.77230167388916,
-1.77346301078796,
-1.77462482452393,
-1.77578711509705,
-1.77694988250732,
-1.77811300754547,
-1.77927660942078,
-1.78044056892395,
-1.78160512447357,
-1.78277003765106,
-1.78393554687500,
-1.78510153293610,
-1.78626787662506,
-1.78743481636047,
-1.78860223293304,
-1.78977000713348,
-1.79093813896179,
-1.79210686683655,
-1.79327595233917,
-1.79444551467896,
-1.79561555385590,
-1.79678606987000,
-1.79795718193054,
-1.79912865161896,
-1.80030059814453,
-1.80147302150726,
-1.80264580249786,
-1.80381906032562,
-1.80499279499054,
-1.80616688728333,
-1.80734157562256,
-1.80851674079895,
-1.80969238281250,
-1.81086838245392,
-1.81204497814178,
-1.81322205066681,
-1.81439936161041,
-1.81557726860046,
-1.81675553321838,
-1.81793427467346,
-1.81911361217499,
-1.82029330730438,
-1.82147347927094,
-1.82265424728394,
-1.82383537292480,
-1.82501697540283,
-1.82619893550873,
-1.82738125324249,
-1.82856392860413,
-1.82974720001221,
-1.83093094825745,
-1.83211505413055,
-1.83329975605011,
-1.83448493480682,
-1.83567047119141,
-1.83685660362244,
-1.83804297447205,
-1.83922982215881,
-1.84041726589203,
-1.84160506725311,
-1.84279334545136,
-1.84398210048676,
-1.84517133235931,
-1.84636116027832,
-1.84755134582520,
-1.84874200820923,
-1.84993302822113,
-1.85112440586090,
-1.85231637954712,
-1.85350883007050,
-1.85470175743103,
-1.85589504241943,
-1.85708892345428,
-1.85828328132629,
-1.85947811603546,
-1.86067330837250,
-1.86186897754669,
-1.86306500434875,
-1.86426150798798,
-1.86545848846436,
-1.86665606498718,
-1.86785399913788,
-1.86905241012573,
-1.87025129795074,
-1.87145078182220,
-1.87265062332153,
-1.87385082244873,
-1.87505137920380,
-1.87625253200531,
-1.87745416164398,
-1.87865626811981,
-1.87985873222351,
-1.88106179237366,
-1.88226532936096,
-1.88346934318542,
-1.88467383384705,
-1.88587856292725,
-1.88708376884460,
-1.88828945159912,
-1.88949573040009,
-1.89070236682892,
-1.89190948009491,
-1.89311695098877,
-1.89432489871979,
-1.89553332328796,
-1.89674222469330,
-1.89795148372650,
-1.89916110038757,
-1.90037131309509,
-1.90158188343048,
-1.90279304981232,
-1.90400457382202,
-1.90521669387817,
-1.90642929077148,
-1.90764224529266,
-1.90885579586029,
-1.91006958484650,
-1.91128385066986,
-1.91249859333038,
-1.91371381282806,
-1.91492950916290,
-1.91614568233490,
-1.91736233234406,
-1.91857945919037,
-1.91979706287384,
-1.92101514339447,
-1.92223346233368,
-1.92345237731934,
-1.92467164993286,
-1.92589151859283,
-1.92711174488068,
-1.92833256721497,
-1.92955374717712,
-1.93077552318573,
-1.93199765682220,
-1.93322014808655,
-1.93444311618805,
-1.93566656112671,
-1.93689036369324,
-1.93811464309692,
-1.93933928012848,
-1.94056451320648,
-1.94179022312164,
-1.94301640987396,
-1.94424295425415,
-1.94546985626221,
-1.94669735431671,
-1.94792520999908,
-1.94915354251862,
-1.95038235187531,
-1.95161163806915,
-1.95284152030945,
-1.95407176017761,
-1.95530247688293,
-1.95653367042542,
-1.95776522159576,
-1.95899713039398,
-1.96022963523865,
-1.96146261692047,
-1.96269595623016,
-1.96392989158630,
-1.96516418457031,
-1.96639907360077,
-1.96763443946838,
-1.96887004375458,
-1.97010612487793,
-1.97134268283844,
-1.97257959842682,
-1.97381687164307,
-1.97505474090576,
-1.97629308700562,
-1.97753190994263,
-1.97877120971680,
-1.98001098632813,
-1.98125100135803,
-1.98249149322510,
-1.98373246192932,
-1.98497390747070,
-1.98621594905853,
-1.98745834827423,
-1.98870122432709,
-1.98994457721710,
-1.99118852615356,
-1.99243283271790,
-1.99367749691010,
-1.99492251873016,
-1.99616813659668,
-1.99741411209106,
-1.99866068363190,
-1.99990773200989,
-2.00115513801575,
-2.00240278244019,
-2.00365114212036,
-2.00489974021912,
-2.00614881515503,
-2.00739836692810,
-2.00864839553833,
-2.00989866256714,
-2.01114964485168,
-2.01240110397339,
-2.01365303993225,
-2.01490545272827,
-2.01615834236145,
-2.01741147041321,
-2.01866507530212,
-2.01991915702820,
-2.02117371559143,
-2.02242875099182,
-2.02368450164795,
-2.02494049072266,
-2.02619671821594,
-2.02745366096497,
-2.02871060371399,
-2.02996826171875,
-2.03122639656067,
-2.03248476982117,
-2.03374385833740,
-2.03500342369080,
-2.03626322746277,
-2.03752374649048,
-2.03878474235535,
-2.04004597663879,
-2.04130768775940,
-2.04256987571716,
-2.04383254051209,
-2.04509568214417,
-2.04635906219482,
-2.04762315750122,
-2.04888749122620,
-2.05015254020691,
-2.05141782760620,
-2.05268335342407,
-2.05394959449768,
-2.05521607398987,
-2.05648326873779,
-2.05775070190430,
-2.05901861190796,
-2.06028723716736,
-2.06155610084534,
-2.06282544136047,
-2.06409549713135,
-2.06536555290222,
-2.06663632392883,
-2.06790757179260,
-2.06917905807495,
-2.07045078277588,
-2.07172322273254,
-2.07299613952637,
-2.07426953315735,
-2.07554340362549,
-2.07681751251221,
-2.07809209823608,
-2.07936739921570,
-2.08064293861389,
-2.08191895484924,
-2.08319544792175,
-2.08447241783142,
-2.08574986457825,
-2.08702778816223,
-2.08830595016480,
-2.08958435058594,
-2.09086346626282,
-2.09214305877686,
-2.09342288970947,
-2.09470343589783,
-2.09598445892334,
-2.09726572036743,
-2.09854769706726,
-2.09983015060425,
-2.10111260414124,
-2.10239577293396,
-2.10367941856384,
-2.10496330261230,
-2.10624766349793,
-2.10753250122070,
-2.10881805419922,
-2.11010384559631,
-2.11139011383057,
-2.11267662048340,
-2.11396384239197,
-2.11525130271912,
-2.11653923988342,
-2.11782765388489,
-2.11911678314209,
-2.12040615081787,
-2.12169599533081,
-2.12298607826233,
-2.12427663803101,
-2.12556767463684,
-2.12685918807983,
-2.12815117835999,
-2.12944364547730,
-2.13073635101318,
-2.13202977180481,
-2.13332366943359,
-2.13461804389954,
-2.13591265678406,
-2.13720750808716,
-2.13850283622742,
-2.13979887962341,
-2.14109516143799,
-2.14239192008972,
-2.14368939399719,
-2.14498710632324,
-2.14628529548645,
-2.14758419990540,
-2.14888310432434,
-2.15018272399902,
-2.15148234367371,
-2.15278267860413,
-2.15408349037170,
-2.15538477897644,
-2.15668654441834,
-2.15798878669739,
-2.15929126739502,
-2.16059422492981,
-2.16189765930176,
-2.16320157051086,
-2.16450595855713,
-2.16581058502197,
-2.16711568832397,
-2.16842150688171,
-2.16972756385803,
-2.17103409767151,
-2.17234110832214,
-2.17364835739136,
-2.17495608329773,
-2.17626452445984,
-2.17757320404053,
-2.17888236045837,
-2.18019175529480,
-2.18150186538696,
-2.18281245231628,
-2.18412327766418,
-2.18543457984924,
-2.18674635887146,
-2.18805861473084,
-2.18937110900879,
-2.19068431854248,
-2.19199776649475,
-2.19331169128418,
-2.19462633132935,
-2.19594097137451,
-2.19725608825684,
-2.19857192039490,
-2.19988799095154,
-2.20120477676392,
-2.20252156257629,
-2.20383906364441,
-2.20515704154968,
-2.20647549629211,
-2.20779395103455,
-2.20911312103272,
-2.21043276786804,
-2.21175289154053,
-2.21307349205017,
-2.21439433097839,
-2.21571564674377,
-2.21703743934631,
-2.21835994720459,
-2.21968245506287,
-2.22100543975830,
-2.22232913970947,
-2.22365307807922,
-2.22497749328613,
-2.22630238533020,
-2.22762751579285,
-2.22895336151123,
-2.23027968406677,
-2.23160624504089,
-2.23293304443359,
-2.23426055908203,
-2.23558855056763,
-2.23691678047180,
-2.23824548721313,
-2.23957467079163,
-2.24090433120728,
-2.24223446846008,
-2.24356508255005,
-2.24489593505859,
-2.24622726440430,
-2.24755907058716,
-2.24889111518860,
-2.25022387504578,
-2.25155687332153,
-2.25289058685303,
-2.25422453880310,
-2.25555896759033,
-2.25689363479614,
-2.25822877883911,
-2.25956439971924,
-2.26090049743652,
-2.26223707199097,
-2.26357412338257,
-2.26491165161133,
-2.26624965667725,
-2.26758766174316,
-2.26892638206482,
-2.27026534080505,
-2.27160501480103,
-2.27294492721558,
-2.27428531646729,
-2.27562642097473,
-2.27696776390076,
-2.27830934524536,
-2.27965140342712,
-2.28099393844605,
-2.28233695030212,
-2.28368043899536,
-2.28502440452576,
-2.28636860847473,
-2.28771352767944,
-2.28905868530273,
-2.29040431976318,
-2.29175019264221,
-2.29309678077698,
-2.29444360733032,
-2.29579091072083,
-2.29713869094849,
-2.29848670959473,
-2.29983544349670,
-2.30118465423584,
-2.30253410339355,
-2.30388402938843,
-2.30523419380188,
-2.30658483505249,
-2.30793595314026,
-2.30928754806519,
-2.31063961982727,
-2.31199216842651,
-2.31334519386292,
-2.31469821929932,
-2.31605195999146,
-2.31740593910217,
-2.31876063346863,
-2.32011556625366,
-2.32147121429443,
-2.32282710075378,
-2.32418346405029,
-2.32554030418396,
-2.32689714431763,
-2.32825469970703,
-2.32961273193359,
-2.33097124099731,
-2.33232998847961,
-2.33368921279907,
-2.33504891395569,
-2.33640933036804,
-2.33776998519897,
-2.33913087844849,
-2.34049224853516,
-2.34185409545898,
-2.34321618080139,
-2.34457898139954,
-2.34594202041626,
-2.34730577468872,
-2.34866976737976,
-2.35003423690796,
-2.35139894485474,
-2.35276412963867,
-2.35412979125977,
-2.35549592971802,
-2.35686254501343,
-2.35822939872742,
-2.35959696769714,
-2.36096477508545,
-2.36233282089233,
-2.36370134353638,
-2.36507058143616,
-2.36643981933594,
-2.36780977249146,
-2.36918020248413,
-2.37055087089539,
-2.37192225456238,
-2.37329411506653,
-2.37466597557068,
-2.37603831291199,
-2.37741112709045,
-2.37878441810608,
-2.38015818595886,
-2.38153243064880,
-2.38290691375732,
-2.38428211212158,
-2.38565754890442,
-2.38703322410584,
-2.38840961456299,
-2.38978600502014,
-2.39116311073303,
-2.39254069328308,
-2.39391875267029,
-2.39529705047607,
-2.39667606353760,
-2.39805507659912,
-2.39943456649780,
-2.40081453323364,
-2.40219497680664,
-2.40357589721680,
-2.40495729446411,
-2.40633893013001,
-2.40772128105164,
-2.40910387039185,
-2.41048693656921,
-2.41187024116516,
-2.41325402259827,
-2.41463828086853,
-2.41602277755737,
-2.41740798950195,
-2.41879367828369,
-2.42017960548401,
-2.42156600952148,
-2.42295265197754,
-2.42433977127075,
-2.42572736740112,
-2.42711544036865,
-2.42850399017334,
-2.42989277839661,
-2.43128228187561,
-2.43267202377319,
-2.43406224250793,
-2.43545246124268,
-2.43684339523315,
-2.43823480606079,
-2.43962669372559,
-2.44101905822754,
-2.44241166114807,
-2.44380474090576,
-2.44519829750061,
-2.44659209251404,
-2.44798636436462,
-2.44938111305237,
-2.45077610015869,
-2.45217156410217,
-2.45356774330139,
-2.45496416091919,
-2.45636105537415,
-2.45775818824768,
-2.45915555953980,
-2.46055340766907,
-2.46195197105408,
-2.46335077285767,
-2.46475028991699,
-2.46615004539490,
-2.46755003929138,
-2.46895074844360,
-2.47035169601440,
-2.47175312042236,
-2.47315478324890,
-2.47455692291260,
-2.47595953941345,
-2.47736263275147,
-2.47876644134522,
-2.48017024993897,
-2.48157429695129,
-2.48297905921936,
-2.48438405990601,
-2.48578977584839,
-2.48719573020935,
-2.48860192298889,
-2.49000883102417,
-2.49141621589661,
-2.49282360076904,
-2.49423170089722,
-2.49563980102539,
-2.49704885482788,
-2.49845790863037,
-2.49986767768860,
-2.50127768516541,
-2.50268816947937,
-2.50409936904907,
-2.50551056861877,
-2.50692200660706,
-2.50833415985107,
-2.50974678993225,
-2.51115965843201,
-2.51257324218750,
-2.51398682594299,
-2.51540136337280,
-2.51681590080261,
-2.51823067665100,
-2.51964616775513,
-2.52106189727783,
-2.52247810363770,
-2.52389478683472,
-2.52531194686890,
-2.52672958374023,
-2.52814745903015,
-2.52956581115723,
-2.53098440170288,
-2.53240323066711,
-2.53382301330566,
-2.53524279594421,
-2.53666305541992,
-2.53808403015137,
-2.53950500488281,
-2.54092693328857,
-2.54234886169434,
-2.54377102851868,
-2.54519391059876,
-2.54661703109741,
-2.54804039001465,
-2.54946470260620,
-2.55088901519775,
-2.55231404304504,
-2.55373930931091,
-2.55516457557678,
-2.55659079551697,
-2.55801701545715,
-2.55944418907166,
-2.56087160110474,
-2.56229925155640,
-2.56372737884522,
-2.56515574455261,
-2.56658458709717,
-2.56801390647888,
-2.56944346427918,
-2.57087373733521,
-2.57230424880981,
-2.57373523712158,
-2.57516670227051,
-2.57659864425659,
-2.57803058624268,
-2.57946300506592,
-2.58089590072632,
-2.58232927322388,
-2.58376288414001,
-2.58519721031189,
-2.58663201332092,
-2.58806705474854,
-2.58950209617615,
-2.59093785285950,
-2.59237408638001,
-2.59381055831909,
-2.59524750709534,
-2.59668493270874,
-2.59812307357788,
-2.59956121444702,
-2.60099959373474,
-2.60243868827820,
-2.60387802124023,
-2.60531783103943,
-2.60675811767578,
-2.60819864273071,
-2.60963964462280,
-2.61108112335205,
-2.61252307891846,
-2.61396527290344,
-2.61540794372559,
-2.61685085296631,
-2.61829423904419,
-2.61973810195923,
-2.62118220329285,
-2.62262701988220,
-2.62407231330872,
-2.62551736831665,
-2.62696313858032,
-2.62840938568115,
-2.62985610961914,
-2.63130307197571,
-2.63275051116943,
-2.63419866561890,
-2.63564682006836,
-2.63709521293640,
-2.63854432106018,
-2.63999366760254,
-2.64144349098206,
-2.64289379119873,
-2.64434432983398,
-2.64579558372498,
-2.64724707603455,
-2.64869880676270,
-2.65015101432800,
-2.65160369873047,
-2.65305662155151,
-2.65451002120972,
-2.65596389770508,
-2.65741801261902,
-2.65887284278870,
-2.66032791137695,
-2.66178321838379,
-2.66323900222778,
-2.66469502449036,
-2.66615152359009,
-2.66760849952698,
-2.66906595230103,
-2.67052388191223,
-2.67198228836060,
-2.67344069480896,
-2.67489981651306,
-2.67635917663574,
-2.67781877517700,
-2.67927908897400,
-2.68073964118958,
-2.68220067024231,
-2.68366217613220,
-2.68512368202209,
-2.68658566474915,
-2.68804836273193,
-2.68951106071472,
-2.69097447395325,
-2.69243812561035,
-2.69390225410461,
-2.69536685943604,
-2.69683170318604,
-2.69829678535461,
-2.69976234436035,
-2.70122838020325,
-2.70269489288330,
-2.70416164398193,
-2.70562887191772,
-2.70709657669067,
-2.70856428146362,
-2.71003270149231,
-2.71150135993958,
-2.71297049522400,
-2.71444010734558,
-2.71590995788574,
-2.71738028526306,
-2.71885108947754,
-2.72032213211060,
-2.72179341316223,
-2.72326540946960,
-2.72473764419556,
-2.72621011734009,
-2.72768330574036,
-2.72915673255920,
-2.73063063621521,
-2.73210477828980,
-2.73357915878296,
-2.73505401611328,
-2.73652935028076,
-2.73800516128540,
-2.73948121070862,
-2.74095797538757,
-2.74243497848511,
-2.74391198158264,
-2.74538969993591,
-2.74686765670776,
-2.74834609031677,
-2.74982500076294,
-2.75130438804626,
-2.75278401374817,
-2.75426411628723,
-2.75574445724487,
-2.75722503662109,
-2.75870633125305,
-2.76018786430359,
-2.76166963577271,
-2.76315212249756,
-2.76463484764099,
-2.76611804962158,
-2.76760172843933,
-2.76908564567566,
-2.77056956291199,
-2.77205443382263,
-2.77353954315186,
-2.77502489089966,
-2.77651095390320,
-2.77799725532532,
-2.77948379516602,
-2.78097081184387,
-2.78245806694031,
-2.78394579887390,
-2.78543400764465,
-2.78692269325256,
-2.78841137886047,
-2.78990101814270,
-2.79139089584351,
-2.79288077354431,
-2.79437088966370,
-2.79586172103882,
-2.79735302925110,
-2.79884433746338,
-2.80033659934998,
-2.80182886123657,
-2.80332159996033,
-2.80481481552124,
-2.80630803108215,
-2.80780196189880,
-2.80929613113403,
-2.81079077720642,
-2.81228590011597,
-2.81378149986267,
-2.81527733802795,
-2.81677341461182,
-2.81826972961426,
-2.81976652145386,
-2.82126379013062,
-2.82276129722595,
-2.82425951957703,
-2.82575798034668,
-2.82725691795349,
-2.82875609397888,
-2.83025550842285,
-2.83175516128540,
-2.83325576782227,
-2.83475637435913,
-2.83625745773315,
-2.83775877952576,
-2.83926057815552,
-2.84076261520386,
-2.84226512908936,
-2.84376811981201,
-2.84527134895325,
-2.84677505493164,
-2.84827923774719,
-2.84978365898132,
-2.85128831863403,
-2.85279321670532,
-2.85429883003235,
-2.85580468177795,
-2.85731101036072,
-2.85881781578064,
-2.86032485961914,
-2.86183238029480,
-2.86334013938904,
-2.86484813690186,
-2.86635661125183,
-2.86786532402039,
-2.86937475204468,
-2.87088441848755,
-2.87239456176758,
-2.87390518188477,
-2.87541580200195,
-2.87692666053772,
-2.87843799591064,
-2.87995004653931,
-2.88146233558655,
-2.88297486305237,
-2.88448786735535,
-2.88600158691406,
-2.88751506805420,
-2.88902878761292,
-2.89054346084595,
-2.89205813407898,
-2.89357328414917,
-2.89508914947510,
-2.89660501480103,
-2.89812159538269,
-2.89963793754578,
-2.90115499496460,
-2.90267229080200,
-2.90419006347656,
-2.90570831298828,
-2.90722680091858,
-2.90874576568604,
-2.91026496887207,
-2.91178464889526,
-2.91330456733704,
-2.91482472419739,
-2.91634559631348,
-2.91786670684814,
-2.91938829421997,
-2.92091012001038,
-2.92243242263794,
-2.92395496368408,
-2.92547774314880,
-2.92700099945068,
-2.92852473258972,
-2.93004894256592,
-2.93157315254211,
-2.93309807777405,
-2.93462324142456,
-2.93614840507507,
-2.93767404556274,
-2.93920040130615,
-2.94072699546814,
-2.94225382804871,
-2.94378137588501,
-2.94530916213989,
-2.94683694839478,
-2.94836521148682,
-2.94989395141602,
-2.95142316818237,
-2.95295262336731,
-2.95448231697083,
-2.95601272583008,
-2.95754337310791,
-2.95907425880432,
-2.96060514450073,
-2.96213674545288,
-2.96366882324219,
-2.96520113945007,
-2.96673393249512,
-2.96826720237732,
-2.96980071067810,
-2.97133445739746,
-2.97286868095398,
-2.97440314292908,
-2.97593784332275,
-2.97747302055359,
-2.97900891304016,
-2.98054504394531,
-2.98208141326904,
-2.98361778259277,
-2.98515486717224,
-2.98669219017029,
-2.98822999000549,
-2.98976778984070,
-2.99130654335022,
-2.99284553527832,
-2.99438452720642,
-2.99592375755310,
-2.99746370315552,
-2.99900388717651,
-3.00054430961609,
-3.00208520889282,
-3.00362682342529,
-3.00516843795776,
-3.00671029090881,
-3.00825238227844,
-3.00979518890381,
-3.01133823394775,
-3.01288175582886,
-3.01442527770996,
-3.01596975326538,
-3.01751422882080,
-3.01905894279480,
-3.02060389518738,
-3.02214956283569,
-3.02369546890259,
-3.02524161338806,
-3.02678823471069,
-3.02833533287048,
-3.02988290786743,
-3.03143048286438,
-3.03297829627991,
-3.03452658653259,
-3.03607535362244,
-3.03762459754944,
-3.03917384147644,
-3.04072380065918,
-3.04227399826050,
-3.04382419586182,
-3.04537487030029,
-3.04692625999451,
-3.04847788810730,
-3.05002975463867,
-3.05158185958862,
-3.05313444137573,
-3.05468750000000,
-3.05624055862427,
-3.05779409408569,
-3.05934786796570,
-3.06090235710144,
-3.06245708465576,
-3.06401205062866,
-3.06556749343872,
-3.06712317466736,
-3.06867933273315,
-3.07023549079895,
-3.07179212570190,
-3.07334947586060,
-3.07490706443787,
-3.07646489143372,
-3.07802295684814,
-3.07958102226257,
-3.08114004135132,
-3.08269906044006,
-3.08425855636597,
-3.08581852912903,
-3.08737874031067,
-3.08893966674805,
-3.09050035476685,
-3.09206128120422,
-3.09362268447876,
-3.09518480300903,
-3.09674715995789,
-3.09830975532532,
-3.09987258911133,
-3.10143613815308,
-3.10299968719482,
-3.10456371307373,
-3.10612773895264,
-3.10769248008728,
-3.10925745964050,
-3.11082291603088,
-3.11238861083984,
-3.11395454406738,
-3.11552071571350,
-3.11708736419678,
-3.11865425109863,
-3.12022161483765,
-3.12178945541382,
-3.12335753440857,
-3.12492609024048,
-3.12649488449097,
-3.12806367874146,
-3.12963294982910,
-3.13120269775391,
-3.13277292251587,
-3.13434338569641,
-3.13591432571411,
-3.13748502731323,
-3.13905644416809,
-3.14062809944153,
-3.14220023155212,
-3.14377260208130,
-3.14534521102905,
-3.14691853523254,
-3.14849209785461,
-3.15006589889526,
-3.15163969993591,
-3.15321397781372,
-3.15478897094727,
-3.15636396408081,
-3.15793943405151,
-3.15951538085938,
-3.16109156608582,
-3.16266798973084,
-3.16424465179443,
-3.16582179069519,
-3.16739916801453,
-3.16897678375244,
-3.17055511474609,
-3.17213368415833,
-3.17371225357056,
-3.17529129981995,
-3.17687058448792,
-3.17845034599304,
-3.18003058433533,
-3.18161106109619,
-3.18319177627563,
-3.18477296829224,
-3.18635439872742,
-3.18793606758118,
-3.18951821327209,
-3.19110059738159,
-3.19268321990967,
-3.19426655769348,
-3.19585013389587,
-3.19743394851685,
-3.19901776313782,
-3.20060205459595,
-3.20218658447266,
-3.20377182960510,
-3.20535731315613,
-3.20694303512573,
-3.20852923393250,
-3.21011519432068,
-3.21170210838318,
-3.21328902244568,
-3.21487641334534,
-3.21646404266357,
-3.21805214881897,
-3.21964049339294,
-3.22122907638550,
-3.22281789779663,
-3.22440719604492,
-3.22599673271179,
-3.22758650779724,
-3.22917699813843,
-3.23076772689819,
-3.23235893249512,
-3.23394989967346,
-3.23554134368897,
-3.23713326454163,
-3.23872542381287,
-3.24031805992126,
-3.24191117286682,
-3.24350428581238,
-3.24509763717651,
-3.24669122695923,
-3.24828553199768,
-3.24988007545471,
-3.25147485733032,
-3.25306987762451,
-3.25466537475586,
-3.25626111030579,
-3.25785732269287,
-3.25945353507996,
-3.26105022430420,
-3.26264739036560,
-3.26424455642700,
-3.26584219932556,
-3.26744055747986,
-3.26903867721558,
-3.27063727378845,
-3.27223610877991,
-3.27383542060852,
-3.27543473243713,
-3.27703499794006,
-3.27863526344299,
-3.28023600578308,
-3.28183674812317,
-3.28343772888184,
-3.28503918647766,
-3.28664088249207,
-3.28824305534363,
-3.28984570503235,
-3.29144859313965,
-3.29305148124695,
-3.29465460777283,
-3.29625821113586,
-3.29786229133606,
-3.29946660995483,
-3.30107140541077,
-3.30267643928528,
-3.30428147315979,
-3.30588698387146,
-3.30749249458313,
-3.30909895896912,
-3.31070542335510,
-3.31231236457825,
-3.31391954421997,
-3.31552720069885,
-3.31713461875916,
-3.31874251365662,
-3.32035088539124,
-3.32195973396301,
-3.32356882095337,
-3.32517814636230,
-3.32678794860840,
-3.32839751243591,
-3.33000755310059,
-3.33161807060242,
-3.33322906494141,
-3.33484029769897,
-3.33645176887512,
-3.33806371688843,
-3.33967590332031,
-3.34128785133362,
-3.34290075302124,
-3.34451389312744,
-3.34612727165222,
-3.34774088859558,
-3.34935498237610,
-3.35096907615662,
-3.35258340835571,
-3.35419821739197,
-3.35581326484680,
-3.35742878913879,
-3.35904479026794,
-3.36066079139709,
-3.36227726936340,
-3.36389374732971,
-3.36551046371460,
-3.36712765693665,
-3.36874532699585,
-3.37036323547363,
-3.37198162078857,
-3.37360024452209,
-3.37521910667419,
-3.37683796882629,
-3.37845730781555,
-3.38007688522339,
-3.38169693946838,
-3.38331747055054,
-3.38493824005127,
-3.38655924797058,
-3.38818025588989,
-3.38980174064636,
-3.39142322540283,
-3.39304542541504,
-3.39466786384583,
-3.39629077911377,
-3.39791393280029,
-3.39953756332397,
-3.40116095542908,
-3.40278482437134,
-3.40440893173218,
-3.40603351593018,
-3.40765810012817,
-3.40928363800049,
-3.41090917587280,
-3.41253495216370,
-3.41416072845459,
-3.41578698158264,
-3.41741371154785,
-3.41904044151306,
-3.42066764831543,
-3.42229509353638,
-3.42392277717590,
-3.42555069923401,
-3.42717909812927,
-3.42880797386169,
-3.43043684959412,
-3.43206620216370,
-3.43369579315186,
-3.43532586097717,
-3.43695569038391,
-3.43858599662781,
-3.44021654129028,
-3.44184756278992,
-3.44347906112671,
-3.44511079788208,
-3.44674301147461,
-3.44837498664856,
-3.45000743865967,
-3.45164012908936,
-3.45327305793762,
-3.45490622520447,
-3.45653986930847,
-3.45817399024963,
-3.45980834960938,
-3.46144270896912,
-3.46307754516602,
-3.46471261978149,
-3.46634817123413,
-3.46798372268677,
-3.46961975097656,
-3.47125577926636,
-3.47289204597473,
-3.47452878952026,
-3.47616600990295,
-3.47780346870422,
-3.47944140434265,
-3.48107957839966,
-3.48271799087524,
-3.48435640335083,
-3.48599505424500,
-3.48763418197632,
-3.48927354812622,
-3.49091315269470,
-3.49255323410034,
-3.49419355392456,
-3.49583363533020,
-3.49747443199158,
-3.49911570549011,
-3.50075721740723,
-3.50239896774292,
-3.50404095649719,
-3.50568342208862,
-3.50732588768005,
-3.50896835327148,
-3.51061153411865,
-3.51225471496582,
-3.51389837265015,
-3.51554226875305,
-3.51718640327454,
-3.51883101463318,
-3.52047562599182,
-3.52212071418762,
-3.52376627922058,
-3.52541184425354,
-3.52705788612366,
-3.52870416641235,
-3.53035092353821,
-3.53199744224548,
-3.53364443778992,
-3.53529167175293,
-3.53693914413452,
-3.53858685493469,
-3.54023504257202,
-3.54188346862793,
-3.54353189468384,
-3.54518055915833,
-3.54682993888855,
-3.54847955703735,
-3.55012941360474,
-3.55177974700928,
-3.55343031883240,
-3.55508065223694,
-3.55673146247864,
-3.55838251113892,
-3.56003403663635,
-3.56168580055237,
-3.56333780288696,
-3.56499004364014,
-3.56664252281189,
-3.56829500198364,
-3.56994795799255,
-3.57160115242004,
-3.57325482368469,
-3.57490849494934,
-3.57656264305115,
-3.57821750640869,
-3.57987213134766,
-3.58152723312378,
-3.58318257331848,
-3.58483815193176,
-3.58649396896362,
-3.58815026283264,
-3.58980679512024,
-3.59146332740784,
-3.59312009811401,
-3.59477710723877,
-3.59643459320068,
-3.59809231758118,
-3.59975028038025,
-3.60140872001648,
-3.60306692123413,
-3.60472559928894,
-3.60638451576233,
-3.60804367065430,
-3.60970330238342,
-3.61136293411255,
-3.61302304267883,
-3.61468315124512,
-3.61634349822998,
-3.61800432205200,
-3.61966538429260,
-3.62132668495178,
-3.62298846244812,
-3.62465071678162,
-3.62631273269653,
-3.62797522544861,
-3.62963795661926,
-3.63130116462708,
-3.63296461105347,
-3.63462829589844,
-3.63629221916199,
-3.63795638084412,
-3.63962078094482,
-3.64128518104553,
-3.64295005798340,
-3.64461541175842,
-3.64628076553345,
-3.64794659614563,
-3.64961266517639,
-3.65127873420715,
-3.65294504165649,
-3.65461158752441,
-3.65627861022949,
-3.65794587135315,
-3.65961337089539,
-3.66128110885620,
-3.66294908523560,
-3.66461706161499,
-3.66628551483154,
-3.66795420646668,
-3.66962313652039,
-3.67129254341126,
-3.67296218872070,
-3.67463183403015,
-3.67630171775818,
-3.67797183990479,
-3.67964220046997,
-3.68131303787231,
-3.68298411369324,
-3.68465566635132,
-3.68632698059082,
-3.68799853324890,
-3.68967056274414,
-3.69134283065796,
-3.69301533699036,
-3.69468808174133,
-3.69636130332947,
-3.69803452491760,
-3.69970798492432,
-3.70138168334961,
-3.70305562019348,
-3.70473003387451,
-3.70640468597412,
-3.70807957649231,
-3.70975446701050,
-3.71142959594727,
-3.71310496330261,
-3.71478080749512,
-3.71645689010620,
-3.71813321113586,
-3.71981000900269,
-3.72148704528809,
-3.72316384315491,
-3.72484111785889,
-3.72651863098145,
-3.72819662094116,
-3.72987461090088,
-3.73155307769775,
-3.73323178291321,
-3.73491048812866,
-3.73658967018127,
-3.73826885223389,
-3.73994851112366,
-3.74162840843201,
-3.74330854415894,
-3.74498915672302,
-3.74666953086853,
-3.74835014343262,
-3.75003123283386,
-3.75171256065369,
-3.75339436531067,
-3.75507616996765,
-3.75675845146179,
-3.75844073295593,
-3.76012325286865,
-3.76180577278137,
-3.76348853111267,
-3.76517152786255,
-3.76685500144959,
-3.76853871345520,
-3.77022242546082,
-3.77190637588501,
-3.77359056472778,
-3.77527523040772,
-3.77695989608765,
-3.77864503860474,
-3.78033065795898,
-3.78201603889465,
-3.78370165824890,
-3.78538775444031,
-3.78707408905029,
-3.78876066207886,
-3.79044747352600,
-3.79213476181030,
-3.79382181167603,
-3.79550909996033,
-3.79719686508179,
-3.79888486862183,
-3.80057334899902,
-3.80226182937622,
-3.80395078659058,
-3.80563974380493,
-3.80732870101929,
-3.80901789665222,
-3.81070733070374,
-3.81239700317383,
-3.81408715248108,
-3.81577754020691,
-3.81746768951416,
-3.81915831565857,
-3.82084918022156,
-3.82254052162170,
-3.82423210144043,
-3.82592391967773,
-3.82761597633362,
-3.82930803298950,
-3.83100032806397,
-3.83269286155701,
-3.83438587188721,
-3.83607912063599,
-3.83777236938477,
-3.83946585655212,
-3.84115934371948,
-3.84285306930542,
-3.84454703330994,
-3.84624147415161,
-3.84793615341187,
-3.84963107109070,
-3.85132646560669,
-3.85302162170410,
-3.85471701622009,
-3.85641288757324,
-3.85810899734497,
-3.85980534553528,
-3.86150193214417,
-3.86319899559021,
-3.86489558219910,
-3.86659264564514,
-3.86828970909119,
-3.86998724937439,
-3.87168502807617,
-3.87338328361511,
-3.87508153915405,
-3.87677979469299,
-3.87847852706909,
-3.88017749786377,
-3.88187670707703,
-3.88357615470886,
-3.88527607917786,
-3.88697576522827,
-3.88867568969727,
-3.89037561416626,
-3.89207601547241,
-3.89377665519714,
-3.89547753334045,
-3.89717888832092,
-3.89888024330139,
-3.90058183670044,
-3.90228366851807,
-3.90398573875427,
-3.90568804740906,
-3.90739035606384,
-3.90909290313721,
-3.91079592704773,
-3.91249871253967,
-3.91420197486877,
-3.91590547561646,
-3.91760921478272,
-3.91931319236755,
-3.92101764678955,
-3.92272233963013,
-3.92442679405212,
-3.92613148689270,
-3.92783617973328,
-3.92954134941101,
-3.93124699592590,
-3.93295264244080,
-3.93465876579285,
-3.93636465072632,
-3.93807101249695,
-3.93977761268616,
-3.94148445129395,
-3.94319128990173,
-3.94489836692810,
-3.94660592079163,
-3.94831323623657,
-3.95002102851868,
-3.95172882080078,
-3.95343708992004,
-3.95514583587647,
-3.95685458183289,
-3.95856356620789,
-3.96027231216431,
-3.96198129653931,
-3.96369075775147,
-3.96540045738220,
-3.96711039543152,
-3.96882057189941,
-3.97053122520447,
-3.97224164009094,
-3.97395205497742,
-3.97566270828247,
-3.97737383842468,
-3.97908520698547,
-3.98079681396484,
-3.98250889778137,
-3.98422074317932,
-3.98593282699585,
-3.98764491081238,
-3.98935747146606,
-3.99107027053833,
-3.99278306961060,
-3.99449658393860,
-3.99620985984802,
-3.99792337417603,
-3.99963712692261,
-4.00135087966919,
-4.00306510925293,
-4.00477933883667,
-4.00649404525757,
-4.00820875167847,
-4.00992393493652,
-4.01163911819458,
-4.01335430145264,
-4.01506996154785,
-4.01678562164307,
-4.01850175857544,
-4.02021789550781,
-4.02193403244019,
-4.02365064620972,
-4.02536773681641,
-4.02708482742310,
-4.02880191802979,
-4.03051948547363,
-4.03223705291748,
-4.03395462036133,
-4.03567266464233,
-4.03739070892334,
-4.03910923004150,
-4.04082775115967,
-4.04254674911499,
-4.04426574707031,
-4.04598474502564,
-4.04770374298096,
-4.04942369461060,
-4.05114364624023,
-4.05286359786987,
-4.05458354949951,
-4.05630397796631,
-4.05802440643311,
-4.05974483489990,
-4.06146574020386,
-4.06318712234497,
-4.06490802764893,
-4.06662988662720,
-4.06835126876831,
-4.07007312774658,
-4.07179498672485,
-4.07351732254028,
-4.07524013519287,
-4.07696247100830,
-4.07868576049805,
-4.08040857315064,
-4.08213138580322,
-4.08385515213013,
-4.08557844161987,
-4.08730220794678,
-4.08902597427368,
-4.09075069427490,
-4.09247446060181,
-4.09419918060303,
-4.09592390060425,
-4.09764862060547,
-4.09937381744385,
-4.10109901428223,
-4.10282468795776,
-4.10455036163330,
-4.10627555847168,
-4.10800170898438,
-4.10972785949707,
-4.11145401000977,
-4.11318111419678,
-4.11490821838379,
-4.11663484573364,
-4.11836147308350,
-4.12008857727051,
-4.12181615829468,
-4.12354421615601,
-4.12527179718018,
-4.12699937820435,
-4.12872743606567,
-4.13045597076416,
-4.13218450546265,
-4.13391304016113,
-4.13564205169678,
-4.13737106323242,
-4.13910007476807,
-4.14082956314087,
-4.14255905151367,
-4.14428853988648,
-4.14601850509644,
-4.14774894714356,
-4.14947938919067,
-4.15120983123779,
-4.15294027328491,
-4.15467119216919,
-4.15640211105347,
-4.15813302993774,
-4.15986490249634,
-4.16159629821777,
-4.16332769393921,
-4.16505956649780,
-4.16679143905640,
-4.16852378845215,
-4.17025661468506,
-4.17198896408081,
-4.17372179031372,
-4.17545461654663,
-4.17718744277954,
-4.17892122268677,
-4.18065452575684,
-4.18238782882690,
-4.18412208557129,
-4.18585586547852,
-4.18759012222290,
-4.18932437896729,
-4.19105863571167,
-4.19279336929321,
-4.19452810287476,
-4.19626331329346,
-4.19799852371216,
-4.19973373413086,
-4.20146894454956,
-4.20320463180542,
-4.20494079589844,
-4.20667695999146,
-4.20841312408447,
-4.21014976501465,
-4.21188592910767,
-4.21362257003784,
-4.21535921096802,
-4.21709632873535,
-4.21883344650269,
-4.22057104110718,
-4.22230815887451,
-4.22404575347900,
-4.22578334808350,
-4.22752141952515,
-4.22925949096680,
-4.23099803924561,
-4.23273658752441,
-4.23447513580322,
-4.23621368408203,
-4.23795270919800,
-4.23969173431397,
-4.24143075942993,
-4.24317073822022,
-4.24491024017334,
-4.24664974212647,
-4.24838924407959,
-4.25012969970703,
-4.25186967849731,
-4.25361013412476,
-4.25535106658936,
-4.25709199905396,
-4.25883245468140,
-4.26057338714600,
-4.26231479644775,
-4.26405620574951,
-4.26579761505127,
-4.26753950119019,
-4.26928138732910,
-4.27102327346802,
-4.27276515960693,
-4.27450752258301,
-4.27624988555908,
-4.27799224853516,
-4.27973556518555,
-4.28147840499878,
-4.28322124481201,
-4.28496456146240,
-4.28670787811279,
-4.28845167160034,
-4.29019546508789,
-4.29193925857544,
-4.29368352890015,
-4.29542779922485,
-4.29717206954956,
-4.29891633987427,
-4.30066108703613,
-4.30240583419800,
-4.30415105819702,
-4.30589580535889,
-4.30764102935791,
-4.30938625335693,
-4.31113195419312,
-4.31287765502930,
-4.31462335586548,
-4.31636953353882,
-4.31811523437500,
-4.31986141204834,
-4.32160758972168,
-4.32335424423218,
-4.32510089874268,
-4.32684803009033,
-4.32859516143799,
-4.33034181594849,
-4.33208894729614,
-4.33383655548096,
-4.33558416366577,
-4.33733177185059,
-4.33907985687256,
-4.34082794189453,
-4.34257650375366,
-4.34432458877564,
-4.34607267379761,
-4.34782123565674,
-4.34957027435303,
-4.35131931304932,
-4.35306835174561,
-4.35481739044189,
-4.35656642913818,
-4.35831594467163,
-4.36006546020508,
-4.36181545257568,
-4.36356544494629,
-4.36531591415405,
-4.36706590652466,
-4.36881589889526,
-4.37056636810303,
-4.37231683731079,
-4.37406778335571,
-4.37581872940064,
-4.37756967544556,
-4.37932062149048,
-4.38107156753540,
-4.38282299041748,
-4.38457441329956,
-4.38632678985596,
-4.38807868957520,
-4.38983011245728,
-4.39158248901367,
-4.39333438873291,
-4.39508676528931,
-4.39683914184570,
-4.39859199523926,
-4.40034484863281,
-4.40209722518921,
-4.40385055541992,
-4.40560340881348,
-4.40735673904419,
-4.40911006927490,
-4.41086387634277,
-4.41261768341064,
-4.41437149047852,
-4.41612529754639,
-4.41787910461426,
-4.41963338851929,
-4.42138767242432,
-4.42314243316650,
-4.42489719390869,
-4.42665195465088,
-4.42840671539307,
-4.43016147613525,
-4.43191671371460,
-4.43367195129395,
-4.43542718887329,
-4.43718290328980,
-4.43893814086914,
-4.44069337844849,
-4.44244956970215,
-4.44420576095581,
-4.44596195220947,
-4.44771814346314,
-4.44947481155396,
-4.45123100280762,
-4.45298767089844,
-4.45474433898926,
-4.45650100708008,
-4.45825815200806,
-4.46001577377319,
-4.46177244186401,
-4.46353006362915,
-4.46528720855713,
-4.46704483032227,
-4.46880245208740,
-4.47056055068970,
-4.47231864929199,
-4.47407674789429,
-4.47583484649658,
-4.47759294509888,
-4.47935152053833,
-4.48111009597778,
-4.48286914825439,
-4.48462772369385,
-4.48638629913330,
-4.48814535140991,
-4.48990440368652,
-4.49166393280029,
-4.49342298507690,
-4.49518299102783,
-4.49694252014160,
-4.49870157241821,
-4.50046157836914,
-4.50222158432007,
-4.50398159027100,
-4.50574207305908,
-4.50750255584717,
-4.50926256179810,
-4.51102304458618,
-4.51278400421143,
-4.51454448699951,
-4.51630544662476,
-4.51806688308716,
-4.51982831954956,
-4.52158927917481,
-4.52335023880005,
-4.52511167526245,
-4.52687311172485,
-4.52863502502441,
-4.53039693832398,
-4.53215885162354,
-4.53392076492310,
-4.53568267822266,
-4.53744506835938,
-4.53920745849609,
-4.54096984863281,
-4.54273271560669,
-4.54449510574341,
-4.54625749588013,
-4.54802036285400,
-4.54978322982788,
-4.55154657363892,
-4.55330944061279,
-4.55507326126099,
-4.55683660507202,
-4.55859947204590,
-4.56036329269409,
-4.56212711334229,
-4.56389093399048,
-4.56565523147583,
-4.56741905212402,
-4.56918287277222,
-4.57094717025757,
-4.57271146774292,
-4.57447576522827,
-4.57624053955078,
-4.57800531387329,
-4.57977056503296,
-4.58153486251831,
-4.58329963684082,
-4.58506488800049,
-4.58683013916016,
-4.58859539031982,
-4.59036064147949,
-4.59212589263916,
-4.59389114379883,
-4.59565687179565,
-4.59742259979248,
-4.59918832778931,
-4.60095453262329,
-4.60272073745728,
-4.60448646545410,
-4.60625267028809,
-4.60801887512207,
-4.60978507995606,
-4.61155176162720,
-4.61331844329834,
-4.61508512496948,
-4.61685180664063,
-4.61861848831177,
-4.62038564682007,
-4.62215280532837,
-4.62391996383667,
-4.62568712234497,
-4.62745475769043,
-4.62922191619873,
-4.63098955154419,
-4.63275671005249,
-4.63452482223511,
-4.63629245758057,
-4.63806056976318,
-4.63982820510864,
-4.64159631729126,
-4.64336442947388,
-4.64513254165649,
-4.64690113067627,
-4.64866924285889,
-4.65043830871582,
-4.65220642089844,
-4.65397500991821,
-4.65574359893799,
-4.65751266479492,
-4.65928173065186,
-4.66105031967163,
-4.66281986236572,
-4.66458892822266,
-4.66635799407959,
-4.66812753677368,
-4.66989660263062,
-4.67166662216187,
-4.67343616485596,
-4.67520570755005,
-4.67697572708130,
-4.67874526977539,
-4.68051528930664,
-4.68228530883789,
-4.68405532836914,
-4.68582582473755,
-4.68759584426880,
-4.68936586380005,
-4.69113636016846,
-4.69290685653687,
-4.69467735290527,
-4.69644832611084,
-4.69821882247925,
-4.69998979568481,
-4.70176029205322,
-4.70353126525879,
-4.70530223846436,
-4.70707321166992,
-4.70884466171265,
-4.71061611175537,
-4.71238756179810,
-4.71415853500366,
-4.71592998504639,
-4.71770143508911,
-4.71947288513184,
-4.72124528884888,
-4.72301673889160,
-4.72478818893433,
-4.72656011581421,
-4.72833204269409,
-4.73010396957398,
-4.73187637329102,
-4.73364877700806,
-4.73542070388794,
-4.73719310760498,
-4.73896551132202,
-4.74073791503906,
-4.74251031875610,
-4.74428319931030,
-4.74605607986450,
-4.74782896041870,
-4.74960136413574,
-4.75137424468994,
-4.75314712524414,
-4.75492048263550,
-4.75669336318970,
-4.75846672058106,
-4.76023960113525,
-4.76201295852661,
-4.76378631591797,
-4.76555967330933,
-4.76733350753784,
-4.76910734176636,
-4.77088069915772,
-4.77265405654907,
-4.77442789077759,
-4.77620172500610,
-4.77797555923462,
-4.77974987030029,
-4.78152418136597,
-4.78329753875732,
-4.78507184982300,
-4.78684568405151,
-4.78861999511719,
-4.79039430618286,
-4.79216861724854,
-4.79394340515137,
-4.79571771621704,
-4.79749202728272,
-4.79926633834839,
-4.80104112625122,
-4.80281591415405,
-4.80459070205689,
-4.80636548995972,
-4.80814027786255,
-4.80991506576538,
-4.81169033050537,
-4.81346511840820,
-4.81524085998535,
-4.81701612472534,
-4.81879091262817,
-4.82056617736816,
-4.82234144210815,
-4.82411718368530,
-4.82589244842529,
-4.82766819000244,
-4.82944393157959,
-4.83121919631958,
-4.83299446105957,
-4.83477020263672,
-4.83654594421387,
-4.83832168579102,
-4.84009742736816,
-4.84187364578247,
-4.84364938735962,
-4.84542512893677,
-4.84720134735107,
-4.84897708892822,
-4.85075330734253,
-4.85253000259399,
-4.85430574417114,
-4.85608196258545,
-4.85785818099976,
-4.85963439941406,
-4.86141061782837,
-4.86318731307983,
-4.86496400833130,
-4.86674070358276,
-4.86851692199707,
-4.87029361724854,
-4.87207031250000,
-4.87384700775147,
-4.87562417984009,
-4.87740135192871,
-4.87917804718018,
-4.88095474243164,
-4.88273143768311,
-4.88450860977173,
-4.88628578186035,
-4.88806247711182,
-4.88984012603760,
-4.89161682128906,
-4.89339399337769,
-4.89517116546631,
-4.89694881439209,
-4.89872598648071,
-4.90050363540649,
-4.90228080749512,
-4.90405797958374,
-4.90583562850952,
-4.90761280059814,
-4.90939044952393,
-4.91116809844971,
-4.91294574737549,
-4.91472339630127,
-4.91650104522705,
-4.91827869415283,
-4.92005634307861,
-4.92183446884155,
-4.92361211776733,
-4.92539024353027,
-4.92716789245606,
-4.92894554138184,
-4.93072366714478,
-4.93250131607056,
-4.93427944183350,
-4.93605756759644,
-4.93783569335938,
-4.93961381912231,
-4.94139146804810,
-4.94316959381104,
-4.94494771957398,
-4.94672632217407,
-4.94850492477417,
-4.95028305053711,
-4.95206069946289,
-4.95383882522583,
-4.95561742782593,
-4.95739603042603,
-4.95917463302612,
-4.96095275878906,
-4.96273088455200,
-4.96450948715210,
-4.96628808975220,
-4.96806621551514,
-4.96984481811523,
-4.97162389755249,
-4.97340250015259,
-4.97518062591553,
-4.97695922851563,
-4.97873735427856,
-4.98051643371582,
-4.98229551315308,
-4.98407459259033,
-4.98585271835327,
-4.98763132095337,
-4.98940992355347,
-4.99118900299072,
-4.99296760559082,
-4.99474668502808,
-4.99652528762817,
-4.99830436706543,
-5.00008296966553,
-5.00186204910278,
-5.00364065170288,
-5.00541973114014,
-5.00719881057739,
-5.00897836685181,
-5.01075696945190,
-5.01253557205200,
-5.01431465148926,
-5.01609373092651,
-5.01787281036377,
-5.01965236663818,
-5.02143096923828,
-5.02320957183838,
-5.02498865127564,
-5.02676820755005,
-5.02854728698731,
-5.03032636642456,
-5.03210544586182,
-5.03388452529907,
-5.03566360473633,
-5.03744268417358,
-5.03922176361084,
-5.04100084304810,
-5.04278087615967,
-5.04456043243408,
-5.04633951187134,
-5.04811811447144,
-5.04989719390869,
-5.05167627334595,
-5.05345582962036,
-5.05523538589478,
-5.05701446533203,
-5.05879306793213,
-5.06057214736939,
-5.06235170364380,
-5.06413125991821,
-5.06591033935547,
-5.06768989562988,
-5.06946897506714,
-5.07124805450439,
-5.07302761077881,
-5.07480716705322,
-5.07658624649048,
-5.07836580276489,
-5.08014488220215,
-5.08192396163940,
-5.08370351791382,
-5.08548259735107,
-5.08726215362549,
-5.08904123306274,
-5.09082078933716,
-5.09260034561157,
-5.09437942504883,
-5.09615850448608,
-5.09793758392334,
-5.09971666336060,
-5.10149621963501,
-5.10327625274658,
-5.10505533218384,
-5.10683441162109,
-5.10861301422119,
-5.11039209365845,
-5.11217164993286,
-5.11395120620728,
-5.11573076248169,
-5.11750984191895,
-5.11928892135620,
-5.12106752395630,
-5.12284708023071,
-5.12462663650513,
-5.12640571594238,
-5.12818527221680,
-5.12996387481689,
-5.13174295425415,
-5.13352203369141,
-5.13530158996582,
-5.13708066940308,
-5.13886022567749,
-5.14063882827759,
-5.14241743087769,
-5.14419651031494,
-5.14597606658936,
-5.14775514602661,
-5.14953422546387,
-5.15131330490112,
-5.15309190750122,
-5.15487098693848,
-5.15665006637573,
-5.15842914581299,
-5.16020822525024,
-5.16198730468750,
-5.16376590728760,
-5.16554498672485,
-5.16732406616211,
-5.16910314559937,
-5.17088174819946,
-5.17266082763672,
-5.17443943023682,
-5.17621803283691,
-5.17799663543701,
-5.17977571487427,
-5.18155431747437,
-5.18333292007446,
-5.18511152267456,
-5.18689060211182,
-5.18866920471191,
-5.19044780731201,
-5.19222640991211,
-5.19400501251221,
-5.19578361511231,
-5.19756221771240,
-5.19934082031250,
-5.20111942291260,
-5.20289802551270,
-5.20467615127564,
-5.20645475387573,
-5.20823335647583,
-5.21001148223877,
-5.21178960800171,
-5.21356773376465,
-5.21534633636475,
-5.21712446212769,
-5.21890258789063,
-5.22068119049072,
-5.22245931625366,
-5.22423696517944,
-5.22601509094238,
-5.22779846191406,
-5.23049259185791,
-5.23128509521484,
-5.23532867431641,
-5.23456478118897,
-5.24057531356812,
-5.23722219467163,
-5.24134778976440,
-5.23859834671021,
-5.23510694503784,
-5.23889064788818,
-5.21802043914795,
-5.23799991607666,
-5.18568801879883,
-5.23689317703247,
-5.13208770751953,
-5.23012447357178,
-5.14520883560181,
-5.25729274749756,
-5.11474180221558,
-5.28632688522339,
-5.09200954437256,
-5.42192268371582,
-5.08283662796021,
-5.25474309921265,
-5.00170660018921,
-5.35484743118286,
-5.25959491729736,
-5.20737934112549,
-5.86766290664673,
-5.03213834762573,
-6.69971656799316,
-4.97603464126587,
-6.51251840591431,
-5.12299919128418,
-7.13586759567261,
-5.53422832489014,
-7.90243721008301,
-6.41802453994751,
-10.6019515991211,
-6.82497549057007,
33.1978225708008,
-9.66641521453857,
-37.5254058837891,
-14.8991260528564,
-3.79583954811096,
16.4838237762451,
13.4833536148071,
59.7543601989746,
40.5096168518066,
-19.3894863128662,
-0.429540872573853,
-0.961202561855316,
-17.1116428375244,
-17.3420219421387,
-66.8547592163086,
0.972260117530823,
73.3756713867188,
-54.4821701049805,
-19.7678146362305,
7.01152896881104,
2.67027688026428,
5.94766902923584,
-17.6949539184570,
39.1751213073731,
-33.6451759338379,
29.4297695159912,
15.6194610595703,
-64.2730407714844,
-18.9644069671631,
-13.5047531127930,
-18.5988464355469,
-64.5209350585938,
51.0063514709473,
38.1700477600098,
-40.2093505859375,
49.0820236206055,
38.0025749206543,
-28.0351905822754,
-67.2158966064453,
-8.68502998352051,
-22.0369567871094,
-18.2142848968506,
44.5766601562500,
-53.7355499267578,
-37.3336334228516,
6.16938638687134,
-43.6734352111816,
-5.80642604827881,
22.7053699493408,
-29.8952178955078,
0.0637274980545044,
60.6618537902832,
25.2705345153809,
50.1082801818848,
59.9894104003906,
67.0321884155273,
40.4744186401367,
-33.3396148681641,
-20.5240573883057,
6.88310050964356,
18.1657409667969,
18.5009326934814,
78.8490753173828,
-16.0670452117920,
5.90121889114380,
65.7405548095703,
-72.9150314331055,
12.0054378509521,
33.7683258056641,
35.3321456909180,
14.2086057662964,
-24.2394866943359,
58.5855484008789,
-21.4226398468018,
-60.3691940307617,
-14.7555904388428,
3.00824189186096,
63.7593498229981,
7.74946308135986,
-54.6538314819336,
36.1558189392090,
15.9385290145874,
-38.9520187377930,
-2.80210876464844,
38.8286933898926,
30.5303115844727,
-27.3159065246582,
37.4168357849121,
-14.2492017745972,
-28.4515838623047,
56.2191276550293,
-35.2391090393066,
36.3062973022461,
29.3300781250000,
-48.0863838195801,
6.66316270828247,
-45.9831008911133,
-9.54656696319580,
78.7801742553711,
-2.05814290046692,
5.02997732162476,
26.6008892059326,
-49.9871788024902,
19.4818897247314,
33.9472351074219,
31.7115097045898,
32.9484596252441,
-16.8051242828369,
8.64315605163574,
-12.9996089935303,
25.9124317169189,
42.7756996154785,
-56.7802047729492,
43.7423095703125,
36.6373214721680,
-25.3397731781006,
57.8327789306641,
-39.4388275146484,
-17.3328189849854,
11.9537668228149,
-56.9870147705078,
-18.8904743194580,
88.0877761840820,
-2.13946318626404,
-38.3947219848633,
77.9635848999023,
-2.57099175453186,
34.5604019165039,
4.11260557174683,
-17.4170207977295,
59.4251556396484,
53.6906356811523,
-16.2721595764160,
-4.71926879882813,
23.2015838623047,
-64.9056015014648,
-33.9311180114746,
8.04700469970703,
35.8909606933594,
11.4700918197632,
20.8073921203613,
-12.1971912384033,
5.06617641448975,
12.3197898864746,
-45.2749557495117,
19.5522651672363,
-28.3042926788330,
-12.2026729583740,
-11.5550928115845,
26.7808971405029,
54.1720733642578,
-13.5157051086426,
67.9375305175781,
-11.7539358139038,
-27.0390090942383,
108.141288757324,
-6.57281351089478,
-44.7432250976563,
-13.9304342269897,
-1.75268125534058,
60.6490516662598,
20.8220462799072,
32.7565994262695,
44.9942283630371,
-12.0255784988403,
-69.4570693969727,
29.3226871490479,
9.76781272888184,
-45.1487159729004,
77.9070053100586,
3.53256869316101,
-24.3467922210693,
6.69786548614502,
-3.13764762878418,
11.4549312591553,
9.33519554138184,
37.9603500366211,
56.0392532348633,
-8.76451969146729,
21.0510768890381,
40.3092269897461,
-65.6785888671875,
34.6200752258301,
64.3350524902344,
11.0666713714600,
-14.3659162521362,
-44.0153121948242,
54.7746582031250,
-11.6997985839844,
-77.0076599121094,
27.8728389739990,
56.2644767761231,
-1.79159808158875,
21.9306678771973,
-38.7388114929199,
-35.5281791687012,
70.0832748413086,
-67.6559829711914,
46.2323913574219,
40.3242073059082,
-14.7781829833984,
38.1171836853027,
-60.6582031250000,
23.2172107696533,
-3.20177030563355,
46.4551315307617,
1.56185710430145,
-14.8003559112549,
56.4831695556641,
-32.7735824584961,
-23.9024143218994,
-30.0049667358398,
37.1030197143555,
41.2666511535645,
-3.96679186820984,
-14.7679138183594,
-12.3199367523193,
26.6830120086670,
28.6641731262207,
6.16778707504273,
-53.1585845947266,
4.68997383117676,
10.7507467269897,
-66.3530883789063,
-13.8652191162109,
33.6226615905762,
20.2462482452393,
8.02377128601074,
55.3839492797852,
-6.49423789978027,
-38.0157165527344,
56.7978096008301,
11.5355806350708,
8.73983001708984,
31.8294296264648,
-53.2135353088379,
18.9280548095703,
48.1781616210938,
-61.1871032714844,
12.1138887405396,
36.5568771362305,
-2.25415539741516,
-22.7559261322022,
-50.0366249084473,
-16.2789115905762,
-34.7165374755859,
-35.2057838439941,
21.2557353973389,
1.33447122573853,
-60.8290214538574,
28.8983783721924,
-23.5847702026367,
-71.3672180175781,
85.5951843261719,
18.2977828979492,
10.7055416107178,
-18.5772590637207,
-3.09329223632813,
43.6553001403809,
-61.3128242492676,
68.0710067749023,
36.3282394409180,
-51.5249252319336,
5.68952274322510,
4.57800197601318,
-42.9737663269043,
-21.5165176391602,
19.8115081787109,
35.0824813842773,
33.8718757629395,
5.58738613128662,
38.6587829589844,
-31.3279018402100,
27.1094017028809,
7.03605890274048,
-31.6186885833740,
42.9520874023438,
25.7433052062988,
57.7511329650879,
-11.2148962020874,
-2.16235256195068,
72.6293182373047,
22.4003543853760,
-30.7711601257324,
24.8457622528076,
-20.2350082397461,
-39.9819869995117,
64.7493667602539,
-32.5978813171387,
-34.7058906555176,
-24.7767944335938,
-9.57128429412842,
46.6326408386231,
-18.3886260986328,
5.64688396453857,
-41.8353691101074,
13.4878997802734,
18.0417175292969,
10.2957210540771,
69.7742614746094,
-65.2382431030273,
48.6511726379395,
41.0595321655273,
-3.84959769248962,
26.6603813171387,
-56.5036621093750,
39.4025192260742,
-24.9393692016602,
16.8276844024658,
38.8875846862793,
-78.0092773437500,
-23.6270198822022,
25.8200225830078,
34.0142173767090,
-73.2981948852539,
-38.7098541259766,
-14.2440900802612,
-42.2492332458496,
20.1064834594727,
9.12325668334961,
-11.9975767135620,
-1.07645046710968,
74.5634841918945,
-10.3673982620239,
-39.1240882873535,
42.1351890563965,
-6.49497032165527,
-15.4909896850586,
-21.3782615661621,
21.7507057189941,
46.4245071411133,
18.3584384918213,
-26.1086139678955,
11.5551443099976,
9.33989334106445,
-56.6083221435547,
75.0902938842773,
33.2356147766113,
-25.3643150329590,
22.5087451934814,
-24.8982009887695,
25.2631206512451,
12.0041742324829,
-75.4632949829102,
6.20219612121582,
-2.65899133682251,
-55.8205032348633,
56.5637435913086,
-2.58828401565552,
-1.36293375492096,
-12.0456781387329,
-63.2559356689453,
37.5852661132813,
-36.3308982849121,
27.8405570983887,
5.04931974411011,
-46.3842430114746,
38.8850021362305,
-38.4843025207520,
46.4255638122559,
40.3407363891602,
-13.4648942947388,
0.800641119480133,
22.8562393188477,
46.9403076171875,
2.47047758102417,
38.3638877868652,
10.4629335403442,
-44.2806320190430,
11.4019403457642,
32.6211318969727,
-64.1767501831055,
-9.76977443695068,
-14.6239356994629,
-80.2506713867188,
6.69973230361939,
7.61401748657227,
-31.3731307983398,
18.2535514831543,
35.8319091796875,
-67.3216323852539,
-19.2715530395508,
50.1722717285156,
6.34368658065796,
27.9968204498291,
64.4382095336914,
8.95486259460449,
-22.0293617248535,
100.572845458984,
11.1373996734619,
-34.6561088562012,
52.4573593139648,
-48.4725418090820,
-17.4496974945068,
4.60370492935181,
-9.47225666046143,
12.0026102066040,
-15.1642923355103,
1.31969070434570,
56.2806358337402,
-4.56334877014160,
-26.2022476196289,
71.5632781982422,
-64.4417800903320,
-27.7465782165527,
83.9777679443359,
14.9396905899048,
-18.9316196441650,
-40.1088752746582,
-32.2631225585938,
-16.3091278076172,
76.7480773925781,
2.11790132522583,
-57.2168006896973,
47.3679618835449,
35.2687873840332,
-12.3578319549561,
-11.7859125137329,
49.8608589172363,
-21.3814563751221,
-17.9341926574707,
53.0495758056641,
-52.6736831665039,
30.0437850952148,
40.7717475891113,
-57.4010658264160,
-35.1962585449219,
-22.5976715087891,
38.0424957275391,
13.2482776641846,
36.9541931152344,
28.2888145446777,
-11.9979982376099,
51.2181358337402,
-33.0463600158691,
-10.7103939056396,
-0.894707739353180,
-59.6361885070801,
7.95266294479370,
-34.5565795898438,
-46.8966026306152,
19.0636329650879,
32.7401123046875,
-2.45088005065918,
10.5618505477905,
-3.26857137680054,
-49.5032463073731,
-18.3708744049072,
39.8896179199219,
20.1789836883545,
-68.1619033813477,
23.2530555725098,
2.73275303840637,
5.39656686782837,
51.9263114929199,
-31.6528739929199,
28.7923030853272,
-8.47624015808106,
17.5382099151611,
45.4528617858887,
-13.3458528518677,
-29.1897354125977,
1.35151529312134,
14.2223768234253,
-36.8479804992676,
23.3980884552002,
-53.5244483947754,
-37.7540855407715,
54.5738639831543,
-17.1847248077393,
44.9828872680664,
9.52105426788330,
-49.9488105773926,
17.5789794921875,
-45.0303688049316,
-16.1904640197754,
0.474797874689102,
4.60163688659668,
49.5089950561523,
33.9187660217285,
53.5088958740234,
-22.9917774200439,
-20.0190544128418,
-33.0185737609863,
16.4903316497803,
33.0548667907715,
6.73020076751709,
53.8879356384277,
-22.0065116882324,
9.01470756530762,
0.546408891677856,
-38.6601409912109,
9.00841808319092,
-5.59678983688355,
-73.9043350219727,
38.4999771118164,
7.04108047485352,
-38.9116439819336,
24.5194492340088,
-56.4915428161621,
3.53865337371826,
-26.2746124267578,
3.92729783058167,
47.5369567871094,
29.7076473236084,
26.3320369720459,
7.26682329177856,
54.4688796997070,
22.0013103485107,
32.7580070495606,
42.3009490966797,
-6.55741024017334,
-42.5459327697754,
-13.3195066452026,
-12.4920387268066,
-41.9214591979981,
-39.6148681640625,
-29.5049686431885,
-5.94527769088745,
-15.9488649368286,
-52.8075866699219,
-3.61644244194031,
4.65624427795410,
1.70652735233307,
52.3782882690430,
-13.6542434692383,
35.1435585021973,
20.2065181732178,
19.9260005950928,
53.3873634338379,
-3.55785131454468,
30.1035442352295,
46.3420486450195,
-13.4113054275513,
-32.9855880737305,
70.1295394897461,
5.98101139068604,
-3.49472951889038,
12.5718441009521,
10.5529975891113,
18.8527812957764,
-28.5757846832275,
-7.56277942657471,
-41.6028137207031,
14.1959533691406,
-34.2911758422852,
-57.2343559265137,
-0.796233415603638,
-17.9099082946777,
36.5602035522461,
-9.71606731414795,
-33.3843040466309,
69.3317184448242,
-8.85242652893066,
-43.8089675903320,
54.4730911254883,
-45.6184768676758,
-9.55883979797363,
57.7298431396484,
-14.7509241104126,
33.4353179931641,
9.44063377380371,
-28.7915325164795,
14.8077125549316,
22.8228626251221,
-17.9796581268311,
-37.3453254699707,
48.5178871154785,
14.8367919921875,
-38.9339904785156,
17.2635669708252,
14.4973831176758,
-3.51628541946411,
-19.6861820220947,
46.7425842285156,
39.3533897399902,
35.4766120910645,
15.7811880111694,
-42.4361000061035,
29.1029758453369,
-22.5361843109131,
13.6698875427246,
36.4399909973145,
26.8295230865479,
8.63103580474854,
-18.9839782714844,
14.7608566284180,
-21.6106662750244,
37.5852088928223,
-20.8578987121582,
-40.9388771057129,
33.4858131408691,
15.4059057235718,
-43.7124748229981,
-2.28433918952942,
41.0581092834473,
-12.4021654129028,
-6.38958168029785,
39.1591644287109,
17.4146385192871,
-50.0528869628906,
38.2527923583984,
5.18085813522339,
-23.2924728393555,
-15.4862613677979,
-24.1688499450684,
37.7812271118164,
12.0746879577637,
14.2080831527710,
-41.5220909118652,
31.5226612091064,
15.8989477157593,
-55.9686584472656,
26.7581138610840,
-39.1703186035156,
18.5872936248779,
20.1445980072022,
-49.9872055053711,
-0.394193083047867,
24.4242401123047,
-9.77887535095215,
-48.3950843811035,
-32.1757392883301,
-2.19093418121338,
6.53294658660889,
-66.9795837402344,
53.9520874023438,
1.19041776657105,
-31.6954441070557,
50.6379165649414,
-68.1844100952148,
7.63305282592773,
43.2498550415039,
-17.1052932739258,
-51.1386146545410,
50.7337913513184,
11.9357137680054,
-33.4330825805664,
5.71447753906250,
6.07217311859131,
29.8185672760010,
-33.6229438781738,
45.1868019104004,
-15.6563310623169,
-36.1909751892090,
18.3628005981445,
16.1875228881836,
39.3396835327148,
17.8168544769287,
18.5976505279541,
-53.7112808227539,
-19.8416328430176,
-10.2971925735474,
-13.9922428131104,
55.8911743164063,
27.1762332916260,
36.6184387207031,
7.15268945693970,
-6.40040731430054,
19.7359867095947,
-28.2066307067871,
-28.5272045135498,
-12.7424545288086,
-0.257941335439682,
-13.9939002990723,
-0.758831799030304,
49.5601158142090,
-5.97515726089478,
3.87996912002563,
58.3558197021484,
11.8413467407227,
-20.5965633392334,
-48.2604751586914,
3.57008790969849,
34.8635330200195,
-51.9655609130859,
35.7022819519043,
63.4015541076660,
-49.1675148010254,
38.4671287536621,
70.1178283691406,
-19.5777873992920,
-17.6210842132568,
3.84144473075867,
44.2181777954102,
40.4880027770996,
-52.9839401245117,
-24.2238273620605,
33.4645576477051,
-38.9644699096680,
-50.2559852600098,
-12.8533763885498,
-32.8947525024414,
-55.4139633178711,
-30.2197723388672,
-15.5547819137573,
-11.9441432952881,
11.5520267486572,
-21.5887088775635,
6.22249031066895,
-34.2732048034668,
-55.6620178222656,
65.7560348510742,
-9.93038940429688,
12.7296123504639,
11.6481847763062,
-18.2316684722900,
39.9033546447754,
-43.4891929626465,
1.85967838764191,
19.8637065887451,
-4.17075443267822,
-33.6368522644043,
13.5511131286621,
28.7742671966553,
-27.6036510467529,
28.8739089965820,
13.3561239242554,
48.7162513732910,
25.7813301086426,
-8.92962646484375,
24.4692249298096,
43.1832160949707,
56.9098320007324,
2.69010210037231,
5.52678012847900,
22.5355167388916,
-13.6779375076294,
-8.91315841674805,
30.6995582580566,
-13.5851211547852,
-60.1051330566406,
-7.00819349288940,
-20.1082401275635,
-37.6439323425293,
0.435294419527054,
24.3401641845703,
40.7272338867188,
23.8708152770996,
10.6065568923950,
-30.0709056854248,
7.99261856079102,
-11.3226652145386,
-47.7675094604492,
30.4035758972168,
20.5722866058350,
39.1741485595703,
32.3233222961426,
37.4554901123047,
10.8289613723755,
22.8675861358643,
16.5590362548828,
-43.0730781555176,
41.4778022766113,
0.758259892463684,
-1.61338996887207,
44.7878913879395,
48.5422706604004,
-30.3899230957031,
-16.8823490142822,
12.8710098266602,
-38.1455993652344,
60.3702430725098,
0.589805960655212,
2.86515092849731,
-23.3744239807129,
-37.5025138854981,
3.59428834915161,
-28.3988342285156,
69.4674377441406,
-38.5134544372559,
-18.0577774047852,
50.9940643310547,
-42.6490478515625,
64.9125289916992,
34.4206962585449,
-23.6332302093506,
16.0259246826172,
7.88730573654175,
38.2431831359863,
32.9348449707031,
1.70412802696228,
23.7071094512939,
42.3110809326172,
27.1528453826904,
28.5834426879883,
-5.16251182556152,
28.7841949462891,
31.2215862274170,
-50.6304702758789,
-26.2419033050537,
30.2594032287598,
14.9319934844971,
0.748410344123840,
11.8811454772949,
-61.9522171020508,
-28.7130451202393,
58.3588562011719,
38.1415481567383,
37.2712631225586,
-22.8537235260010,
-50.7760353088379,
21.6719913482666,
53.5736923217773,
21.3508567810059,
-35.2750854492188,
-14.9516401290894,
40.2975349426270,
24.7105636596680,
-16.7083911895752,
60.6900062561035,
53.3868751525879,
-62.7163505554199,
38.3630409240723,
56.9617004394531,
-43.1207122802734,
-20.6663246154785,
-17.2029113769531,
22.1877899169922,
29.9427032470703,
-38.3299674987793,
-25.9656753540039,
7.77024078369141,
-37.8271064758301,
-31.4777908325195,
55.4357872009277,
-18.4833145141602,
-14.2747945785522,
61.9466361999512,
26.5338001251221,
18.6922721862793,
26.5397377014160,
17.6005611419678,
-29.4410247802734,
22.1887302398682,
-4.42572355270386,
8.53335475921631,
32.0422782897949,
-35.1988372802734,
69.8407669067383,
18.3456344604492,
-54.0079307556152,
25.7569847106934,
48.1200447082520,
-10.0661745071411,
10.8301897048950,
61.1848678588867,
-10.7385425567627,
60.0754661560059,
17.0862770080566,
-15.2464981079102,
29.1898441314697,
-37.7255935668945,
45.2573471069336,
5.49331569671631,
-48.3992156982422,
11.8959646224976,
34.5515747070313,
-19.9653015136719,
23.8703556060791,
34.0890998840332,
-26.1627178192139,
46.0228500366211,
18.4762401580811,
38.1881599426270,
-4.68968009948731,
-5.31003427505493,
31.1854782104492,
-31.8709774017334,
1.80613923072815,
9.84785175323486,
21.4847393035889,
-3.56278157234192,
-10.6422300338745,
48.1542282104492,
31.5279655456543,
-10.6464309692383,
-16.2717533111572,
-9.55655574798584,
23.2314720153809,
17.1207942962647,
9.49153709411621,
68.8637542724609,
18.3528213500977,
-43.8865699768066,
-7.48158836364746,
45.6029357910156,
49.4522094726563,
13.3032169342041,
0.115310072898865,
-34.2246398925781,
16.8860359191895,
5.38293218612671,
-27.1131458282471,
47.8439254760742,
43.4717102050781,
11.5827646255493,
-36.1417999267578,
4.19307708740234,
26.6641178131104,
-24.8301143646240,
30.4208641052246,
26.4531631469727,
5.94827651977539,
49.6804466247559,
10.0229597091675,
-43.4065704345703,
60.9001693725586,
35.3140144348145,
-60.8713531494141,
36.0761070251465,
2.72263526916504,
1.56395995616913,
7.55288743972778,
-19.4912910461426,
15.3177862167358,
-35.5219154357910,
-4.69674634933472,
54.4998359680176,
36.0637207031250,
-51.2627334594727,
-44.9527397155762,
33.6136054992676,
34.8751525878906,
-32.9073829650879,
-13.5235233306885,
36.9821548461914,
-38.7030906677246,
14.0864915847778,
55.8142089843750,
-8.74973678588867,
17.3948040008545,
25.7049732208252,
23.6037483215332,
46.6007614135742,
7.03555393218994,
14.0450925827026,
64.6031799316406,
5.10544013977051,
-23.7271747589111,
74.9521560668945,
5.82297849655151,
-46.4624099731445,
67.0680084228516,
-23.4617271423340,
-37.9899787902832,
47.9099197387695,
50.0489311218262,
10.3171787261963,
-47.8049736022949,
-24.5287475585938,
-9.43583011627197,
38.7970466613770,
-23.0632152557373,
-52.1537322998047,
50.4689712524414,
1.48521745204926,
-38.9797210693359,
26.8120574951172,
-4.35648965835571,
-29.0737018585205,
26.3238506317139,
18.6879806518555,
18.4965171813965,
-33.8372535705566,
-20.0715389251709,
33.1462516784668,
0.302526146173477,
24.4837303161621,
39.9309997558594,
12.5895509719849,
-15.7476024627686,
9.59563732147217,
4.73912906646729,
41.3208656311035,
58.7326507568359,
-6.15525054931641,
49.5866508483887,
24.9373874664307,
5.18294000625610,
-23.6766376495361,
-14.0280408859253,
50.0900001525879,
-14.7392301559448,
31.9160976409912,
-23.2714824676514,
-6.67581939697266,
50.7425575256348,
-28.6131114959717,
12.5074558258057,
35.3765907287598,
59.1793365478516,
-21.1466312408447,
-31.8172245025635,
12.2899456024170,
-25.3591041564941,
16.6879940032959,
-29.2554492950439,
-31.3655052185059,
22.9406490325928,
12.0027456283569,
-35.5096054077148,
-47.4510116577148,
-12.2088327407837,
19.8594017028809,
4.30841016769409,
-7.50652313232422,
58.8809852600098,
5.93805646896362,
-10.8046522140503,
-20.5362567901611,
14.4920501708984,
78.6649398803711,
-18.5258712768555,
-7.52860498428345,
19.9458446502686,
-1.84639668464661,
24.1872348785400,
8.40562438964844,
-26.8371372222900,
39.0913124084473,
16.8748703002930,
-38.1490020751953,
-5.48626518249512,
-53.7594871520996,
-18.9679908752441,
-25.5688533782959,
-24.9921131134033,
44.0236511230469,
-10.0830354690552,
-3.38761854171753,
1.09301459789276,
15.2667131423950,
-12.2068099975586,
-49.9666557312012,
9.20098972320557,
17.8215389251709,
23.7266292572022,
-44.4799156188965,
11.3203954696655,
43.3892478942871,
-51.0005874633789,
16.8056354522705,
10.5281524658203,
25.9497814178467,
1.36318135261536,
-34.9670295715332,
48.2642211914063,
-56.4065704345703,
-24.3993625640869,
32.7820854187012,
-52.8781166076660,
-11.7037677764893,
-10.9637889862061,
12.3153419494629,
39.8207740783691,
40.1001243591309,
-21.9474620819092,
-24.6038074493408,
7.19004344940186,
-38.8383522033691,
26.1295204162598,
-36.7621994018555,
-56.4289855957031,
43.2038955688477,
31.3180217742920,
-3.84739685058594,
3.20573449134827,
39.1757774353027,
38.3289031982422,
1.28264069557190,
-28.9014949798584,
-12.8684139251709,
23.7617683410645,
-6.30763673782349,
-47.0791130065918,
42.9196166992188,
19.4998950958252,
-21.6451148986816,
-3.31494021415710,
-21.5681743621826,
-12.1310586929321,
-43.2396430969238,
-2.81734085083008,
-35.1215553283691,
-20.4952888488770,
44.1237144470215,
-14.3361129760742,
14.3184499740601,
23.8292961120605,
-16.7768440246582,
-10.2458181381226,
-4.34635114669800,
-21.4763774871826,
-20.2776165008545,
1.39926624298096,
-37.7630691528320,
-23.5692234039307,
38.7739524841309,
25.1237030029297,
-2.08842849731445,
-54.7700042724609,
20.3437881469727,
19.4352149963379,
-52.1078529357910,
62.2663383483887,
6.54956579208374,
-59.4567565917969,
7.02766561508179,
9.69390964508057,
-29.1305561065674,
-26.3529338836670,
-5.82154846191406,
-24.8342247009277,
28.0069103240967,
12.4618577957153,
-35.5886573791504,
-11.3770809173584,
-23.4959907531738,
-20.8649139404297,
-20.3425559997559,
-37.8787918090820,
-28.3344440460205,
-6.37633657455444,
-17.7989788055420,
-9.35177326202393,
-2.64448523521423,
-22.7545299530029,
-12.3372077941895,
-30.6830196380615,
-7.57718229293823,
1.45293653011322,
-29.2139568328857,
-33.9445877075195,
-33.0373420715332,
35.1098518371582,
-16.8670387268066,
-53.6207656860352,
46.1243400573731,
16.2706451416016,
-5.16729593276978,
14.0088777542114,
-27.7269172668457,
-21.7340545654297,
-1.47214102745056,
-58.5607910156250,
-23.5069942474365,
37.3163833618164,
17.0281028747559,
15.3918590545654,
-18.1778526306152,
4.73547267913818,
-9.72891998291016,
-32.6923027038574,
-7.25730705261231,
3.13127899169922,
-20.2553253173828,
-56.1004028320313,
-13.7254209518433,
14.3332281112671,
27.3534774780273,
22.1461963653564,
45.2539939880371,
-6.26394224166870,
-30.5163688659668,
1.26698708534241,
-31.5513057708740,
6.19447612762451,
42.2779808044434,
4.76911640167236,
-2.68792843818665,
58.5035972595215,
-32.4721984863281,
-23.3346366882324,
48.5893096923828,
-1.75134110450745,
13.0017910003662,
-8.70049667358398,
-29.5541496276855,
-15.1209840774536,
-10.0634632110596,
-29.7107486724854,
6.50338697433472,
44.1653327941895,
-39.4755401611328,
-27.7967720031738,
65.0276947021484,
-9.14956951141357,
-40.0154876708984,
55.3112220764160,
-30.0012435913086,
-36.7765426635742,
49.5013809204102,
3.07809281349182,
25.7126274108887,
-15.4364805221558,
-30.3333015441895,
20.6055812835693,
25.6635608673096,
18.7083549499512,
-9.87398433685303,
29.4959754943848,
8.77398395538330,
6.48356914520264,
17.2783222198486,
36.8438529968262,
45.2652549743652,
-37.3277854919434,
24.3058414459229,
9.16310501098633,
-51.4048728942871,
-23.1328620910645,
-18.8957347869873,
-22.9529705047607,
-0.358069270849228,
20.6977996826172,
4.32809257507324,
33.0529937744141,
-19.5938682556152,
20.4099769592285,
8.98251152038574,
-4.65621185302734,
22.9196281433105,
-44.8309288024902,
40.9892272949219,
8.60838890075684,
15.5862035751343,
57.1406097412109,
-8.67877388000488,
-30.0970993041992,
-32.2707405090332,
11.8405427932739,
22.8543815612793,
18.5322437286377,
-8.14905834197998,
-28.0896224975586,
21.2416687011719,
28.1583614349365,
36.5862846374512,
32.6542015075684,
-22.7649078369141,
-21.8330993652344,
-4.44428443908691,
62.4469680786133,
-5.04630470275879,
-16.7823333740234,
52.0977783203125,
-50.7998809814453,
-26.6385269165039,
-18.6123142242432,
-22.0216102600098,
2.30667257308960,
-43.1409797668457,
-42.1423912048340,
-7.78857898712158,
-31.9247684478760,
-34.8152732849121,
11.3279104232788,
-17.0527763366699,
7.69992113113403,
1.57694637775421,
7.55149078369141,
27.5784378051758,
16.5508594512939,
19.4547557830811,
-37.9385414123535,
0.172097966074944,
-6.48848867416382,
-34.5817680358887,
5.34419250488281,
-46.4923362731934,
25.7622127532959,
49.0465507507324,
-45.1336250305176,
46.8760833740234,
0.774808883666992,
-54.4254684448242,
-11.6420650482178,
-36.4853668212891,
15.1847705841064,
-29.8279953002930,
23.2537612915039,
56.7088775634766,
-36.1324424743652,
13.6101789474487,
-23.3122558593750,
-17.8673610687256,
27.5751419067383,
-2.10712075233459,
9.56053924560547,
3.66970968246460,
-22.9728775024414,
-8.06701087951660,
32.8180084228516,
11.9559211730957,
25.0465507507324,
4.14509439468384,
21.5443954467773,
45.9305305480957,
-37.0987396240234,
-16.5753688812256,
44.2082977294922,
17.6563968658447,
-3.30337166786194,
45.5233726501465,
-3.67483997344971,
-1.09573805332184,
46.8792572021484,
14.2145824432373,
7.25457668304443,
10.0578289031982,
-7.70980167388916,
-24.8716907501221,
1.39351892471313,
12.2543716430664,
31.9589042663574,
22.3997325897217,
44.4086341857910,
-1.98539769649506,
-49.2928085327148,
59.2892456054688,
-6.06667804718018,
-35.0290451049805,
63.1961898803711,
20.8067436218262,
-39.8974876403809,
-13.5705671310425,
9.17763042449951,
-12.4787349700928,
-5.40087604522705,
-11.1470775604248,
39.4486351013184,
18.6176052093506,
7.17428350448608,
16.8511009216309,
-36.2173767089844,
42.6246757507324,
-35.2033882141113,
-8.10208225250244,
56.4946060180664,
-39.5239639282227,
-1.97241306304932,
17.4108600616455,
24.9081287384033,
-26.8878536224365,
23.2881031036377,
28.0652561187744,
-55.0891647338867,
12.2444849014282,
-22.6768074035645,
10.8291845321655,
28.6125335693359,
17.7815399169922,
66.3974151611328,
3.65934109687805,
-37.7142372131348,
2.98813343048096,
14.6336336135864,
-50.4670143127441,
4.51627731323242,
26.5228080749512,
-41.4061546325684,
-41.9559593200684,
-5.44829082489014,
-11.4799737930298,
-4.69091939926148,
20.0996322631836,
-1.74550044536591,
4.55458593368530,
-1.83900725841522,
45.4242248535156,
24.5655403137207,
21.7082881927490,
55.5421295166016,
13.6452589035034,
54.4909133911133,
21.5440979003906,
7.74630117416382,
43.4108314514160,
-23.5752353668213,
32.0314178466797,
52.8281059265137,
-45.2949523925781,
-18.0757560729980,
12.6135320663452,
-3.98355865478516,
4.10988759994507,
44.6585922241211,
21.3917503356934,
-9.58360004425049,
9.28512954711914,
13.5124216079712,
3.08142733573914,
-37.4060745239258,
18.1455268859863,
5.22065639495850,
-47.1632156372070,
50.7050247192383,
14.1224060058594,
-39.6791038513184,
42.1768760681152,
42.9985847473145,
19.1764278411865,
22.8860187530518,
-10.1107540130615,
38.1245727539063,
61.8169250488281,
-13.7149114608765,
-26.9799175262451,
-20.4772605895996,
-9.37142467498779,
-1.58150768280029,
-22.3190994262695,
-31.9031829833984,
-12.8494081497192,
-41.2281837463379,
-51.2116622924805,
44.1902885437012,
1.22403478622437,
-46.5150032043457,
13.7615442276001,
-29.5781288146973,
-16.9996891021729,
23.7574539184570,
2.37514734268188,
8.89303970336914,
22.8151912689209,
-7.76227855682373,
-5.32889890670776,
39.4157485961914,
-9.98790168762207,
7.07763290405273,
-13.5298528671265,
-27.4455032348633,
15.0360603332520,
-23.0132331848145,
-0.956893801689148,
-24.6794548034668,
6.91793251037598,
21.7030982971191,
-34.3249931335449,
-21.0632076263428,
9.18263912200928,
-2.74844074249268,
-1.19712746143341,
35.7286834716797,
31.4570713043213,
-11.0092306137085,
-19.0409717559814,
57.5521316528320,
-7.50090408325195,
11.3175382614136,
34.1026077270508,
-4.04755830764771,
34.2593574523926,
-12.6006975173950,
1.42572605609894,
-20.8535881042480,
35.0469589233398,
10.4757814407349,
-50.0953102111816,
37.1648559570313,
-9.55156803131104,
-14.5932531356812,
16.8604984283447,
35.0663566589356,
28.1725845336914,
-29.6497058868408,
13.6397066116333,
31.8276500701904,
1.05729353427887,
-16.3877086639404,
-26.5977439880371,
40.2334327697754,
1.22689783573151,
-62.2958030700684,
3.45971584320068,
46.0876960754395,
16.5552005767822,
16.8432674407959,
2.29864788055420,
-30.7279796600342,
26.3582992553711,
-15.6602010726929,
-15.5231027603149,
-2.34686923027039,
-57.7021179199219,
-14.3270244598389,
30.6651039123535,
21.7303466796875,
13.9761381149292,
28.5437164306641,
-42.5302543640137,
6.61401081085205,
71.6863327026367,
-17.1821708679199,
-39.1856956481934,
-9.68546867370606,
19.6830730438232,
-6.61495161056519,
-1.82614636421204,
18.9733409881592,
-12.2562818527222,
-43.1544876098633,
-38.8078575134277,
7.37379455566406,
18.2347965240479,
45.7769889831543,
0.301674664020538,
-37.1640396118164,
-10.0540733337402,
1.67646729946136,
3.60369825363159,
-4.13601541519165,
44.3386688232422,
21.7322463989258,
-4.20841312408447,
-14.2016572952271,
34.0169410705566,
10.1816492080688,
-13.7475967407227,
28.4375305175781,
-35.0648040771484,
34.9544219970703,
3.38660979270935,
-27.2126331329346,
-11.8802223205566,
-29.9770202636719,
46.2747573852539,
2.77680087089539,
1.68148767948151,
23.1945972442627,
-23.4961833953857,
-13.2406444549561,
8.95480632781982,
-21.2847213745117,
7.08126640319824,
7.93234825134277,
-49.6518173217773,
23.8752593994141,
-18.6280918121338,
-23.7137088775635,
36.3630561828613,
-66.4750366210938,
-16.7182369232178,
26.6574020385742,
-41.4330482482910,
-20.8120861053467,
-0.721129477024078,
0.977861225605011,
12.4799928665161,
-19.8493499755859,
-46.5657844543457,
-8.19257164001465,
-5.95396041870117,
-49.0103225708008,
27.3336563110352,
37.9920921325684,
-43.1842613220215,
26.7566871643066,
29.6318988800049,
21.8410663604736,
-5.09712314605713,
-33.2762413024902,
29.3867340087891,
-10.8267393112183,
48.2654571533203,
18.0002422332764,
-51.4417839050293,
16.3384151458740,
23.0620841979980,
-8.59460830688477,
-58.1017875671387,
33.9916458129883,
-12.8016939163208,
-45.0821914672852,
15.6584367752075,
-9.26290607452393,
17.7004737854004,
-11.7200918197632,
20.0959930419922,
-23.3512783050537,
-35.1905288696289,
-27.1784133911133,
15.7926311492920,
16.2357673645020,
-18.7228832244873,
37.5918540954590,
-27.2081375122070,
33.5735702514648,
21.4845714569092,
-15.2870082855225,
-16.9266052246094,
-34.2345504760742,
-28.0036220550537,
-16.5301551818848,
17.5547351837158,
-10.2554206848145,
15.3138685226440,
-40.9027595520020,
20.7348041534424,
52.8580589294434,
-21.6667041778564,
15.2484264373779,
15.6195507049561,
54.4484939575195,
-7.01472949981689,
-5.15486621856689,
54.3036499023438,
-17.7432098388672,
-45.9271507263184,
-23.6184730529785,
20.9963703155518,
-0.995890438556671,
10.4610490798950,
-8.38274478912354,
-6.11234998703003,
12.8760309219360,
-75.0194168090820,
20.9354915618897,
34.1980857849121,
-53.1377067565918,
-21.5144958496094,
2.10518598556519,
10.1155815124512,
-31.3765010833740,
29.7242603302002,
42.7263336181641,
2.58425593376160,
34.8080711364746,
-40.8988380432129,
27.1530570983887,
31.0228996276855,
-45.5873603820801,
12.4397745132446,
-18.0133991241455,
-2.26537322998047,
-32.1379280090332,
-13.2929096221924,
5.65052413940430,
-40.0184516906738,
-36.7351684570313,
-29.1222476959229,
12.8411512374878,
-37.6578559875488,
-24.1354808807373,
28.9119586944580,
34.6614379882813,
-26.9844303131104,
-2.00739622116089,
60.9548912048340,
-0.813469707965851,
-6.49128293991089,
-23.0128078460693,
-7.79549360275269,
47.0802650451660,
23.0181846618652,
-40.7940750122070,
6.23124694824219,
17.9617595672607,
-42.8864288330078,
-20.9695758819580,
24.2689094543457,
23.3986549377441,
-5.48257398605347,
-37.8963470458984,
-7.62202262878418,
50.7977676391602,
-8.61952400207520,
7.55708456039429,
1.43366658687592,
-27.1688270568848,
-17.9836616516113,
-31.7751903533936,
46.8779220581055,
10.8431463241577,
-18.5403327941895,
10.2108783721924,
16.0589237213135,
40.7023925781250,
0.452456235885620,
29.5532798767090,
-5.92858695983887,
-36.4678955078125,
35.5076217651367,
-18.9568386077881,
-8.97403526306152,
-6.83744525909424,
-43.2007293701172,
-6.33036994934082,
6.37434196472168,
35.8781814575195,
2.58174300193787,
17.8904476165772,
45.6699905395508,
17.7699947357178,
42.9499969482422,
37.6535797119141,
-28.5062751770020,
-1.07284128665924,
42.0978507995606,
-20.1477909088135,
8.97522163391113,
-22.6726188659668,
-2.77356314659119,
43.8374938964844,
-6.02242326736450,
-12.5075645446777,
-19.1257324218750,
24.4098606109619,
-8.18019580841065,
32.8814392089844,
43.1947174072266,
-8.08916759490967,
29.7441673278809,
-5.36643218994141,
29.1644725799561,
9.27036857604981,
-4.64161062240601,
41.6718597412109,
-26.4469909667969,
-33.7164649963379,
-7.31031799316406,
23.9064292907715,
-29.8112030029297,
-55.0621070861816,
26.2071952819824,
-36.6189651489258,
-15.5108852386475,
48.3632583618164,
-11.0625047683716,
19.2912063598633,
9.25288105010986,
-17.2914924621582,
-13.9175529479980,
-11.2025833129883,
44.7656745910645,
-30.3925209045410,
7.98960494995117,
18.7878513336182,
-40.5683250427246,
3.63986706733704,
-32.7457733154297,
-2.45402717590332,
25.9458713531494,
14.1191463470459,
-8.38275432586670,
-6.57265377044678,
-18.0797061920166,
25.2781505584717,
7.93627548217773,
-49.3482780456543,
-2.59662175178528,
-34.4325637817383,
16.7486343383789,
-21.9054718017578,
-20.1887397766113,
46.6272354125977,
-36.3877220153809,
-1.64235389232636,
22.2439384460449,
13.0181713104248,
22.0756015777588,
-24.9024791717529,
7.68303871154785,
47.1038627624512,
-15.7970838546753,
-2.07666897773743,
-8.98120117187500,
-26.0166110992432,
53.7414932250977,
-14.1436862945557,
-20.2867431640625,
32.1473007202148,
-19.6377124786377,
-3.44643330574036,
-7.65592288970947,
-24.8423500061035,
-25.7643928527832,
-27.5670089721680,
-36.4176445007324,
-25.9235191345215,
-30.8216533660889,
-14.7190103530884,
12.9192819595337,
-20.0884304046631,
-30.9833774566650,
-17.7482242584229,
28.9965114593506,
18.1124229431152,
7.30819082260132,
9.05364227294922,
-10.4946737289429,
10.7744588851929,
52.5533027648926,
3.81494045257568,
0.432887375354767,
43.6631050109863,
-32.8672027587891,
-4.03007555007935,
-14.3737630844116,
10.2223205566406,
37.8605194091797,
-31.3814964294434,
19.7184028625488,
18.2777175903320,
-28.5289001464844,
-18.3180751800537,
-7.78744649887085,
7.14260196685791,
24.5807418823242,
-24.6508369445801,
-18.2678813934326,
9.56804084777832,
-15.3940973281860,
-20.9943618774414,
4.16542720794678,
24.6411094665527,
-37.9873542785645,
-18.9202175140381,
9.23921775817871,
-10.8959369659424,
22.5698032379150,
-27.0437717437744,
-37.1855773925781,
2.93060827255249,
-19.4032478332520,
12.1754512786865,
-1.76821827888489,
-21.7618694305420,
8.53138542175293,
6.95765161514282,
26.6797008514404,
13.7932138442993,
-6.94843626022339,
10.8300457000732,
18.3330001831055,
-25.1188602447510,
0.941851556301117,
57.4180107116699,
-17.8133220672607,
-17.9716300964355,
22.3310699462891,
-22.3531494140625,
-5.05639076232910,
28.5740814208984,
-0.0385491512715817,
0.239660620689392,
46.9354400634766,
-12.5912475585938,
-30.8055362701416,
36.6208877563477,
15.5779170989990,
-12.9046220779419,
3.08149790763855,
35.0461158752441,
26.2131919860840,
35.5258674621582,
27.5726013183594,
38.7222290039063,
19.9222030639648,
-23.5376148223877,
-3.20420122146606,
-2.36059808731079,
43.3360061645508,
10.8552417755127,
3.59321737289429,
7.57251882553101,
-27.9330558776855,
10.9255876541138,
-16.8872413635254,
19.7681236267090,
4.75287771224976,
-21.0607643127441,
53.6281356811523,
31.1773128509522,
-9.36104488372803,
-26.6192893981934,
23.2889404296875,
17.4296989440918,
19.9922275543213,
41.8036613464356,
13.1787080764771,
39.5649070739746,
19.7847194671631,
-19.6488456726074,
-16.6612854003906,
34.2937011718750,
-5.08141660690308,
-41.5807151794434,
21.9303226470947,
26.6707210540772,
-7.57835102081299,
-10.6920833587646,
0.653505504131317,
-33.4389915466309,
-3.37352538108826,
26.8477725982666,
-35.0578041076660,
-36.5274124145508,
37.9431266784668,
7.25494527816773,
-50.2607002258301,
10.3677892684937,
-14.7389478683472,
9.12152290344238,
9.03133392333984,
-17.7408199310303,
-3.05672073364258,
-29.5576496124268,
44.0851783752441,
11.1938343048096,
15.5273590087891,
21.3172149658203,
12.5891742706299,
0.0549328587949276,
-27.4950351715088,
-0.253694713115692,
-27.5650062561035,
31.3328895568848,
22.8166103363037,
-11.5004024505615,
-27.1956424713135,
-4.95970010757446,
-28.8901844024658,
-3.39086532592773,
30.7533092498779,
-37.3169059753418,
49.5680656433106,
5.42428636550903,
10.2736558914185,
48.1009635925293,
3.43527984619141,
43.6805000305176,
2.75487828254700,
32.0551719665527,
52.9089164733887,
20.5553703308105,
31.2199192047119,
16.8205394744873,
-15.5686626434326,
-17.5912570953369,
-7.04707670211792,
-36.9272003173828,
14.9018888473511,
-14.2897148132324,
-59.2141113281250,
3.77308869361877,
-11.9242095947266,
-10.6947154998779,
-16.5226650238037,
37.4798469543457,
24.7709636688232,
-50.3503227233887,
23.6398792266846,
14.5024881362915,
7.89380264282227,
21.4842891693115,
31.1736068725586,
29.2936248779297,
6.30447959899902,
23.6496505737305,
12.6771097183228,
45.0002059936523,
17.5190086364746,
-16.6570339202881,
12.1536912918091,
12.8603076934814,
-31.0787677764893,
-9.38326358795166,
48.8886413574219,
-22.9420108795166,
-27.4966945648193,
5.89750289916992,
-20.1671867370605,
17.6325473785400,
18.6514625549316,
-37.4997367858887,
-7.98517847061157,
18.5401248931885,
-7.88084936141968,
7.36005544662476,
-16.9036464691162,
-23.5142402648926,
26.8775806427002,
24.7076797485352,
24.8844661712647,
-15.7615375518799,
-39.1614036560059,
10.4723138809204,
34.9039573669434,
14.5607624053955,
-4.09095382690430,
17.1873512268066,
13.0296745300293,
12.8983249664307,
29.7927398681641,
41.4859848022461,
8.10179710388184,
15.6265020370483,
40.7175369262695,
-19.4406528472900,
6.29751920700073,
38.8868598937988,
11.1036100387573,
-60.3119239807129,
-1.57452607154846,
33.7457427978516,
-41.6864776611328,
36.2452583312988,
-5.06177520751953,
9.07662296295166,
33.4433441162109,
7.18511581420898,
49.0618400573731,
9.44254970550537,
-30.9381122589111,
3.71299672126770,
31.0653228759766,
-39.6202621459961,
30.1970558166504,
36.6228942871094,
-15.6003360748291,
13.7100877761841,
48.5010566711426,
-5.09098196029663,
-25.3091335296631,
12.0473003387451,
-26.8303966522217,
38.5272140502930,
-37.9374465942383,
-24.4276256561279,
31.6435985565186,
-44.6683959960938,
-6.38145494461060,
4.84069871902466,
9.46351337432861,
2.99132418632507,
-25.5410137176514,
10.2749223709106,
-0.726517796516419,
-10.7424640655518,
29.4496078491211,
27.1249294281006,
36.3389434814453,
11.5914831161499,
11.3251523971558,
-36.9916992187500,
8.77327251434326,
36.6447105407715,
-41.4632110595703,
16.0618457794189,
1.05391895771027,
25.5081405639648,
-15.4987907409668,
-13.6585378646851,
12.1773748397827,
-33.6977081298828,
-8.15436935424805,
-29.2634544372559,
59.3474922180176,
11.4253597259521,
-36.7619056701660,
27.9107952117920,
-14.0341005325317,
-12.4385519027710,
-30.3638458251953,
-11.0452241897583,
-6.27556991577148,
-10.2923393249512,
37.9282684326172,
-7.41422176361084,
37.3851661682129,
31.0194263458252,
-29.8212242126465,
40.6010627746582,
16.5985908508301,
-7.93067789077759,
-25.8547935485840,
-3.92810630798340,
35.1041564941406,
22.7168254852295,
20.3704948425293,
-39.9520416259766,
-10.2832698822021,
20.9994983673096,
-11.0614395141602,
-21.8817443847656,
-27.5892009735107,
-26.5626277923584,
-16.5889968872070,
36.8560600280762,
-3.99888396263123,
-32.3639793395996,
30.6166229248047,
-12.8083534240723,
10.2726812362671,
42.0604667663574,
-31.4736061096191,
8.64343833923340,
50.1120910644531,
4.23445034027100,
-13.4781999588013,
9.33269500732422,
42.0245208740234,
1.25601875782013,
15.6158857345581,
49.9145889282227,
-12.6748342514038,
-15.3248805999756,
-22.6563720703125,
-2.11333632469177,
-8.86059093475342,
-15.9177322387695,
3.54069256782532,
17.3928833007813,
9.62762069702148,
-34.7257995605469,
14.4756078720093,
5.15458917617798,
28.1956386566162,
-14.8272457122803,
-23.1629505157471,
31.9270248413086,
-39.4970054626465,
21.1219997406006,
33.0416336059570,
8.66677188873291,
9.31205940246582,
-4.91172170639038,
37.3093490600586,
36.3727798461914,
12.0394334793091,
-27.1859111785889,
-12.9419956207275,
-13.3512210845947,
-29.2756443023682,
-9.71936893463135,
33.3306121826172,
21.8707809448242,
-36.6062164306641,
35.5551071166992,
-0.142304539680481,
-30.2486610412598,
45.6633148193359,
8.23095893859863,
-38.8760948181152,
31.6374301910400,
27.3466720581055,
-0.800831556320190,
30.0582942962647,
-6.18576622009277,
23.7319393157959,
-11.6646394729614,
8.43601417541504,
49.3648414611816,
28.5196361541748,
-9.05348587036133,
-12.3015995025635,
45.5609817504883,
-43.4187088012695,
-12.5955238342285,
22.4257259368897,
-4.66416406631470,
13.2919731140137,
-15.2841596603394,
-3.80575895309448,
16.3395748138428,
-12.4530858993530,
-31.5315837860107,
2.32243728637695,
-30.4445533752441,
1.50946187973022,
36.6197509765625,
1.58185470104218,
30.5307979583740,
-17.3023586273193,
-24.4514484405518,
12.6694383621216,
-10.9881410598755,
-31.7931919097900,
-15.2145242691040,
37.3057174682617,
-39.2192459106445,
-37.7522811889648,
52.9412612915039,
-12.9992752075195,
-22.5026855468750,
-1.37962460517883,
16.5472316741943,
4.11930036544800,
-43.4981498718262,
54.5149955749512,
21.3920288085938,
-44.0837059020996,
-8.03339862823486,
-31.6301460266113,
11.5731363296509,
4.65435552597046,
-23.4623641967773,
-18.9900989532471,
1.07826876640320,
-18.6207733154297,
-12.5312376022339,
30.7037582397461,
-14.8437662124634,
14.8125648498535,
-32.5639762878418,
8.85624027252197,
74.5051269531250,
-35.8675155639648,
-4.80896711349487,
22.4177265167236,
-40.2750396728516,
-23.8771095275879,
-6.54133033752441,
-40.0784721374512,
-5.24154424667358,
-0.225512430071831,
-13.5815525054932,
26.5088558197022,
17.0209846496582,
-9.39623260498047,
2.04764604568481,
-7.59255790710449,
-16.3406829833984,
-16.2651309967041,
-30.1690387725830,
-5.40741920471191,
-21.9405231475830,
-4.17014884948731,
25.3802204132080,
-11.4433956146240,
18.7834033966064,
31.2297210693359,
-22.4154167175293,
-4.55772209167481,
-15.1064910888672,
-10.9940719604492,
10.6659421920776,
-37.1724510192871,
12.5592727661133,
-5.86482238769531,
-5.72852849960327,
4.29291820526123,
-43.6821517944336,
-26.9477653503418,
-7.74763536453247,
36.0550003051758,
-5.96304988861084,
-27.8914680480957,
-5.14434528350830,
-18.7096080780029,
-10.4437847137451,
26.5498867034912,
2.32072162628174,
-9.09551525115967,
25.0212173461914,
7.24724960327148,
-15.0775432586670,
-13.9278850555420,
-6.29338312149048,
-20.6590099334717,
13.5227327346802,
-10.8485813140869,
-27.1963615417480,
-30.2956085205078,
-26.5661907196045,
-20.0296096801758,
-19.3415412902832,
11.6472311019897,
-23.0843143463135,
3.83851790428162,
-18.6402854919434,
3.61521196365356,
42.9350929260254,
5.17150974273682,
-26.7762031555176,
-9.52454376220703,
13.0875205993652,
-42.4511413574219,
-20.3791637420654,
6.97961759567261,
24.8615207672119,
17.3693084716797,
-6.55451393127441,
-24.1326427459717,
20.7139129638672,
18.5571632385254,
8.82409572601318,
12.5650043487549,
-18.0755176544189,
37.8599052429199,
-35.0525093078613,
-32.9750785827637,
13.8426733016968,
5.16831350326538,
14.2390871047974,
-0.411822378635407,
50.3194580078125,
8.35631084442139,
-27.0998477935791,
33.2913780212402,
-1.94983851909637,
-35.9735755920410,
41.0831031799316,
-0.345307409763336,
-46.8943557739258,
41.6753311157227,
9.77535152435303,
-35.6717872619629,
7.77549695968628,
22.1736621856689,
-28.4479598999023,
-11.2669954299927,
39.5079765319824,
-43.0097770690918,
-20.0955390930176,
38.9877738952637,
-1.49753129482269,
-22.9849014282227,
-39.8519477844238,
10.4614276885986,
19.9862804412842,
-64.6659698486328,
-14.8240804672241,
11.7097282409668,
-17.4923477172852,
22.4426403045654,
-15.7671022415161,
3.14626240730286,
8.13570022583008,
5.51454687118530,
23.7838668823242,
23.5691394805908,
29.7500896453857,
-27.7898921966553,
33.1532669067383,
44.9795494079590,
-1.11360859870911,
-0.538894534111023,
-12.6662778854370,
-1.20559179782867,
-4.55489873886108,
29.3021831512451,
9.61583995819092,
0.687260627746582,
24.8305511474609,
-26.5790538787842,
-5.83551263809204,
44.3963088989258,
28.9944267272949,
4.33051538467407,
-13.6204805374146,
27.5521659851074,
27.7557678222656,
-19.8879528045654,
8.64060115814209,
-21.2537021636963,
-25.3037185668945,
26.9289932250977,
16.4875507354736,
-10.3928537368774,
-14.9979753494263,
31.6149272918701,
-16.0222835540772,
-21.0660667419434,
63.2795753479004,
13.3332672119141,
-30.7518196105957,
2.50445485115051,
29.8600311279297,
2.90281414985657,
8.78733253479004,
42.8778152465820,
25.7068519592285,
8.32223510742188,
1.74737083911896,
-17.6913089752197,
-27.9932327270508,
-8.97988319396973,
10.2673921585083,
19.7252941131592,
-17.4789485931397,
12.8384351730347,
15.5169963836670,
-39.1878852844238,
-13.4920434951782,
6.81678962707520,
44.9434776306152,
6.81363773345947,
-26.0514926910400,
23.5645713806152,
-16.0508251190186,
18.3774700164795,
51.6315689086914,
-10.5541982650757,
17.7992420196533,
4.90346384048462,
8.63084793090820,
12.4680948257446,
-12.8069620132446,
21.7392673492432,
-26.0396671295166,
-18.4384593963623,
29.3126964569092,
31.2343940734863,
-12.9140024185181,
-41.9402580261231,
11.2320880889893,
-13.4443130493164,
-10.1053724288940,
-16.1559085845947,
-27.7745819091797,
-18.8837928771973,
-14.0774602890015,
33.6716384887695,
-18.3991069793701,
17.2222518920898,
15.8504810333252,
-30.2103137969971,
16.8484420776367,
22.2709388732910,
13.4258003234863,
-39.2771568298340,
-0.193566933274269,
-11.1266593933105,
-38.9978981018066,
10.2500152587891,
-1.79606962203980,
10.9706144332886,
-16.9794139862061,
-25.2393951416016,
-10.5540409088135,
-11.3098306655884,
15.0777940750122,
-0.869257748126984,
-15.2157220840454,
-6.78598785400391,
17.6222610473633,
12.9215555191040,
22.3729114532471,
33.4950981140137,
-7.32960939407349,
19.4073734283447,
40.9770774841309,
5.04345798492432,
-27.5465278625488,
27.0861110687256,
30.1073055267334,
-42.9235229492188,
27.8757495880127,
18.0915260314941,
-26.5140857696533,
22.1238632202148,
5.85070705413818,
24.1908817291260,
26.8938217163086,
23.2929382324219,
-10.2638292312622,
-32.4434738159180,
44.0103797912598,
27.4056053161621,
22.7975635528564,
-12.0860319137573,
-12.4288721084595,
34.4975433349609,
30.3656101226807,
26.0414485931397,
6.16343641281128,
18.8608493804932,
-28.2363376617432,
14.6515140533447,
28.9474716186523,
1.89795351028442,
26.0606136322022,
-41.2707748413086,
-3.64585375785828,
17.4573497772217,
-37.0676193237305,
26.1158485412598,
10.1893692016602,
-49.4713134765625,
31.8559722900391,
17.5845966339111,
7.16634464263916,
23.8950576782227,
-28.8386516571045,
9.59716129302979,
27.3900165557861,
9.51884937286377,
-11.6409769058228,
-16.4686698913574,
17.8845672607422,
33.6248016357422,
-15.1935968399048,
4.64526844024658,
38.2624130249023,
-26.1489543914795,
9.02851676940918,
46.5695686340332,
26.5920772552490,
15.3468723297119,
-20.2899093627930,
-7.72971057891846,
34.8299598693848,
11.9759502410889,
14.1732368469238,
41.2327194213867,
18.0833930969238,
-11.1004705429077,
-16.6119232177734,
46.0420303344727,
27.9604053497314,
-34.8333129882813,
36.5206832885742,
7.26155710220337,
-35.4244651794434,
34.9963455200195,
10.0410690307617,
-3.45217370986938,
3.02426314353943,
0.0132321445271373,
2.91524100303650,
-30.0694408416748,
-1.65815794467926,
12.4286317825317,
-28.5618209838867,
-23.8109569549561,
-6.29429578781128,
-17.7697963714600,
-21.8683795928955,
16.8359985351563,
17.7372055053711,
4.52308082580566,
18.4917068481445,
-28.1163940429688,
-24.0025844573975,
7.28488636016846,
19.2824916839600,
28.4343605041504,
-26.3915309906006,
-3.25610566139221,
28.5759792327881,
13.5248384475708,
30.4617652893066,
-16.3457183837891,
-11.5374078750610,
15.2778816223145,
-19.6967544555664,
7.45686531066895,
-1.78377223014832,
-32.1636352539063,
-23.5285530090332,
-17.6806144714355,
-22.1003189086914,
-30.8807773590088,
-21.8040637969971,
-19.5172042846680,
-31.2076168060303,
6.53088712692261,
36.3771476745606,
-28.0376205444336,
-0.267573833465576,
33.2039222717285,
7.55253601074219,
6.34864521026611,
19.1113224029541,
36.3907012939453,
7.69090604782105,
20.9138965606689,
2.04254102706909,
-12.5686445236206,
-10.1998424530029,
23.1994037628174,
7.27666616439819,
-48.4601097106934,
-9.91419219970703,
-16.1376037597656,
22.9948139190674,
9.67905521392822,
-7.63198614120483,
28.7836704254150,
-7.07011795043945,
-3.59912276268005,
30.7672233581543,
13.2253885269165,
-32.5454139709473,
-5.26397800445557,
44.5439643859863,
16.5689067840576,
-22.7577152252197,
12.0111980438232,
0.549745261669159,
-7.78720045089722,
14.3753442764282,
11.0116481781006,
33.8729438781738,
1.81982374191284,
-1.78935420513153,
23.9262256622314,
12.7345266342163,
15.9941673278809,
-7.97344493865967,
-19.5765628814697,
0.0776306167244911,
17.2067298889160,
12.3198575973511,
1.58615207672119,
34.8991470336914,
4.46923875808716,
-36.7881507873535,
28.8522586822510,
36.9372596740723,
-32.3389129638672,
24.3023414611816,
11.3778905868530,
-40.1768989562988,
48.0933914184570,
-6.15051698684692,
-19.4377136230469,
52.8733901977539,
14.5491504669189,
-34.8383598327637,
14.8958702087402,
48.8295669555664,
-39.7252349853516,
13.2864551544189,
36.3528213500977,
-27.5610275268555,
-38.5382270812988,
0.612359881401062,
30.2803688049316,
-32.7988052368164,
13.0941152572632,
21.6818847656250,
-9.89714050292969,
5.01282024383545,
23.2301025390625,
17.7978763580322,
-38.0810852050781,
-3.95224213600159,
22.7258129119873,
3.17437386512756,
0.611265778541565,
12.8265113830566,
-7.96545600891113,
4.95624780654907,
9.18110179901123,
-6.32189464569092,
41.9146690368652,
-21.1367797851563,
-12.2444295883179,
44.3027687072754,
5.25104618072510,
-0.101904667913914,
6.73009872436523,
36.0535240173340,
-13.2904491424561,
-15.7344875335693,
36.6585540771484,
-17.2266254425049,
-49.8696174621582,
6.46255826950073,
20.0545253753662,
-9.70818042755127,
17.5344181060791,
-13.4201202392578,
-11.6891136169434,
16.3464584350586,
17.3855457305908,
32.2477149963379,
21.1685256958008,
31.3699588775635,
28.4960575103760,
10.9891119003296,
26.7366657257080,
22.4847240447998,
-31.1256275177002,
10.9494981765747,
40.4906768798828,
-25.9574108123779,
0.945153951644898,
8.99514293670654,
-31.1094131469727,
-15.7277479171753,
-7.27432060241699,
-17.4369659423828,
-13.7894887924194,
4.54517936706543,
21.8238830566406,
-11.6835641860962,
-34.5559539794922,
21.4284801483154,
-8.67303276062012,
-18.4366874694824,
7.86018133163452,
-25.4232349395752,
4.18113327026367,
38.8589248657227,
12.2232770919800,
-30.2154808044434,
4.73428201675415,
-9.42853260040283,
-21.0658435821533,
-4.09140968322754,
-44.7428207397461,
-3.83501577377319,
5.11987304687500,
-16.8109703063965,
8.50979232788086,
6.60340452194214,
11.0801095962524,
-5.18262720108032,
-20.4560298919678,
-2.86176204681397,
-33.7854003906250,
-0.834759473800659,
42.6921195983887,
4.12193107604981,
-15.7484169006348,
7.67095994949341,
4.65117835998535,
-29.2812938690186,
-1.83252775669098,
28.2236957550049,
29.4311466217041,
-14.9295129776001,
-27.7081909179688,
6.19510030746460,
22.0707187652588,
-16.8049297332764,
-19.8331050872803,
17.5346260070801,
-2.26484465599060,
12.8355598449707,
-24.0266036987305,
-9.26936340332031,
11.2368144989014,
3.67237901687622,
3.53052663803101,
-9.46247673034668,
39.0425567626953,
-5.39155387878418,
7.77253866195679,
14.3300142288208,
-4.35456609725952,
-6.34127473831177,
-19.0713081359863,
47.9202766418457,
-9.03919792175293,
0.600556492805481,
26.7235774993897,
-23.9206752777100,
14.1537084579468,
30.7133502960205,
29.9014682769775,
-12.3605213165283,
5.31078243255615,
8.75975322723389,
-43.8789901733398,
17.4783267974854,
46.6899108886719,
11.8628149032593,
-10.1634941101074,
-14.4760198593140,
-15.4036378860474,
2.62026643753052,
21.4273986816406,
11.0290822982788,
2.92626500129700,
3.19758915901184,
3.54365348815918,
-22.2059478759766,
-0.546314477920532,
22.2163238525391,
-10.6589279174805,
5.93106317520142,
34.5662498474121,
-9.68225002288818,
-19.0919456481934,
28.5388584136963,
-8.20840454101563,
-33.6392288208008,
16.7298908233643,
38.5445747375488,
4.32470178604126,
-37.3300552368164,
-6.70534324645996,
1.20909011363983,
8.52724838256836,
31.9017505645752,
-0.353282094001770,
17.5186519622803,
-14.6989927291870,
-22.7453269958496,
0.382377475500107,
-6.60848045349121,
39.0453872680664,
-18.1815109252930,
-24.8498725891113,
11.4216394424438,
-14.8179931640625,
25.2690582275391,
-5.54724168777466,
-39.3524436950684,
24.7674789428711,
12.4577493667603,
-38.2653579711914,
-14.5681734085083,
35.4425506591797,
-1.96168911457062,
-46.1442947387695,
13.5438480377197,
7.51662349700928,
-18.9570426940918,
21.6314430236816,
-8.43882656097412,
-34.7665443420410,
3.74085283279419,
-33.9947166442871,
-25.3184642791748,
17.7435302734375,
-19.9726123809814,
12.9797315597534,
9.10889911651611,
17.4570884704590,
10.2945079803467,
-40.0193481445313,
31.6500301361084,
0.288049072027206,
-19.8046073913574,
40.2237014770508,
7.02033519744873,
-24.8948802947998,
-25.9776229858398,
5.93864917755127,
26.8113803863525,
-0.474661231040955,
-27.1709327697754,
19.7081642150879,
11.1768569946289,
-29.5134525299072,
21.1738071441650,
29.9279136657715,
4.27259349822998,
-30.3500728607178,
2.28946304321289,
45.8371887207031,
14.3192720413208,
21.1838836669922,
10.5261335372925,
-35.1474723815918,
-12.6242837905884,
43.9822235107422,
-5.08072090148926,
-16.0855274200439,
24.4984874725342,
-22.7654113769531,
-26.0399951934814,
12.9074335098267,
37.1948699951172,
11.1576652526855,
-5.98070287704468,
14.4994611740112,
27.1246623992920,
27.8690166473389,
16.5957298278809,
-0.0881865024566650,
-2.70435500144959,
15.2874898910522,
-24.3304538726807,
18.2073020935059,
1.75682079792023,
-14.4271135330200,
17.0931053161621,
-32.8657112121582,
21.7533645629883,
-16.3889579772949,
12.1821975708008,
49.0640945434570,
-4.78446722030640,
26.6135807037354,
-2.06749820709229,
-11.0458879470825,
2.48385596275330,
34.3937149047852,
-16.2518386840820,
-34.3866577148438,
2.03443956375122,
-28.1541061401367,
15.6445226669312,
10.7035512924194,
7.26260423660278,
9.44036483764648,
-24.2925472259522,
-19.7965660095215,
25.6415042877197,
23.4642467498779,
-40.7834510803223,
-10.9486036300659,
22.1092433929443,
33.8287048339844,
-1.97127187252045,
-12.7881851196289,
-3.18232369422913,
-14.3588008880615,
19.3540458679199,
-4.31701135635376,
32.7427597045898,
6.71550369262695,
-34.5015068054199,
14.1613063812256,
-17.4402809143066,
5.13644218444824,
41.0713844299316,
-0.398344069719315,
-18.4884796142578,
-11.4688596725464,
2.63958907127380,
11.4646415710449,
-30.2771987915039,
-21.0322856903076,
8.53752517700195,
9.52868652343750,
28.8212356567383,
-8.91525840759277,
-3.07199835777283,
-8.27201271057129,
-23.0949344635010,
28.8361358642578,
-23.4925193786621,
-20.0172424316406,
28.3748779296875,
-13.8788967132568,
0.341412752866745,
16.2153739929199,
-3.19973659515381,
-20.9169826507568,
-15.8371009826660,
-4.36615896224976,
7.40629768371582,
24.1292152404785,
3.27802944183350,
19.1816406250000,
18.5209960937500,
-24.9202919006348,
-12.9922809600830,
19.8273429870605,
26.5225677490234,
3.04836106300354,
-14.5079412460327,
1.35125994682312,
17.8553867340088,
11.3756027221680,
-0.386778503656387,
7.09140014648438,
-4.08723449707031,
-32.4957313537598,
-6.52288055419922,
33.4872703552246,
0.253668934106827,
-34.2360382080078,
30.6956176757813,
6.31040000915527,
-35.1844062805176,
29.5256843566895,
-5.80156183242798,
0.202654048800468,
14.3849430084229,
-15.4762926101685,
9.03829097747803,
-13.0445461273193,
-22.1255874633789,
-6.12983369827271,
-24.4613151550293,
-34.1501235961914,
-26.9614429473877,
-33.1429138183594,
-15.8559741973877,
-8.02709674835205,
11.6715898513794,
-10.1169357299805,
-19.5020542144775,
37.9177818298340,
-1.25326120853424,
7.79214906692505,
34.5355606079102,
-12.2545509338379,
16.2421627044678,
50.1131248474121,
-5.56498003005981,
11.8088626861572,
35.7359390258789,
-18.6295070648193,
-17.4032936096191,
10.0346021652222,
2.70508956909180,
-33.8699874877930,
1.48729193210602,
3.12246894836426,
-17.8282585144043,
8.94549179077148,
-24.3599433898926,
-1.02241873741150,
4.26576852798462,
-23.1168956756592,
12.6948080062866,
3.26439857482910,
1.79880642890930,
29.3934059143066,
27.4693851470947,
18.7232227325439,
-5.05343723297119,
-36.9944229125977,
10.1541576385498,
21.2088680267334,
-37.3929557800293,
-21.6423778533936,
2.96084737777710,
-3.10760068893433,
20.8419246673584,
9.56902503967285,
-32.5125656127930,
19.8531036376953,
22.6743240356445,
18.5174827575684,
-2.88315463066101,
-15.0822315216064,
15.3570299148560,
-25.4171695709229,
15.4516859054565,
6.54719543457031,
-32.4173736572266,
-26.8944129943848,
10.9989624023438,
-4.20636653900147,
-22.7976970672607,
16.9679260253906,
-1.97096145153046,
-6.68492269515991,
-27.1932640075684,
-8.49231338500977,
-16.3780727386475,
4.53772544860840,
5.38966274261475,
-27.0316963195801,
1.81698882579803,
-24.8387851715088,
12.9540004730225,
25.2408084869385,
5.93639039993286,
5.16703939437866,
19.9013175964355,
29.2806587219238,
-18.1445903778076,
-11.5784597396851,
-8.39513683319092,
0.586539328098297,
-24.9358005523682,
-4.90988874435425,
14.5603551864624,
-39.6212921142578,
-11.3906621932983,
-8.96525096893311,
-34.7977333068848,
-20.0786857604980,
27.9514331817627,
4.94637918472290,
24.4303131103516,
1.16475713253021,
-12.0607919692993,
9.87583065032959,
-25.3496398925781,
22.7834968566895,
-14.4726858139038,
12.3259420394897,
-14.5188302993774,
-8.69413089752197,
18.1966037750244,
-22.0156860351563,
31.7576293945313,
7.66221857070923,
-7.89448881149292,
-30.1216506958008,
0.642630159854889,
16.7099018096924,
-0.851865351200104,
22.3483695983887,
23.7117519378662,
-18.6913890838623,
-6.51368188858032,
53.9563407897949,
-5.55520057678223,
-4.50895261764526,
39.1663894653320,
25.6103477478027,
9.92652320861816,
-2.75146460533142,
-15.9853448867798,
4.45337772369385,
12.2806930541992,
-10.0938835144043,
18.1936550140381,
19.5703029632568,
1.00224566459656,
-26.7876815795898,
-2.33909368515015,
19.6898040771484,
-27.6060981750488,
12.0873651504517,
8.58300495147705,
-30.5410385131836,
-10.5505599975586,
15.6999950408936,
6.42710304260254,
-31.0935745239258,
12.8458633422852,
33.1475982666016,
7.09364700317383,
-13.7837009429932,
9.64437580108643,
22.4970474243164,
4.50927305221558,
37.8940353393555,
10.9739084243774,
-16.8655319213867,
23.2636089324951,
25.0881919860840,
-25.1129055023193,
-14.2114200592041,
31.6852302551270,
18.4327640533447,
4.46138191223145,
18.8501415252686,
6.45464181900024,
-9.26924419403076,
-5.84327077865601,
2.26711463928223,
9.19649505615234,
-22.1746120452881,
-18.7694625854492,
22.5938568115234,
-1.25701570510864,
-3.37899780273438,
-2.70878553390503,
-10.8580541610718,
47.5868988037109,
-8.62774753570557,
-21.7719917297363,
29.6471061706543,
-34.2081565856934,
-29.7079734802246,
-16.1435050964355,
4.82861757278442,
19.2196731567383,
-30.6745872497559,
-22.6533527374268,
4.41509580612183,
-3.17649078369141,
-20.9041843414307,
-23.4563694000244,
2.18282103538513,
10.2583026885986,
-27.0415554046631,
-18.6152400970459,
1.36975431442261,
13.2832393646240,
4.42517995834351,
-28.2910270690918,
23.5049343109131,
24.6025581359863,
16.1588516235352,
9.23380947113037,
-0.0411111116409302,
26.5294284820557,
-24.6952819824219,
14.1911191940308,
12.2111196517944,
-33.2158851623535,
-10.7036476135254,
-36.5723037719727,
-21.9253845214844,
17.4661693572998,
20.4162349700928,
3.82234358787537,
15.7426185607910,
12.7613077163696,
8.54984664916992,
17.0072879791260,
18.5991916656494,
-14.3791608810425,
-15.5854167938232,
47.7824935913086,
24.3223400115967,
13.0988759994507,
3.33672332763672,
-23.4814262390137,
25.7060604095459,
20.1315402984619,
-30.3294391632080,
17.9912338256836,
22.4697074890137,
-15.1380853652954,
2.10838937759399,
-14.3152666091919,
-5.91825103759766,
-20.0417938232422,
2.02819705009460,
7.46972990036011,
-37.8385047912598,
19.3198223114014,
-7.50746631622314,
-22.8979721069336,
24.7601737976074,
-22.8777370452881,
-29.0426273345947,
-27.4332523345947,
-27.5984573364258,
16.0589733123779,
21.0895195007324,
5.11637544631958,
-22.5646572113037,
-19.1789302825928,
2.19368028640747,
7.58502149581909,
-0.00143754936289042,
30.9161014556885,
-1.96230304241180,
-27.7579669952393,
33.2439651489258,
-13.2346296310425,
12.5587949752808,
29.5671043395996,
14.3326930999756,
10.3873891830444,
-12.6271333694458,
23.2129077911377,
1.91580271720886,
-33.0194282531738,
-20.0421352386475,
28.1036262512207,
-29.4700508117676,
-9.62427806854248,
14.9432277679443,
-20.9654293060303,
38.6564826965332,
-24.9738044738770,
11.1340827941895,
14.5254764556885,
-27.4104118347168,
13.8307762145996,
-29.9081535339355,
18.8934459686279,
17.9422798156738,
6.47493648529053,
-3.46145772933960,
-14.2376651763916,
16.4938964843750,
-20.3614253997803,
8.05983543395996,
2.05856442451477,
-11.8274431228638,
-20.5829925537109,
-15.4316577911377,
-10.6792993545532,
-27.4932346343994,
15.5181999206543,
-24.3337898254395,
-26.8648815155029,
-20.6928234100342,
-25.0770568847656,
-12.3488779067993,
-3.38976716995239,
13.4771308898926,
-27.5009632110596,
18.9642047882080,
1.11395144462585,
5.33127832412720,
5.42323970794678,
-22.7359752655029,
19.7185611724854,
-24.9417343139648,
26.6298065185547,
30.1345577239990,
-10.1179580688477,
-8.02957534790039,
9.62141418457031,
7.16439247131348,
-43.2506980895996,
21.0993652343750,
21.6867961883545,
-35.8644218444824,
-12.6173419952393,
-23.6020412445068,
-12.2113037109375,
22.3404998779297,
-22.9241027832031,
-9.14805793762207,
-14.9672183990479,
-3.74244070053101,
8.85451126098633,
-13.5806417465210,
26.1782341003418,
-15.3396062850952,
-1.25035297870636,
15.0909452438355,
-22.5807495117188,
-6.97230243682861,
-13.9866199493408,
-15.0761146545410,
18.0184841156006,
-3.25846719741821,
-31.3470249176025,
10.8548536300659,
-1.13525903224945,
-18.0344467163086,
17.0641403198242,
-1.71524322032928,
-2.65254950523376,
28.2827224731445,
-3.43465209007263,
4.91166591644287,
1.32245886325836,
-19.0836906433105,
8.69983005523682,
-20.5806751251221,
-3.58645176887512,
8.05655860900879,
-14.8186540603638,
17.2919979095459,
26.8744373321533,
8.86228466033936,
-2.90993118286133,
19.7389888763428,
2.05794858932495,
-18.4214687347412,
-3.89970088005066,
-20.4647369384766,
-9.24400043487549,
-23.8164310455322,
-22.3000335693359,
30.5448970794678,
-8.91989135742188,
-28.0237808227539,
24.6887016296387,
-8.36292552947998,
-26.1054401397705,
24.6697921752930,
16.0266475677490,
13.9967184066772,
4.66105747222900,
0.332176506519318,
26.5747051239014,
-10.7285099029541,
-15.0964126586914,
4.63415670394898,
0.945755720138550,
7.74087190628052,
-14.4993982315063,
-7.84961080551148,
-12.4330863952637,
-32.3877906799316,
-21.4362049102783,
-11.4925823211670,
12.6977281570435,
-31.9536991119385,
-7.55315303802490,
16.4961071014404,
-39.2677688598633,
-4.16365718841553,
4.55637598037720,
10.6238746643066,
23.6459598541260,
12.9207286834717,
-6.27499771118164,
-0.972785353660584,
5.44523239135742,
-14.9432029724121,
21.0569915771484,
20.6941337585449,
-32.0028648376465,
9.88490676879883,
21.7998771667480,
-26.1667804718018,
11.9860906600952,
-10.4873304367065,
-12.4181213378906,
-10.7451572418213,
-12.4588804244995,
17.2208423614502,
6.20272731781006,
9.09977340698242,
-17.9116001129150,
20.1641159057617,
18.0668411254883,
-4.96313667297363,
-12.3284387588501,
-25.6053581237793,
8.65025043487549,
-20.0435562133789,
-21.7468738555908,
19.4760150909424,
13.8485507965088,
-23.6313591003418,
-21.0246620178223,
10.9219856262207,
26.0071048736572,
-7.84352731704712,
-5.55696630477905,
33.6771240234375,
0.344093531370163,
-0.515560507774353,
-28.0989055633545,
-1.60441935062408,
16.5476608276367,
-38.6105422973633,
15.6812038421631,
-14.4131612777710,
-12.8505744934082,
14.9721279144287,
-18.6745071411133,
8.09883022308350,
13.3245363235474,
12.2064743041992,
-1.49987447261810,
-18.6997966766357,
-17.4515552520752,
18.4576187133789,
-3.56824064254761,
-28.7805442810059,
4.28110551834106,
-4.14887571334839,
-3.37061214447022,
5.18401288986206,
-5.90300989151001,
-22.4358463287354,
-26.5049495697022,
-24.9957580566406,
14.8527326583862,
0.333351343870163,
-11.1001062393188,
44.1502494812012,
-17.9893989562988,
-18.8261833190918,
26.2734889984131,
-34.9380416870117,
-11.3412818908691,
22.7750873565674,
1.56538748741150,
15.6769857406616,
-4.78402471542358,
-29.2889537811279,
-4.08860111236572,
-2.02425813674927,
-3.20517206192017,
34.2790298461914,
7.83971691131592,
-7.68853330612183,
35.7311172485352,
5.08200597763062,
-10.7977161407471,
3.62767100334168,
4.21016931533814,
20.3933963775635,
-15.2165069580078,
-19.8094177246094,
27.8119468688965,
-1.44237756729126,
-20.5643863677979,
-10.9800348281860,
-7.92266511917114,
-3.31091141700745,
-24.1190223693848,
-5.11665773391724,
25.3661670684814,
-14.2544498443604,
-34.3246536254883,
33.0230598449707,
4.50281381607056,
-23.7316799163818,
19.4604663848877,
14.1409807205200,
8.33534908294678,
-10.9357395172119,
18.2782936096191,
22.4503021240234,
26.7349472045898,
-6.09768247604370,
-13.9916048049927,
15.6144475936890,
-25.3974685668945,
0.168135121464729,
-8.78742122650147,
20.0906906127930,
16.4239921569824,
-3.57160735130310,
8.06251335144043,
6.21539497375488,
19.9665355682373,
-8.01841735839844,
7.35344552993774,
6.86075401306152,
6.04974508285523,
-10.2932968139648,
24.6837615966797,
21.3047676086426,
-17.0232257843018,
28.4209575653076,
-1.48077344894409,
1.51941776275635,
-4.32283782958984,
6.04712772369385,
1.14026129245758,
-24.7546710968018,
20.6981296539307,
-6.43531179428101,
14.4707422256470,
-8.59122943878174,
-26.8045272827148,
-0.0377286151051521,
-20.3161697387695,
-6.89129877090454,
-12.2970657348633,
-12.6170444488525,
-1.75302016735077,
-0.374833852052689,
-32.3774986267090,
14.9946470260620,
36.7467155456543,
-14.9234542846680,
-31.8292560577393,
18.9376506805420,
19.2537250518799,
-17.3887310028076,
29.8600425720215,
-10.7253351211548,
-30.2064590454102,
-9.89843940734863,
18.7459125518799,
-14.5398244857788,
-15.4513711929321,
17.4499568939209,
-34.5468482971191,
-2.27357888221741,
6.11098432540894,
9.57804393768311,
11.0018415451050,
-9.30159664154053,
22.3845157623291,
23.3864212036133,
-1.81999683380127,
26.2816085815430,
14.1944236755371,
-18.2781848907471,
31.6613788604736,
4.68530654907227,
-12.7971057891846,
35.5508689880371,
8.34074783325195,
17.5532779693604,
24.5517597198486,
2.95666694641113,
26.9204845428467,
21.6522293090820,
-8.96233654022217,
-10.4237108230591,
26.0317478179932,
7.27494096755981,
7.57488059997559,
16.2558498382568,
-15.9359588623047,
15.0370941162109,
-14.6569547653198,
-0.298075675964355,
37.0434379577637,
13.9846849441528,
21.0238323211670,
-1.90081131458282,
0.192105934023857,
13.8877420425415,
-2.23875570297241,
-26.8155364990234,
16.4000701904297,
25.8692226409912,
-21.5418663024902,
-13.6691827774048,
-10.6583309173584,
-14.3551111221313,
-4.28114891052246,
14.4496059417725,
-13.2878189086914,
1.35218834877014,
3.55556988716126,
-32.2926025390625,
10.0335817337036,
-1.02146363258362,
-11.2816267013550,
-0.865216195583344,
1.22166883945465,
17.1621208190918,
-3.60858702659607,
-11.9905691146851,
-21.0767459869385,
-6.17277240753174,
-0.249894261360168,
2.64022159576416,
24.2323570251465,
9.80699634552002,
-18.0533008575439,
-17.9622364044189,
-5.37394380569458,
-6.36622095108032,
24.0009822845459,
23.8940849304199,
19.8296413421631,
-1.57826042175293,
-25.3956031799316,
9.30631732940674,
14.8580293655396,
4.66014003753662,
15.6360416412354,
22.5537757873535,
-1.13037323951721,
17.3941154479980,
25.0518894195557,
-23.8824424743652,
7.72076654434204,
14.2538089752197,
-29.2453193664551,
-4.02334547042847,
8.83682727813721,
33.4760246276856,
0.556798756122589,
-8.55740451812744,
19.1089305877686,
-19.9025936126709,
26.0420436859131,
9.37463283538818,
-4.90031623840332,
17.7622947692871,
-27.6876068115234,
-7.23010396957398,
11.8909959793091,
-13.8110694885254,
-7.59025287628174,
17.0704994201660,
-5.79934406280518,
13.5666904449463,
28.6914501190186,
-8.26761722564697,
15.1130571365356,
2.09088516235352,
-7.95709228515625,
18.2263946533203,
26.3717117309570,
4.22112417221069,
21.7769260406494,
20.7041549682617,
-15.4830856323242,
24.8289165496826,
-4.91173028945923,
10.5913276672363,
14.8637790679932,
8.06098842620850,
13.8839988708496,
-32.2044639587402,
7.43597841262817,
-10.7055149078369,
14.9050674438477,
-5.15843343734741,
-35.4184455871582,
32.9837455749512,
-5.15597963333130,
-24.1048641204834,
-20.3423576354980,
0.946358203887940,
-13.9656686782837,
-31.1457405090332,
-3.57233381271362,
8.10407257080078,
21.3589668273926,
-20.3788013458252,
2.99781465530396,
-7.40329933166504,
-5.36411046981812,
39.5504226684570,
-0.235914349555969,
6.89485311508179,
22.0344009399414,
21.5159225463867,
-7.12524986267090,
12.3262138366699,
16.7736949920654,
-21.2346286773682,
13.7077369689941,
0.567478179931641,
1.52295100688934,
8.48620700836182,
0.692824721336365,
-5.98564338684082,
-27.5291175842285,
-19.6831321716309,
-24.4350700378418,
14.2786159515381,
23.9131717681885,
-15.0554256439209,
-12.0244636535645,
-8.04517650604248,
-25.4234256744385,
-9.33314037322998,
9.58222961425781,
-20.7774200439453,
-23.5910530090332,
13.8576927185059,
24.7138175964355,
-10.0906038284302,
19.1985607147217,
0.0918249785900116,
-25.3875732421875,
16.8374462127686,
14.7375888824463,
20.9513206481934,
-8.55035591125488,
-17.6120586395264,
-4.05933570861816,
16.9742832183838,
20.7980003356934,
-1.96362698078156,
-10.4667015075684,
-25.7866420745850,
-23.8157024383545,
-24.7160968780518,
-4.43239593505859,
19.6425609588623,
0.152455434203148,
-17.2631187438965,
-1.44207477569580,
12.0740308761597,
14.1812248229980,
6.94061040878296,
-0.603748738765717,
1.53843677043915,
20.8344154357910,
14.1802701950073,
6.41176891326904,
32.4230575561523,
-10.6152896881104,
-4.22898149490356,
28.1872539520264,
8.98420619964600,
8.23327255249023,
-7.69501256942749,
20.4300231933594,
14.0572929382324,
-1.88424599170685,
31.2791576385498,
27.6490554809570,
-11.4748830795288,
-20.3866138458252,
20.2736568450928,
-11.6014003753662,
-7.53917741775513,
19.3355350494385,
2.11226963996887,
-10.6245212554932,
-20.1795883178711,
28.3053264617920,
-6.48655033111572,
-8.64759349822998,
38.5954513549805,
-13.4827527999878,
-27.8526763916016,
10.0570478439331,
33.3083801269531,
11.7622575759888,
17.4425640106201,
6.83068132400513,
-24.1703453063965,
24.9535446166992,
11.4449329376221,
-13.7339992523193,
33.2361831665039,
-4.33516359329224,
-3.92650771141052,
21.8136596679688,
-2.65678739547730,
28.1603431701660,
-13.1532640457153,
-27.5445709228516,
26.4366722106934,
-14.9533882141113,
-7.62124633789063,
1.67193830013275,
-24.1260776519775,
32.1508026123047,
0.188397064805031,
-12.9206933975220,
7.65204715728760,
-24.6662788391113,
12.3766908645630,
-4.39251279830933,
9.82643127441406,
4.65710973739624,
-40.4368782043457,
14.9482135772705,
14.9650020599365,
23.8255176544189,
2.49639034271240,
-8.37303256988525,
-1.11634612083435,
-8.24216079711914,
32.9099884033203,
-8.73560619354248,
-20.2476215362549,
-5.52011013031006,
24.3019046783447,
-1.48362362384796,
10.6109981536865,
13.2202692031860,
-25.7206745147705,
27.3096618652344,
-26.2661991119385,
12.4328804016113,
10.2962303161621,
-33.6879615783691,
19.4189548492432,
4.24211406707764,
-18.7397766113281,
-6.85643529891968,
21.0964469909668,
-0.368064790964127,
-16.9485759735107,
-19.9031162261963,
8.36935710906982,
-7.45246648788452,
-19.5736217498779,
14.1715679168701,
-12.5195789337158,
10.3285350799561,
-13.4356384277344,
-16.8385715484619,
35.7100944519043,
0.522211492061615,
6.42036056518555,
22.0991554260254,
-11.8651504516602,
-19.7291698455811,
20.0816078186035,
13.1843986511230,
-6.59588623046875,
4.01377868652344,
4.65098905563355,
-2.68815398216248,
0.573758721351624,
21.9102897644043,
-4.83070182800293,
15.2352523803711,
4.16230058670044,
-32.5788879394531,
8.05866241455078,
23.6409931182861,
8.52495956420898,
-36.9233322143555,
4.51769828796387,
29.6644706726074,
-28.1094341278076,
1.31539022922516,
-8.78763294219971,
-33.3881187438965,
0.190581977367401,
-12.4018287658691,
-6.76194524765015,
29.0117931365967,
4.21596097946167,
8.57906723022461,
14.4222612380981,
-9.32635021209717,
18.6661071777344,
5.67711877822876,
16.2914810180664,
0.549726486206055,
-31.1873817443848,
2.17107081413269,
-20.2370853424072,
-1.52700591087341,
-8.18674659729004,
-24.2923107147217,
-18.7935314178467,
-31.5822143554688,
16.8503513336182,
6.13690090179443,
15.6040544509888,
-3.26556658744812,
-29.5253086090088,
26.8293895721436,
-11.2255020141602,
-17.4696674346924,
11.4252462387085,
-6.97611856460571,
-12.0114459991455,
-3.79010677337647,
17.8174419403076,
7.28921937942505,
-22.6437015533447,
-7.56647729873657,
-5.28239536285400,
-32.3395195007324,
-3.51949691772461,
-4.11779451370239,
-25.8980331420898,
2.39336991310120,
4.15372800827026,
-18.9955635070801,
-20.3170623779297,
18.3190364837647,
18.3934516906738,
-6.16725730895996,
-5.68223476409912,
-22.3699417114258,
-2.52390623092651,
22.7877407073975,
20.1812763214111,
3.44378042221069,
-13.7508964538574,
-15.7335834503174,
-7.62638902664185,
18.7008724212647,
17.4570808410645,
-0.270043134689331,
-7.42402458190918,
7.92286396026611,
-3.79248452186584,
-17.4105663299561,
27.8165302276611,
-3.56274986267090,
-38.4379653930664,
11.1145334243774,
20.0579910278320,
11.9702329635620,
3.02342629432678,
20.8324985504150,
18.2021064758301,
-30.7872161865234,
15.6015129089355,
37.6613731384277,
-0.282816201448441,
-2.97327589988709,
-16.8322219848633,
-19.3628387451172,
0.975640475749970,
10.3704795837402,
-3.71790218353272,
-27.2728729248047,
-22.9918537139893,
-14.7098321914673,
15.2960186004639,
13.1331663131714,
-28.9870586395264,
-6.61617183685303,
-4.90986633300781,
7.74289369583130,
4.21275329589844,
-7.36348009109497,
13.9692029953003,
-16.9127712249756,
19.8985519409180,
21.3792743682861,
5.14394092559814,
25.6515140533447,
-9.38750267028809,
8.77223587036133,
6.91683006286621,
0.867252469062805,
1.14284384250641,
-19.6846809387207,
29.6952724456787,
18.6933994293213,
-30.2399063110352,
20.2564392089844,
20.8861865997314,
-17.4148616790772,
15.5644702911377,
29.8195552825928,
13.8721342086792,
-5.04317378997803,
-3.27423715591431,
-0.520283639431000,
-10.4671955108643,
18.3994235992432,
21.3933582305908,
-9.52312755584717,
-13.3951196670532,
-15.2891731262207,
-6.82379198074341,
-4.55163240432739,
4.60021305084229,
13.6312913894653,
2.14720916748047,
-8.93512439727783,
-6.17260456085205,
10.5978727340698,
-13.3697204589844,
12.7799320220947,
18.9779644012451,
0.291616737842560,
31.9058971405029,
-3.64358258247376,
10.4872455596924,
13.3228082656860,
9.74615955352783,
11.5154953002930,
-23.1183910369873,
28.1235904693604,
7.90949535369873,
10.0021438598633,
1.66409361362457,
-15.4452323913574,
9.73046398162842,
-2.82605695724487,
-4.46143579483032,
-14.4705600738525,
7.50386285781860,
-25.5008087158203,
13.5277404785156,
6.96473932266235,
-2.60203313827515,
18.3312911987305,
-13.3378820419312,
12.8679199218750,
-21.8366775512695,
8.01418113708496,
22.5181808471680,
19.5422782897949,
-13.9560794830322,
-14.9667901992798,
16.5372066497803,
-19.0860137939453,
31.2892055511475,
-6.36365747451782,
-22.0181465148926,
17.2975292205811,
-18.3074111938477,
-15.9449672698975,
-6.25794506072998,
-5.35200262069702,
-30.0009231567383,
-4.27525854110718,
35.7674331665039,
5.62284088134766,
13.7169523239136,
1.75493037700653,
3.01038050651550,
19.0218467712402,
-8.39385032653809,
-18.2909564971924,
3.92852163314819,
31.7269630432129,
-16.8444519042969,
-2.48413252830505,
35.6211967468262,
-6.85415220260620,
-13.7164392471313,
21.3822231292725,
24.2249679565430,
-1.75205588340759,
9.62611103057861,
5.95454311370850,
19.4229106903076,
2.75406002998352,
2.82199692726135,
14.1288499832153,
6.60006618499756,
19.3828697204590,
-21.5991401672363,
6.70231723785400,
-1.93942928314209,
7.66877603530884,
35.3175277709961,
-25.0827407836914,
4.82835769653320,
28.0475311279297,
9.10477924346924,
15.3914937973022,
29.8721523284912,
18.7650108337402,
-26.9578723907471,
-7.60919427871704,
29.8077068328857,
5.79776763916016,
7.79309654235840,
0.606126010417938,
-34.5103302001953,
17.1598091125488,
8.83300018310547,
-18.1446380615234,
7.63492441177368,
-28.6522293090820,
-5.14206123352051,
12.9894828796387,
-5.04174232482910,
5.26430416107178,
21.1370506286621,
-9.54742527008057,
-8.31088352203369,
13.5809259414673,
-28.6151294708252,
11.1258249282837,
25.1407203674316,
7.11698818206787,
3.66925740242004,
-21.4472351074219,
-15.7894592285156,
-20.4071617126465,
-11.2200202941895,
11.2062368392944,
-2.75702381134033,
-2.17841982841492,
12.3293123245239,
-18.7166786193848,
-6.94948673248291,
23.0724792480469,
1.30201840400696,
5.11293458938599,
8.91902923583984,
19.4584503173828,
19.9052925109863,
5.46820354461670,
6.15364646911621,
-19.8104972839355,
19.1023368835449,
20.4939842224121,
-16.6066722869873,
8.69542407989502,
-9.42644500732422,
3.85920166969299,
6.44551658630371,
-5.57789468765259,
35.4377937316895,
7.11737489700317,
-14.8940353393555,
10.5464363098145,
-2.65497994422913,
-10.5640411376953,
2.20411920547485,
-5.25965595245361,
-6.90945005416870,
27.6877384185791,
-3.62806177139282,
-25.9920864105225,
33.3692131042481,
3.47761464118958,
-16.1622676849365,
26.2258377075195,
0.106320530176163,
3.26133394241333,
4.04668855667114,
-23.0383872985840,
13.4473524093628,
23.2032470703125,
5.01966619491577,
8.43256378173828,
-12.0746479034424,
-12.8303050994873,
13.9410724639893,
-10.7924261093140,
-20.3179664611816,
10.2712144851685,
-1.04710996150970,
-12.9361295700073,
8.75697994232178,
28.7784881591797,
11.2068490982056,
-8.17003917694092,
18.2429199218750,
29.1077098846436,
-10.2172851562500,
-12.0503044128418,
23.3468933105469,
-9.04949092864990,
-5.79069566726685,
16.6695842742920,
-4.73803949356079,
-20.3326358795166,
-13.6689958572388,
19.8842277526855,
-17.3964824676514,
-24.0907611846924,
-6.45304965972900,
-21.4403724670410,
-1.28435337543488,
-3.91841077804565,
-9.53448772430420,
3.78115367889404,
-13.4990520477295,
-15.2375335693359,
1.84109568595886,
-12.8168716430664,
-11.1183271408081,
4.98537683486939,
11.8886899948120,
-6.33382892608643,
7.81690788269043,
13.3287830352783,
-24.1355133056641,
-23.5761985778809,
1.48148190975189,
15.2316408157349,
-6.55698442459106,
10.3593912124634,
24.1393260955811,
3.74074482917786,
6.67864322662354,
17.6907825469971,
26.9619827270508,
0.163914278149605,
-26.3559741973877,
-0.729355931282044,
7.19540691375732,
5.27733802795410,
5.88599252700806,
-19.2183227539063,
8.95624351501465,
4.61729955673218,
-19.0662174224854,
20.2215061187744,
20.8125419616699,
4.85642337799072,
-15.3416481018066,
-0.462109267711639,
25.9270725250244,
-21.2495765686035,
-27.9225254058838,
5.91081762313843,
8.38543605804443,
9.32600879669190,
3.09307599067688,
20.9187183380127,
19.0256347656250,
-15.8676452636719,
-5.91844606399536,
-9.02760314941406,
-3.28787827491760,
-4.59294223785400,
-29.1846008300781,
4.26329088211060,
9.58828163146973,
-2.32905936241150,
12.3262939453125,
-8.35315704345703,
27.7980155944824,
16.5863857269287,
-32.4147109985352,
28.6248817443848,
12.6738862991333,
7.34408569335938,
22.5825481414795,
-23.4142379760742,
-4.68924236297607,
-12.4657745361328,
-21.6986541748047,
1.41956412792206,
-23.3018226623535,
-26.5638694763184,
4.44047689437866,
-17.9417762756348,
-32.2747116088867,
5.27740669250488,
7.51149892807007,
6.46787357330322,
-1.98798191547394,
-11.8779687881470,
-0.992505311965942,
8.44562149047852,
9.23121452331543,
-20.9028148651123,
13.3230171203613,
14.7098550796509,
-29.7634525299072,
-13.9179773330688,
-11.3041038513184,
-5.89850378036499,
-21.7249908447266,
-0.00393467117100954,
10.3540430068970,
-12.2972221374512,
0.941759169101715,
-0.784362196922302,
19.5017204284668,
-15.9798288345337,
6.20710039138794,
18.5366802215576,
-11.7463588714600,
32.5171928405762,
-3.01819944381714,
-5.69594621658325,
-15.7664270401001,
-28.9840373992920,
19.6407852172852,
19.9925670623779,
-8.48721122741699,
5.97084474563599,
21.7838115692139,
-9.27689933776856,
26.1027202606201,
18.5717296600342,
-10.8419609069824,
21.5570716857910,
0.176809966564178,
-16.4654445648193,
-0.469881266355515,
13.5149631500244,
22.9808750152588,
8.42692756652832,
-3.71860480308533,
4.66631269454956,
1.68195247650146,
-2.79683399200439,
-13.2033958435059,
-19.4351654052734,
-8.99984359741211,
-27.0980434417725,
-6.60610723495483,
-3.60464167594910,
-11.4437799453735,
17.0796070098877,
-0.295973658561707,
22.0171203613281,
16.0975513458252,
-13.4961738586426,
-10.7298326492310,
-13.1922760009766,
-3.51946640014648,
-20.6279621124268,
-14.6655178070068,
12.2515115737915,
17.9922084808350,
-7.17733860015869,
-16.3101863861084,
2.22085118293762,
8.06768703460693,
13.7704048156738,
-14.3343801498413,
-2.27221918106079,
14.6635198593140,
1.03178381919861,
5.86264610290527,
-1.30918705463409,
-0.117708392441273,
-0.899395167827606,
21.6051044464111,
-8.70476150512695,
-15.7362537384033,
33.2152214050293,
-14.0511989593506,
-5.28806543350220,
6.77640390396118,
-33.8534889221191,
-0.153466612100601,
-5.78566646575928,
-20.8761558532715,
17.3053455352783,
13.4160270690918,
-1.59285914897919,
5.84237051010132,
9.80221652984619,
-8.10615730285645,
-26.0944786071777,
-12.0508642196655,
4.59739923477173,
10.7784776687622,
-14.6371688842773,
0.123281426727772,
22.8792095184326,
-5.34928512573242,
14.0664520263672,
12.4881563186646,
14.1613216400146,
5.39453411102295,
12.7945175170898,
15.0127372741699,
-14.7469959259033,
25.2342720031738,
10.1273536682129,
-15.6597805023193,
-1.01932454109192,
18.8511848449707,
6.31393289566040,
-10.4257049560547,
-16.7909946441650,
-11.5027980804443,
-20.6708488464355,
-11.8286275863647,
21.9614505767822,
-19.1504878997803,
8.52635669708252,
-18.0007648468018,
-4.39299011230469,
31.3665657043457,
-37.6300239562988,
11.6242609024048,
13.3873853683472,
1.42604935169220,
16.5269908905029,
-13.4821586608887,
22.3635921478272,
17.0196228027344,
-5.33038425445557,
24.0581722259522,
27.4950523376465,
8.29490566253662,
7.22575616836548,
13.5276403427124,
1.22910594940186,
15.3405418395996,
22.6608848571777,
19.2348880767822,
3.26148462295532,
-13.3720731735230,
-3.00339508056641,
-20.7680797576904,
6.40321159362793,
35.2882995605469,
1.08216667175293,
-0.676487386226654,
5.92151069641113,
-8.98608779907227,
16.9180145263672,
25.2118930816650,
9.42304229736328,
20.4085884094238,
-7.57971286773682,
8.79069328308106,
10.8109970092773,
-0.563441634178162,
19.4842052459717,
-20.7533206939697,
-10.3420295715332,
4.10839891433716,
18.4495773315430,
18.7546157836914,
-24.7668533325195,
-5.38853311538696,
24.8998794555664,
2.97947287559509,
-19.9152755737305,
-11.4802179336548,
-7.92871141433716,
-14.2955951690674,
-1.29408121109009,
-8.51408195495606,
-15.0137310028076,
0.569567561149597,
-12.6144294738770,
9.01567745208740,
-16.2177429199219,
-7.92757320404053,
22.2314205169678,
-16.6855278015137,
-0.999287068843842,
-1.63438498973846,
6.93100500106812,
12.6062555313110,
10.1890783309937,
14.0513267517090,
11.9852724075317,
22.0637550354004,
17.6995792388916,
15.2760372161865,
20.5819854736328,
15.5056457519531,
-16.0618782043457,
0.906356632709503,
1.17519688606262,
-11.6841239929199,
-6.88371276855469,
-28.3682041168213,
6.56475687026978,
-8.42406463623047,
-23.3709602355957,
11.8716535568237,
10.9840116500855,
1.38827359676361,
-2.43442797660828,
23.6509723663330,
7.87743616104126,
-0.591735959053040,
-9.41720008850098,
-8.20167064666748,
18.5848274230957,
8.97678279876709,
5.26982116699219,
2.60110855102539,
-1.35821092128754,
10.2755670547485,
17.6139888763428,
-21.1447944641113,
3.74955344200134,
22.8955898284912,
-12.8836507797241,
0.632754206657410,
5.65944719314575,
-7.73139333724976,
-8.04318141937256,
25.7945404052734,
17.4281864166260,
-10.9473962783813,
17.4335536956787,
5.13484048843384,
-18.1734027862549,
12.5634546279907,
19.0796833038330,
11.0131101608276,
10.4416084289551,
19.3823299407959,
19.4109477996826,
-16.7764453887939,
5.51829195022583,
18.6635227203369,
-1.39087986946106,
9.31348609924316,
0.240906581282616,
4.37179565429688,
10.8861484527588,
-7.28016662597656,
-10.8031444549561,
-17.9556083679199,
-12.8716726303101,
5.25755023956299,
-23.0218982696533,
-12.2274961471558,
13.9385652542114,
11.8096036911011,
12.3090629577637,
-7.41919040679932,
-10.9696245193481,
12.9369125366211,
20.8801002502441,
13.6578340530396,
18.8678379058838,
-4.79812860488892,
11.2447452545166,
27.1995143890381,
-12.8844413757324,
0.230519577860832,
26.9343509674072,
-5.10071754455566,
4.67284631729126,
24.7734603881836,
-15.3011398315430,
-20.5449180603027,
4.95597600936890,
22.5659999847412,
1.12769067287445,
0.319641739130020,
-9.61391067504883,
5.24496841430664,
15.0463161468506,
-3.90428209304810,
1.52566027641296,
-16.8880844116211,
16.8522338867188,
-5.16850900650024,
0.247315883636475,
2.18966412544251,
-8.06823539733887,
25.5906829833984,
-15.9448652267456,
-0.421222537755966,
12.7682275772095,
14.0097208023071,
-7.18281793594360,
-3.89667153358459,
26.6096553802490,
-6.06015300750732,
-14.8328065872192,
-9.37955188751221,
28.8020915985107,
-0.585082948207855,
-26.4673862457275,
13.4705686569214,
-24.2514915466309,
-26.2368602752686,
-12.9130973815918,
-2.45564365386963,
7.41424131393433,
1.11970376968384,
18.9687919616699,
-31.3529148101807,
5.32613658905029,
20.2756576538086,
-29.7407951354980,
-0.0341851562261581,
-15.1332502365112,
13.0129985809326,
-12.1779642105103,
-38.8653373718262,
18.6989383697510,
17.1750907897949,
-5.70717668533325,
-4.90467214584351,
18.9661731719971,
-3.41112947463989,
-16.5413627624512,
24.1959266662598,
25.9338722229004,
-2.70001697540283,
-0.0302014779299498,
-10.1741971969605,
-4.09228563308716,
29.5811996459961,
-0.117914400994778,
-26.9234123229980,
17.8269710540772,
17.2516880035400,
-15.4021377563477,
24.4269542694092,
-0.625773251056671,
-27.6849403381348,
6.94326162338257,
-2.76025795936584,
-3.92632675170898,
-9.85756015777588,
-12.4381113052368,
-10.0355653762817,
-25.4700012207031,
-12.8001537322998,
12.1250095367432,
15.4902248382568,
5.21703767776489,
20.4325904846191,
5.15192604064941,
-13.0666007995605,
21.4479885101318,
-4.84783172607422,
-11.9639406204224,
12.0347080230713,
13.2478923797607,
12.0205039978027,
-21.3409080505371,
1.68361401557922,
13.5330219268799,
7.22787189483643,
9.04528903961182,
19.2595367431641,
13.9806795120239,
1.95353996753693,
21.7960681915283,
2.78765845298767,
3.68960499763489,
-11.5427360534668,
-4.75774002075195,
1.87976133823395,
1.40832293033600,
-3.80093240737915,
6.31638765335083,
15.4006690979004,
-19.0435237884522,
-10.3755178451538,
-15.7341384887695,
6.22290945053101,
-15.6125164031982,
2.58240747451782,
22.7186222076416,
-11.3405485153198,
18.4390754699707,
20.6533203125000,
-7.00991868972778,
-15.0190343856812,
17.1328697204590,
-15.4380254745483,
-13.5015621185303,
26.0047702789307,
-4.47312116622925,
-3.80049204826355,
3.64863324165344,
8.46854686737061,
21.5038814544678,
13.4952812194824,
15.0553903579712,
3.41560912132263,
-3.42005205154419,
27.4221000671387,
1.63323450088501,
-13.9472637176514,
-0.179366707801819,
-16.8626194000244,
-2.84086465835571,
11.8046007156372,
17.7637424468994,
-2.13709259033203,
-7.60079765319824,
8.79161548614502,
-17.8006172180176,
4.51402997970581,
26.0509567260742,
-10.1591796875000,
-16.4385700225830,
2.20650768280029,
8.89561462402344,
12.0319643020630,
15.9675321578980,
10.8423080444336,
-16.8259544372559,
-9.06159877777100,
2.35189175605774,
-18.1290779113770,
14.7830514907837,
-10.4929351806641,
-18.2396984100342,
14.2707405090332,
-9.95264625549316,
-3.97713398933411,
-3.43220901489258,
-9.29983520507813,
-7.38602495193481,
19.4284286499023,
3.14116287231445,
6.27621555328369,
23.0823516845703,
-21.0921974182129,
-1.05810093879700,
21.4471645355225,
4.71789741516113,
-16.3128337860107,
2.42987227439880,
5.16267108917236,
-19.0686073303223,
-9.02028369903565,
-6.20608520507813,
-3.79294848442078,
-13.1626615524292,
-18.6204586029053,
-0.204151526093483,
7.13574028015137,
17.7190055847168,
12.2434310913086,
7.21132659912109,
23.5998630523682,
-10.1457700729370,
-20.9555568695068,
-10.6096935272217,
-12.6389141082764,
-6.14979791641235,
4.24863862991333,
3.56886816024780,
-24.9734725952148,
-14.1393070220947,
-14.4707832336426,
5.66297435760498,
25.9198532104492,
-22.9094963073730,
-13.6037569046021,
25.1363468170166,
15.4792041778564,
12.1562967300415,
7.64394521713257,
12.5104494094849,
22.9355392456055,
-5.19483089447022,
17.6592483520508,
10.0523042678833,
-30.9394054412842,
10.5595512390137,
18.0953063964844,
11.7974386215210,
10.1332998275757,
-5.04205894470215,
8.91794395446777,
-21.3674316406250,
-13.1006698608398,
4.95584917068481,
-23.8916244506836,
10.2199077606201,
-4.29548835754395,
-17.6191730499268,
-18.0592784881592,
-10.0183963775635,
19.3933830261230,
-19.9224109649658,
-6.46033763885498,
10.0751876831055,
6.89029312133789,
-13.6894378662109,
-23.9587821960449,
-9.74865531921387,
-6.61667203903198,
23.6289672851563,
5.93526506423950,
-20.3550167083740,
-8.01454448699951,
21.9674587249756,
-3.12549972534180,
-7.24104928970337,
23.4514541625977,
-15.9802961349487,
-15.3888168334961,
-6.27655267715454,
1.62491679191589,
18.1560707092285,
-20.9709129333496,
3.76073145866394,
23.9306983947754,
-10.1715335845947,
10.3706026077271,
23.1635036468506,
2.44486713409424,
-28.7904644012451,
8.57470226287842,
18.6526985168457,
-22.4469661712647,
1.83873653411865,
-6.64582633972168,
-24.5743942260742,
2.32594037055969,
19.1447601318359,
-14.8875923156738,
-24.0562267303467,
-11.5609693527222,
0.348684757947922,
-1.96826636791229,
-4.91228723526001,
10.2085113525391,
-12.1250114440918,
-4.65635776519775,
-4.47353506088257,
-2.28475189208984,
16.6581001281738,
-7.19684839248657,
-33.5363845825195,
8.82329559326172,
10.8104867935181,
-18.3041763305664,
15.4537887573242,
8.95059204101563,
12.5520200729370,
-19.1756229400635,
3.68157029151917,
36.7982025146484,
-1.54281783103943,
16.4673576354980,
-7.35659456253052,
0.365705639123917,
0.180551439523697,
-8.25336647033691,
24.4298820495605,
11.9101829528809,
7.56046676635742,
-9.41052055358887,
-11.0191183090210,
-2.48169827461243,
2.16308522224426,
5.89605569839478,
-10.9466934204102,
4.98006820678711,
5.07778310775757,
2.38144540786743,
7.59668350219727,
9.30776882171631,
10.5067949295044,
1.68599867820740,
18.7067203521729,
2.90148353576660,
-15.0404691696167,
-8.24881839752197,
-12.3378314971924,
0.675969958305359,
11.4947004318237,
12.1473569869995,
-7.66005516052246,
1.95180165767670,
20.9540233612061,
-26.8147201538086,
3.63700914382935,
23.0937824249268,
-16.6493930816650,
-6.89379215240479,
12.4082403182983,
19.8929157257080,
6.87345218658447,
18.5537242889404,
6.99134969711304,
8.53010463714600,
6.26935148239136,
-12.8603172302246,
-0.588943064212799,
17.4229202270508,
6.97689628601074,
-6.04624891281128,
17.5653953552246,
-9.14617347717285,
-12.1244249343872,
5.51222991943359,
8.07398128509522,
-4.04879665374756,
-13.9587144851685,
-4.46925687789917,
-17.1527042388916,
8.22920513153076,
15.3071508407593,
-18.2109069824219,
-23.2588062286377,
10.1739091873169,
0.406555861234665,
-27.9096794128418,
-4.52571058273315,
-4.72099637985230,
-7.30143737792969,
-11.9390697479248,
-0.385359734296799,
19.7328243255615,
5.93269968032837,
-1.18802773952484,
-14.1358575820923,
13.4408655166626,
27.9551410675049,
-16.2178459167480,
-14.0081481933594,
1.94978559017181,
-20.0069370269775,
-23.0247726440430,
1.80854296684265,
-4.19077205657959,
1.86440598964691,
13.7582445144653,
-8.80486488342285,
-22.7058639526367,
-3.54696536064148,
14.6534385681152,
-8.96711730957031,
24.7420806884766,
11.4550485610962,
-26.4526500701904,
1.72918379306793,
7.66520977020264,
20.9726467132568,
-0.00830799713730812,
10.4347677230835,
-6.57306385040283,
-3.91526508331299,
8.34635543823242,
-13.1440496444702,
9.24168586730957,
-6.46936178207398,
-6.49715423583984,
-13.5714178085327,
7.82853555679321,
2.90206575393677,
-2.13528394699097,
18.5425472259522,
-4.28746652603149,
-8.85913276672363,
2.91454339027405,
21.5403213500977,
-9.81588268280029,
-12.0293979644775,
-8.45334434509277,
-22.6611976623535,
-9.31936740875244,
3.89847636222839,
5.84689140319824,
-16.1428871154785,
14.5276470184326,
0.378917098045349,
-26.5780181884766,
13.6319055557251,
7.10582208633423,
9.72482299804688,
-3.12316679954529,
-17.1181201934814,
10.2109889984131,
6.70801496505737,
-1.03705775737762,
-3.97107720375061,
-8.34234142303467,
-8.59613895416260,
-9.74724292755127,
-7.08062171936035,
16.7178134918213,
-5.73592042922974,
-33.0857887268066,
3.92601871490479,
17.1976509094238,
2.49262380599976,
-22.0629405975342,
6.54514503479004,
-4.52672767639160,
-11.4393892288208,
25.7542304992676,
-4.03793811798096,
8.45717811584473,
-11.9566564559937,
7.74303627014160,
16.6251068115234,
-6.15165805816650,
7.37611055374146,
-27.5562191009522,
15.7385177612305,
17.6209125518799,
0.548461616039276,
21.1649074554443,
18.9889774322510,
13.5100898742676,
-19.6114902496338,
5.21236753463745,
33.2427520751953,
-4.38602685928345,
-24.1487445831299,
13.3144321441650,
-5.37137794494629,
-12.8364410400391,
25.9478836059570,
-1.91995596885681,
15.7332229614258,
-0.260298401117325,
-8.20605182647705,
20.8626937866211,
3.43165397644043,
1.94014513492584,
-25.0965080261230,
-13.5509500503540,
-15.0597448348999,
2.61754560470581,
22.5613327026367,
-6.84441614151001,
18.7897605895996,
-3.39098262786865,
-3.01543760299683,
22.9713096618652,
7.32512426376343,
14.9781475067139,
-11.9811725616455,
24.5271072387695,
17.3983402252197,
-23.9236526489258,
18.4778938293457,
-1.96523582935333,
15.4842462539673,
-5.98198223114014,
-2.99740242958069,
15.0821380615234,
-13.4412012100220,
21.5803737640381,
-9.72645473480225,
7.92076826095581,
3.42830562591553,
-6.01194047927856,
25.8472290039063,
-10.3999805450439,
-17.3241348266602,
-10.1933746337891,
25.0316276550293,
7.25329256057739,
-15.6637916564941,
-12.1682033538818,
-15.5331192016602,
-4.16272830963135,
-17.0392456054688,
15.9598903656006,
-8.03927898406982,
-30.6003742218018,
-13.6832523345947,
-4.95384597778320,
13.2929983139038,
5.92003059387207,
-3.35610771179199,
-23.8896560668945,
20.2289161682129,
16.3184528350830,
7.28666496276856,
15.3454217910767,
-23.5236015319824,
12.7983865737915,
-1.79044961929321,
-20.7277984619141,
-5.08987426757813,
-20.3059272766113,
-17.5745258331299,
1.70560479164124,
18.5300540924072,
-9.87084007263184,
-27.8033180236816,
-2.80089426040649,
6.32665157318115,
1.89275300502777,
-12.7736158370972,
-0.695707380771637,
15.4606580734253,
-5.92179965972900,
-11.2869853973389,
1.37826132774353,
6.81527662277222,
-15.1228904724121,
-13.0226736068726,
-6.73495149612427,
10.7688970565796,
9.26662635803223,
-16.1759357452393,
-1.24422657489777,
4.12157249450684,
18.1742324829102,
-14.5250749588013,
-24.7015724182129,
-1.46034753322601,
-5.18207788467407,
-6.26757574081421,
2.19699835777283,
10.5942134857178,
-20.2243041992188,
-13.6318674087524,
-5.18548631668091,
-9.12209701538086,
-12.5133724212646,
-0.177153006196022,
-2.69819474220276,
-18.2158184051514,
5.08938169479370,
-13.7246532440186,
1.24289822578430,
-3.81823611259460,
-18.3351078033447,
11.7949142456055,
-16.0591106414795,
0.199888765811920,
9.90738677978516,
-9.53557491302490,
3.20832228660584,
11.3708477020264,
5.37669706344605,
-4.54445648193359,
11.4381761550903,
-11.6769256591797,
-6.88406085968018,
22.5655975341797,
7.60998487472534,
6.72288465499878,
7.29322242736816,
-0.0164565425366163,
5.48972511291504,
7.17919874191284,
7.21251201629639,
1.58182024955750,
5.72209692001343,
7.60086917877197,
-18.7158432006836,
-2.58281874656677,
-2.65363717079163,
-0.551289141178131,
-2.61411476135254,
-7.67522525787354,
27.7808341979980,
1.51619958877563,
-5.36351060867310,
3.09523010253906,
-18.4408874511719,
-13.1791877746582,
-0.309266090393066,
-4.18588161468506,
-13.3380899429321,
5.00647926330566,
15.7931070327759,
-5.76498365402222,
-15.4870862960815,
6.27600145339966,
-1.36817133426666,
-1.88209688663483,
-11.7726926803589,
-28.2167663574219,
18.7874011993408,
-8.90421772003174,
-9.37937355041504,
8.41074466705322,
-4.77177715301514,
16.8504886627197,
-26.1980743408203,
0.722024500370026,
11.7738342285156,
-22.1316509246826,
0.490725934505463,
-4.26020526885986,
3.85273408889771,
-9.22000026702881,
-2.28642177581787,
3.28997468948364,
-15.3389530181885,
11.5782289505005,
6.32829332351685,
-6.26223659515381,
6.58104085922241,
-5.76919698715210,
-22.3065567016602,
3.56587290763855,
7.09513998031616,
5.75518369674683,
5.66299104690552,
-4.13691139221191,
11.9876213073730,
11.3540706634521,
15.5025758743286,
-7.35353946685791,
-20.1289062500000,
5.35764789581299,
18.0263938903809,
-9.29254817962647,
-8.04965972900391,
13.0402793884277,
-9.79511737823486,
7.36063098907471,
-10.7468128204346,
-5.64769077301025,
25.8689136505127,
-23.7577095031738,
1.74611937999725,
35.0570869445801,
-1.59157419204712,
4.22511434555054,
3.26312899589539,
-0.550333142280579,
-0.889632403850555,
4.96493911743164,
4.44721126556397,
-15.1368112564087,
13.5265684127808,
4.23333406448364,
-0.597591817378998,
-9.87409019470215,
-7.21238899230957,
21.9043579101563,
-32.9478111267090,
0.770342886447907,
19.5426025390625,
-19.2725734710693,
18.0679779052734,
13.4841547012329,
5.26156044006348,
6.62342977523804,
7.64840030670166,
4.57341051101685,
-26.4238643646240,
1.68131005764008,
17.2562694549561,
-27.3179378509522,
-13.7374553680420,
19.1078128814697,
2.86223983764648,
-20.1318359375000,
1.07832336425781,
22.6050415039063,
7.84862375259399,
10.4965934753418,
1.72366642951965,
6.76770448684692,
-5.27587032318115,
-18.8037185668945,
23.4147853851318,
5.24941730499268,
-0.392378836870194,
1.08291506767273,
-2.77031517028809,
16.4326705932617,
12.6014060974121,
5.68207931518555,
-12.5043783187866,
17.7289810180664,
12.9805355072021,
-22.5480442047119,
3.72850346565247,
15.1375942230225,
-4.72188425064087,
-6.83578968048096,
-9.65443611145020,
-2.54548525810242,
12.3751640319824,
-12.2747344970703,
-5.44423151016235,
7.90767145156860,
-16.2349166870117,
-10.2553730010986,
17.5345554351807,
6.50615596771240,
5.37398624420166,
14.2051219940186,
-13.0191183090210,
-14.9490680694580,
-11.2286586761475,
2.29111433029175,
-10.6610507965088,
-21.0165843963623,
11.6086444854736,
-21.2882041931152,
-8.81852340698242,
11.5195646286011,
-15.3100175857544,
-27.5981369018555,
-6.13356304168701,
12.2465648651123,
-26.2298259735107,
7.05977344512939,
1.68790745735168,
-25.2254257202148,
0.422351062297821,
5.07650136947632,
19.2187614440918,
10.2367010116577,
1.74280500411987,
-2.43297624588013,
-2.82407140731812,
12.6382532119751,
6.26315784454346,
-8.00576877593994,
-11.1122169494629,
-21.8108749389648,
-1.83610558509827,
2.84729290008545,
-5.94244861602783,
0.313286989927292,
10.7461814880371,
13.9726963043213,
-23.3067741394043,
-9.55249881744385,
-7.50841283798218,
-27.0415306091309,
-12.1767206192017,
9.27261638641357,
14.8025512695313,
3.68879342079163,
21.4721126556397,
0.00878773443400860,
-17.7951335906982,
25.0400295257568,
4.90483951568604,
-12.8474292755127,
21.9064311981201,
-6.58537483215332,
-1.36534547805786,
12.3125505447388,
-10.0046596527100,
1.76027369499207,
-5.45851898193359,
-9.69639015197754,
1.46830141544342,
11.0461397171021,
3.66196656227112,
-16.2106971740723,
6.78599834442139,
32.2867774963379,
-20.5891933441162,
-3.90047049522400,
20.4575500488281,
-29.0730857849121,
7.26953315734863,
13.0421638488770,
-9.68792343139648,
-17.0856304168701,
2.73415422439575,
19.3890857696533,
-12.4184083938599,
11.7740240097046,
-0.422578454017639,
-17.9054985046387,
-0.228603139519691,
4.45863771438599,
20.7341594696045,
3.66194796562195,
-4.59748697280884,
10.5912666320801,
2.04863882064819,
-8.61873912811279,
2.82644534111023,
2.98038172721863,
10.6869182586670,
7.46327114105225,
-9.53777980804443,
24.3778076171875,
14.2008018493652,
9.27485656738281,
11.1849803924561,
-11.1362428665161,
6.82265520095825,
-1.17713403701782,
4.34631299972534,
-1.31473779678345,
-14.2701501846313,
7.90949201583862,
3.74013185501099,
-23.3175163269043,
-8.52509593963623,
19.7268657684326,
-5.77799844741821,
9.38212871551514,
10.3746519088745,
-13.1554718017578,
20.0349197387695,
10.8554639816284,
-10.0817909240723,
18.9033870697022,
19.8932781219482,
9.80140113830566,
1.14861059188843,
-18.8536720275879,
4.80715179443359,
-6.12957715988159,
3.33241724967957,
-1.83856594562531,
-9.54883384704590,
11.3255624771118,
-21.3600349426270,
15.8819141387939,
-12.0484704971313,
0.407144010066986,
31.6169433593750,
-26.3930625915527,
8.44781112670898,
19.3569564819336,
-2.09778380393982,
-18.5246791839600,
-4.78475761413574,
19.1997909545898,
8.82198429107666,
-19.6494617462158,
1.32610666751862,
27.7065715789795,
-21.0546150207520,
12.3493661880493,
5.77031564712524,
-17.9714603424072,
29.8108997344971,
14.1899738311768,
14.7949848175049,
-11.6059865951538,
-21.8965644836426,
19.9525394439697,
17.3010768890381,
-1.16669559478760,
-1.21370947360992,
7.01818752288818,
14.9051866531372,
8.38038444519043,
-11.9448852539063,
26.7323551177979,
-4.76768875122070,
-2.66491103172302,
35.5139884948731,
-15.5023031234741,
17.3921871185303,
-0.415739268064499,
-9.99899864196777,
0.487279474735260,
-5.87936973571777,
9.71126270294190,
-23.2516422271729,
12.6797428131104,
-11.1479921340942,
-10.6362962722778,
12.9947509765625,
-3.32704424858093,
23.3291797637939,
-8.98082542419434,
-7.54998540878296,
-14.8162431716919,
3.06398320198059,
-3.75566148757935,
-20.9689044952393,
16.9260768890381,
-11.1967916488647,
11.7803993225098,
0.821936905384064,
-6.26036119461060,
2.20901036262512,
-6.76704883575439,
15.2503337860107,
0.205194160342217,
8.70254898071289,
-11.9431295394897,
11.2089319229126,
16.7095298767090,
-23.9663543701172,
-8.43136978149414,
-7.32973861694336,
2.40240001678467,
4.71879959106445,
13.1459178924561,
2.97896766662598,
-11.8125000000000,
5.31741380691528,
4.00719785690308,
-10.9401550292969,
5.81751012802124,
7.71904659271240,
-24.7084217071533,
16.9854412078857,
4.22706460952759,
-19.1337776184082,
21.5945625305176,
3.77084589004517,
9.94618988037109,
11.1384973526001,
9.34064388275147,
16.6932353973389,
-3.72208023071289,
5.30608081817627,
15.1547651290894,
-2.56938576698303,
1.57817745208740,
3.98283457756043,
-13.2195024490356,
4.78111505508423,
-2.53686809539795,
-21.4017028808594,
-19.7498188018799,
8.20913696289063,
15.1546039581299,
-16.5295829772949,
-6.05288267135620,
-4.53664255142212,
2.58062338829041,
0.615664601325989,
-16.1543922424316,
-12.1717872619629,
-9.10280513763428,
-5.45895242691040,
-13.0578699111938,
2.34008455276489,
8.87492942810059,
-16.5014705657959,
-12.5736265182495,
9.98999023437500,
-10.2163791656494,
-22.9951534271240,
9.31542110443115,
12.6188669204712,
2.12090182304382,
0.686182796955109,
-3.28388714790344,
-17.8817825317383,
-0.151315674185753,
12.9186048507690,
-13.8678989410400,
2.38793635368347,
3.93875384330750,
2.59122633934021,
-5.11967992782593,
2.24098920822144,
30.0208778381348,
-8.27184581756592,
-10.4395132064819,
-9.91821193695068,
-13.5447101593018,
-6.21152448654175,
-8.26899814605713,
-7.43961811065674,
-17.3414955139160,
1.02944922447205,
-0.929444074630737,
-0.663496732711792,
-10.1054325103760,
16.2734718322754,
-0.688442468643189,
-19.5476074218750,
15.3724832534790,
-12.4625015258789,
2.27023148536682,
-1.44227325916290,
12.0383138656616,
4.55966186523438,
5.03598880767822,
3.51187849044800,
-7.86672830581665,
12.6866912841797,
-23.3472080230713,
-17.3497562408447,
-2.18137264251709,
14.3884057998657,
-19.9131603240967,
-2.58917021751404,
30.4288578033447,
-4.72489404678345,
-16.5985946655273,
6.71154785156250,
25.1118907928467,
7.89771366119385,
16.3774356842041,
-11.0279369354248,
-9.51023197174072,
-5.99009084701538,
-19.0481643676758,
-11.9262084960938,
-8.78918075561523,
-23.7985324859619,
-9.57968616485596,
9.49487781524658,
0.595957040786743,
18.0634307861328,
-2.67861771583557,
-19.0716190338135,
-14.6505270004272,
12.3889846801758,
7.12666273117065,
-5.64854717254639,
-9.25631427764893,
-18.9157714843750,
-14.3497810363770,
-8.11893367767334,
5.06933546066284,
-15.7915573120117,
6.26205825805664,
11.3642253875732,
1.74126470088959,
-2.87640094757080,
-2.30282425880432,
3.92401862144470,
-20.4661006927490,
6.68468093872070,
7.47779464721680,
5.70047378540039,
-8.93116569519043,
-18.9331855773926,
-7.46915245056152,
-27.3449916839600,
15.5949449539185,
-0.840401828289032,
-7.63225984573364,
23.5428962707520,
6.01335525512695,
6.91772985458374,
-7.97308015823364,
-2.35811305046082,
-12.1857099533081,
-6.93674707412720,
-10.1884899139404,
-16.2725410461426,
11.0032243728638,
-14.6339302062988,
-12.6519546508789,
-5.75399017333984,
5.58025455474854,
13.7735252380371,
-25.1665019989014,
1.15240776538849,
20.1981124877930,
-20.9958992004395,
7.62956476211548,
24.0972480773926,
-12.3138542175293,
-9.19274806976318,
-10.4318161010742,
4.29953193664551,
4.66203546524048,
-21.6051464080811,
-8.61791515350342,
-12.8580360412598,
-22.9328994750977,
-17.0765933990479,
-6.16697788238525,
-0.291236698627472,
-17.0545425415039,
-23.7027664184570,
0.805502414703369,
0.712448000907898,
-25.1160125732422,
-3.27644014358521,
12.8621520996094,
-5.14219903945923,
-11.5089559555054,
-6.29354763031006,
-9.55434131622315,
5.80042219161987,
12.3375492095947,
-2.78816080093384,
3.90938854217529,
-6.45162487030029,
-10.4027347564697,
11.0849590301514,
23.4066753387451,
-13.7208147048950,
-7.50126171112061,
13.9823722839355,
-26.6295509338379,
0.0118719376623631,
12.3976516723633,
0.604991614818573,
13.3346815109253,
-10.3703107833862,
11.6211299896240,
12.0819034576416,
-21.2845134735107,
10.2225799560547,
0.122850075364113,
-18.0094795227051,
13.1090030670166,
15.1221704483032,
1.28883755207062,
19.1642303466797,
20.3114719390869,
-16.2592239379883,
6.86915159225464,
12.6652450561523,
-6.03191089630127,
0.984592497348785,
-0.436796933412552,
-5.54803991317749,
-18.3003292083740,
12.6446304321289,
-5.00582981109619,
-26.0187149047852,
18.8699493408203,
4.47473955154419,
-8.40136337280273,
13.3080034255981,
-8.84838867187500,
-5.28630304336548,
15.6431255340576,
-14.5917854309082,
5.03715467453003,
20.2728805541992,
7.28868722915649,
14.6491451263428,
-11.3841180801392,
11.4545526504517,
10.7538862228394,
-6.45581340789795,
10.9844818115234,
-21.1238117218018,
-4.67120790481567,
12.2825174331665,
8.17920112609863,
14.4360780715942,
-2.13354682922363,
10.5758171081543,
15.7033414840698,
5.93398523330689,
0.428269088268280,
5.67986583709717,
20.8419799804688,
-17.3216686248779,
-10.0161399841309,
27.8469066619873,
-4.32356119155884,
-7.13166952133179,
9.78790664672852,
0.181835263967514,
-17.7271404266357,
3.09456443786621,
4.14605903625488,
-12.5471067428589,
-2.62518048286438,
-15.8638019561768,
13.3968667984009,
-4.12830066680908,
-15.5378313064575,
18.2557411193848,
-19.0732898712158,
9.39669704437256,
6.84419536590576,
-23.0888175964355,
17.2972278594971,
8.51423263549805,
-3.83320546150208,
10.0425453186035,
17.5337715148926,
1.49036490917206,
-9.77091693878174,
-14.3756237030029,
7.48609352111816,
21.8138713836670,
-18.4317417144775,
-11.7038316726685,
12.9244174957275,
1.58917582035065,
-23.0362777709961,
-3.30844354629517,
24.3000164031982,
-14.5982961654663,
-8.72235965728760,
4.88705682754517,
-15.8765382766724,
2.18824720382690,
-3.50562191009522,
2.63917326927185,
3.01189637184143,
-19.7280139923096,
-5.57341909408569,
10.8089723587036,
18.1312103271484,
-6.47507143020630,
-1.59479808807373,
16.4681491851807,
9.76740837097168,
1.86185908317566,
3.55731201171875,
21.7072353363037,
-3.19356966018677,
-19.7623291015625,
-10.5461444854736,
-2.94166660308838,
-2.67476773262024,
-7.67240333557129,
-19.0804767608643,
-6.75547409057617,
24.6149120330811,
4.75951814651489,
2.22785878181458,
2.30173993110657,
8.17122650146484,
8.45393466949463,
-8.92030429840088,
12.6420478820801,
0.0481488481163979,
7.69426298141480,
11.5407400131226,
-13.0177593231201,
-3.85568404197693,
-14.4619913101196,
-0.605136096477509,
-12.1739511489868,
-22.4092922210693,
0.639689147472382,
-9.10286808013916,
14.2112083435059,
-0.317572236061096,
-9.19659423828125,
-0.342797309160233,
-5.62212944030762,
7.57282400131226,
7.82754468917847,
20.9320011138916,
-12.1267251968384,
-14.8363876342773,
-2.95752358436584,
2.69033193588257,
14.1886568069458,
-19.1055355072022,
1.05314385890961,
-10.5712366104126,
-16.6796646118164,
16.3043136596680,
-17.8936328887939,
-22.1390495300293,
-0.904880583286285,
2.43419957160950,
-8.49969768524170,
-12.1067142486572,
16.3642978668213,
-3.04696416854858,
-5.70817613601685,
3.46039724349976,
2.63047170639038,
17.7135028839111,
-10.4153957366943,
-12.7926921844482,
-2.34385657310486,
9.08910655975342,
1.85355734825134,
6.41322803497314,
12.9283561706543,
-16.1506557464600,
11.4810914993286,
10.9482746124268,
-1.22785770893097,
-10.6644372940063,
-14.0955057144165,
15.4870500564575,
-9.25712585449219,
-23.6418857574463,
5.23377799987793,
-2.28203439712524,
-21.0809936523438,
7.71437931060791,
4.25784301757813,
-3.36674904823303,
-4.48478460311890,
-5.96879816055298,
25.2825698852539,
-9.86691665649414,
-3.71124505996704,
1.12747168540955,
-9.10206508636475,
21.2877712249756,
-11.6839408874512,
-16.9589538574219,
-5.99812507629395,
-11.3883314132690,
-15.3718032836914,
4.67730379104614,
-4.79152679443359,
-30.0902042388916,
-1.11928105354309,
7.26376295089722,
-8.05583667755127,
-17.1129016876221,
-3.90728497505188,
-5.61754465103149,
9.64875793457031,
8.31916332244873,
-12.4465599060059,
0.768177211284638,
4.92934703826904,
14.5390529632568,
5.50990724563599,
-2.87898564338684,
-7.77198314666748,
-9.38867378234863,
-1.98297858238220,
-6.11989879608154,
-10.4792861938477,
-12.0617504119873,
5.73629570007324,
-8.17419052124023,
-2.51889801025391,
23.1050872802734,
5.06989336013794,
14.5107498168945,
3.41523647308350,
-0.956790387630463,
4.88806867599487,
-5.61723089218140,
12.0617618560791,
-6.26734542846680,
-14.1180143356323,
2.52668190002441,
4.09251070022583,
3.06036567687988,
-4.90361022949219,
-11.9872941970825,
-3.96246027946472,
17.3523101806641,
-5.35351133346558,
-19.5919628143311,
11.5556077957153,
7.30318975448608,
-9.91288471221924,
4.39867448806763,
19.2249851226807,
3.89409589767456,
0.510644733905792,
-12.3651027679443,
-15.7878808975220,
16.1803894042969,
-8.28972911834717,
-20.9632606506348,
-13.4434633255005,
-1.05028259754181,
9.23397636413574,
-1.74346768856049,
10.0953092575073,
-12.1180095672607,
0.922256350517273,
12.4483118057251,
-13.8263072967529,
0.192329704761505,
-4.86940050125122,
-0.202733233571053,
5.02822971343994,
0.202239185571671,
-3.10148334503174,
-0.401490688323975,
11.5679683685303,
9.49289417266846,
11.9909925460815,
-0.856192052364349,
3.57382822036743,
1.29161369800568,
-11.0209560394287,
-7.34124898910523,
-7.96214532852173,
-15.7320632934570,
-19.3930664062500,
-5.17983722686768,
-13.1234016418457,
-11.5021743774414,
-6.24388647079468,
-3.63600707054138,
1.90180206298828,
10.2053756713867,
-7.64657402038574,
-14.9665222167969,
13.6600179672241,
-23.8254013061523,
-12.2153854370117,
18.2992477416992,
5.57329273223877,
13.1281614303589,
2.78803682327271,
16.5992927551270,
7.98059415817261,
1.85574090480804,
8.70498847961426,
4.90680456161499,
11.3484201431274,
6.81137657165527,
16.3201274871826,
6.36159133911133,
16.1707153320313,
6.02147340774536,
-11.5794315338135,
2.32117176055908,
12.2287149429321,
1.45446956157684,
-21.7409343719482,
-4.58901691436768,
-1.82590782642365,
11.0599975585938,
15.7256908416748,
4.58339071273804,
7.62615633010864,
5.00244903564453,
8.22729301452637,
8.39834785461426,
2.62158107757568,
3.54248571395874,
0.0344786494970322,
-5.81449317932129,
11.1045475006104,
-0.949545085430145,
7.79178142547607,
19.9700107574463,
-17.1695728302002,
0.709490001201630,
19.0141487121582,
-2.97510242462158,
-15.6964902877808,
13.7153730392456,
17.2235870361328,
-5.69332599639893,
7.83623027801514,
-8.96452808380127,
8.16429138183594,
9.32745838165283,
2.90535712242126,
11.0286788940430,
-5.39339447021484,
16.4089584350586,
18.9783649444580,
13.6696987152100,
12.3807258605957,
-4.12063837051392,
-9.98159694671631,
13.8171825408936,
1.41499829292297,
-15.2153701782227,
23.8286533355713,
0.903553962707520,
-20.6488876342773,
-0.303845882415772,
-6.51534891128540,
1.61201560497284,
-0.652941405773163,
1.74439084529877,
6.27643203735352,
-7.46903657913208,
8.37570095062256,
15.0747900009155,
5.33746194839478,
17.7982482910156,
18.8390998840332,
5.79728794097900,
3.77450871467590,
22.8762626647949,
13.1544132232666,
-14.6317977905273,
-0.641010761260986,
-8.97636222839356,
4.64830923080444,
-2.45757699012756,
-7.28193521499634,
17.7556781768799,
-19.4404926300049,
-0.355495333671570,
8.57216835021973,
-19.8346042633057,
0.731327414512634,
8.06882286071777,
-11.5384922027588,
-2.67364263534546,
2.83626651763916,
-0.659088253974915,
7.71721172332764,
-19.8311100006104,
-14.5947017669678,
-9.79516983032227,
-1.88936030864716,
16.0552062988281,
-3.08292508125305,
7.59930038452148,
3.80944514274597,
-4.47670793533325,
-6.92144727706909,
12.2127075195313,
16.8558349609375,
-8.98393821716309,
-0.700205683708191,
5.23426675796509,
22.2606105804443,
-1.80371582508087,
4.40772676467896,
20.7376003265381,
-5.22892236709595,
-0.839825630187988,
-8.64877414703369,
8.97337055206299,
-15.8656215667725,
-24.5617885589600,
-0.227282077074051,
-15.9652948379517,
0.167177006602287,
-5.09936189651489,
3.01451396942139,
4.19146299362183,
-23.7797927856445,
-10.9818868637085,
13.8099021911621,
15.4937934875488,
-0.404192388057709,
-3.75425624847412,
-9.07670879364014,
-12.7180490493774,
-13.1377515792847,
14.9231166839600,
7.90318441390991,
-26.3806190490723,
3.02838611602783,
6.97959852218628,
-11.5731267929077,
10.9211587905884,
17.3814315795898,
-19.0544815063477,
-2.32520842552185,
16.5750293731689,
13.5819807052612,
-1.78421366214752,
-9.53003406524658,
23.9804267883301,
-8.46333312988281,
-7.00533151626587,
18.2143573760986,
6.35451364517212,
-13.2317190170288,
-9.35569286346436,
15.9851055145264,
-9.72864246368408,
11.0680189132690,
6.24083518981934,
-12.7948284149170,
10.7872123718262,
-18.4889411926270,
-13.8796806335449,
-0.491295218467712,
-0.444772511720657,
13.1109943389893,
1.64874291419983,
2.94930958747864,
-1.40964674949646,
-12.5836849212646,
5.62523794174194,
17.7731800079346,
-11.5775566101074,
-16.4894638061523,
-5.65605926513672,
-7.65528631210327,
1.81118190288544,
-13.5355825424194,
9.41816806793213,
-2.21744251251221,
-19.0749683380127,
5.44875097274780,
-16.5011596679688,
7.29159402847290,
17.6310539245605,
-8.88725757598877,
-12.4405279159546,
1.66037273406982,
-9.68629837036133,
-19.3625831604004,
-7.22192096710205,
-3.22901844978333,
1.49382960796356,
-20.7516384124756,
-16.4027290344238,
-0.709451019763947,
11.4377927780151,
-3.91979622840881,
-18.7056617736816,
-6.67455816268921,
-0.981695055961609,
-1.10486185550690,
-14.7443256378174,
-12.9167003631592,
-15.6942939758301,
-2.69350337982178,
-12.3044176101685,
-20.9963226318359,
-10.6058864593506,
-5.53928232192993,
9.71222591400147,
-19.8411769866943,
-14.9120750427246,
18.4812831878662,
3.52769446372986,
-2.49162960052490,
18.0868453979492,
0.743387281894684,
-23.1056385040283,
13.6667757034302,
3.00738954544067,
-1.49350500106812,
20.6799106597900,
-7.28783464431763,
0.387540668249130,
-2.78921127319336,
8.30669021606445,
1.01124513149261,
-22.4413547515869,
18.9712352752686,
-1.28526437282562,
2.48211669921875,
4.21412897109985,
-9.60992431640625,
23.6496047973633,
5.00721168518066,
11.6145582199097,
-6.55911731719971,
-10.2970151901245,
10.6360788345337,
-14.3290243148804,
12.0387096405029,
-0.825835347175598,
-1.13271224498749,
11.8865289688110,
-13.4247989654541,
10.0042295455933,
-5.28933429718018,
-19.0982303619385,
9.12661361694336,
7.34008789062500,
-9.72071647644043,
-13.0790157318115,
7.89372301101685,
9.35078525543213,
-25.8736553192139,
-3.35641551017761,
14.1677665710449,
-8.89997959136963,
16.1121139526367,
14.3322916030884,
12.9716424942017,
-7.72159910202026,
-22.6601505279541,
-0.743004262447357,
-7.94886589050293,
7.17208909988403,
-19.5952148437500,
-6.56053543090820,
10.9295301437378,
-14.0613260269165,
16.6109733581543,
-8.93202877044678,
2.93154358863831,
2.20515036582947,
-20.7077026367188,
29.4698677062988,
-1.56651902198792,
-11.6715335845947,
14.4589929580688,
0.184026882052422,
1.79498851299286,
1.46902740001678,
4.44161891937256,
12.2187643051147,
-9.85692596435547,
-0.520260930061340,
27.8285369873047,
-8.86148738861084,
1.24048769474030,
20.7704696655273,
-9.95589637756348,
-5.21493959426880,
12.6539335250855,
16.1803188323975,
-10.3659744262695,
-3.22691226005554,
18.3458671569824,
5.06617259979248,
4.18219947814941,
-5.82314062118530,
11.4214820861816,
5.34931325912476,
-11.0002737045288,
7.81972646713257,
3.25852346420288,
-0.0717168152332306,
-6.43564128875732,
14.0793809890747,
4.00394344329834,
-19.1351928710938,
-6.76701593399048,
-7.58455705642700,
-8.86865806579590,
-17.8887844085693,
17.0420837402344,
14.4167480468750,
-23.3169803619385,
12.0406970977783,
7.64596271514893,
-4.55520296096802,
17.9487400054932,
7.88315439224243,
3.60641789436340,
15.0057935714722,
19.2641754150391,
3.31177949905396,
-17.4133052825928,
13.2488193511963,
19.4273834228516,
-11.8545274734497,
19.1343650817871,
8.21587848663330,
-25.8637256622314,
-7.68225669860840,
10.6193161010742,
11.9600324630737,
-11.5394535064697,
-0.224830240011215,
8.14162445068359,
-11.2417449951172,
6.40939331054688,
13.6871767044067,
-7.86548423767090,
5.89770269393921,
6.80252218246460,
-12.9602031707764,
-1.98341155052185,
-4.30429697036743,
-7.19855642318726,
-2.17773342132568,
-7.29447603225708,
-17.4751071929932,
-8.22329139709473,
1.23664283752441,
-0.221830055117607,
2.07733750343323,
16.6320915222168,
11.4607791900635,
-19.7313461303711,
17.8324184417725,
20.5639057159424,
-22.9599399566650,
2.84511041641235,
8.97846889495850,
-31.4084949493408,
0.647261500358582,
9.78771209716797,
-10.5013084411621,
7.58908605575562,
-9.13439273834229,
9.32405281066895,
-9.04821872711182,
-6.31478357315064,
21.0596160888672,
0.351409435272217,
-0.541563749313355,
0.196944743394852,
2.09245252609253,
4.32163667678833,
17.9228057861328,
5.79862833023071,
0.862236857414246,
-2.99491429328918,
6.74960422515869,
11.8521718978882,
-0.702143251895905,
-3.07158994674683,
-18.0974369049072,
-2.16524577140808,
-0.259203106164932,
-4.25065374374390,
12.4108886718750,
-4.90072584152222,
-23.0492725372314,
10.0857229232788,
2.75925254821777,
-7.36768054962158,
24.8423805236816,
-8.65603065490723,
-13.7357196807861,
18.8264484405518,
11.8029441833496,
-13.1622352600098,
-18.0406322479248,
20.2556571960449,
-5.29510068893433,
-29.4934120178223,
15.3076486587524,
17.4274845123291,
-1.05946624279022,
-8.29071331024170,
-0.617962896823883,
-1.30753886699677,
3.29659271240234,
9.33983230590820,
-15.7959690093994,
0.507034659385681,
21.2358055114746,
-3.80885195732117,
-23.2101573944092,
1.61212694644928,
-10.2145957946777,
-18.2709121704102,
-7.46959066390991,
-16.8813381195068,
15.5465517044067,
-5.98434305191040,
-6.93521833419800,
0.507627010345459,
-17.0239582061768,
-12.2448701858521,
-10.4415569305420,
15.3190832138062,
1.87759816646576,
-15.9976167678833,
-14.0502233505249,
-2.86761212348938,
0.910829067230225,
1.15739548206329,
-3.09154558181763,
-2.17359519004822,
0.332403898239136,
-14.5623826980591,
-7.86223173141480,
4.28470182418823,
13.2054290771484,
-19.6181735992432,
-16.8561573028564,
10.6949911117554,
-10.3770704269409,
-20.7753696441650,
-7.49628353118897,
14.4055490493774,
8.61825466156006,
2.34847950935364,
-4.98656463623047,
-11.3695907592773,
8.02951049804688,
-10.8248195648193,
-18.1265888214111,
-1.87136459350586,
-19.6455764770508,
-8.68391323089600,
1.54012608528137,
0.655984342098236,
-3.83717727661133,
0.143440783023834,
7.59712982177734,
3.14324212074280,
18.4727725982666,
1.09445536136627,
5.75834083557129,
-4.90165567398071,
-12.8829040527344,
8.57565975189209,
3.39688491821289,
3.27302384376526,
-18.6383666992188,
7.62223768234253,
17.7271003723145,
-0.367471486330032,
14.0195083618164,
3.75198340415955,
0.205891534686089,
1.67524266242981,
-6.68741607666016,
-8.72920703887940,
7.59481620788574,
-9.78679275512695,
-16.6140651702881,
-8.96617317199707,
-10.6216812133789,
4.66158771514893,
-15.3628473281860,
5.58642959594727,
-1.77058792114258,
-18.3932285308838,
13.7278909683228,
8.48489379882813,
6.66046571731567,
-11.2427444458008,
-0.473893195390701,
-6.76704406738281,
1.67577791213989,
17.5888652801514,
-11.1014404296875,
7.82623338699341,
-5.58982419967651,
2.31770277023315,
4.73085689544678,
-6.15819835662842,
13.1390876770020,
-12.1804504394531,
-2.95149731636047,
10.5924301147461,
7.03922510147095,
5.17536020278931,
-9.35284328460693,
2.71027708053589,
5.45197057723999,
1.45780003070831,
16.9573974609375,
10.9995059967041,
-7.71636056900024,
-0.794032454490662,
-5.31668615341187,
-13.5974254608154,
1.67292475700378,
10.6811552047730,
3.69029974937439,
-8.96002006530762,
-10.9477834701538,
-8.51286983489990,
-5.12216377258301,
5.27182197570801,
3.09102439880371,
-12.9442434310913,
-7.45967197418213,
-0.515651583671570,
7.91900014877319,
8.11241054534912,
9.38945388793945,
12.1929531097412,
-11.1450977325439,
7.46659183502197,
22.4585533142090,
-9.04221248626709,
-13.0587129592896,
-1.84222316741943,
-7.60892295837402,
-9.10823631286621,
-19.1654529571533,
-1.78305113315582,
-3.39981913566589,
-9.04961490631104,
12.8564214706421,
-10.0262603759766,
12.9830665588379,
2.60228419303894,
-11.0787038803101,
15.4212656021118,
-9.78343009948731,
-12.1092548370361,
-15.1309309005737,
-2.48928427696228,
12.5813474655151,
5.83123302459717,
-8.36228275299072,
-10.3986940383911,
17.7862281799316,
-7.67706489562988,
-10.3834476470947,
14.6162719726563,
13.1139640808105,
5.46555852890015,
0.809445083141327,
4.67825365066528,
-12.1199159622192,
10.1363935470581,
9.49260902404785,
-0.660555183887482,
-0.924318850040436,
-0.709350705146790,
26.0604400634766,
-19.3077907562256,
0.822396993637085,
16.3352603912354,
-16.0572147369385,
15.6166267395020,
-5.82133913040161,
10.2777042388916,
26.2325019836426,
-15.8405237197876,
-9.53750133514404,
0.140627503395081,
-8.02367877960205,
7.09079599380493,
-10.0664482116699,
-14.7435083389282,
15.0051345825195,
-15.6261043548584,
-14.1577081680298,
-5.34226226806641,
7.59853601455689,
5.74792861938477,
-7.70336580276489,
24.1729297637939,
-2.52697801589966,
-13.2236175537109,
-5.76699972152710,
16.5256633758545,
3.93221044540405,
-24.0902194976807,
5.17597579956055,
-7.41697359085083,
10.9587602615356,
-9.82494640350342,
-6.73653650283814,
10.7049016952515,
-16.2900066375732,
17.1203632354736,
3.32602763175964,
-13.2541618347168,
-7.09393453598023,
9.34467506408691,
-5.96971940994263,
3.78957056999207,
8.92294597625732,
-7.28977584838867,
11.6284427642822,
-15.2671985626221,
19.1477222442627,
5.83985853195190,
-9.10669422149658,
6.90311479568481,
-3.89340615272522,
19.7111129760742,
-12.3581867218018,
1.31073653697968,
2.70050048828125,
-8.49369430541992,
16.1767215728760,
4.26552772521973,
-7.31008195877075,
-11.2396221160889,
-4.84684848785400,
-10.9897499084473,
14.4600162506104,
-4.04187631607056,
-6.40831708908081,
2.50282621383667,
-17.5950336456299,
5.69347429275513,
-11.7576026916504,
7.36147451400757,
13.1633939743042,
5.29633712768555,
-8.58045482635498,
-17.8714752197266,
1.55384480953217,
-13.4814376831055,
-3.14614844322205,
1.82144498825073,
1.88360202312469,
15.0700082778931,
9.20624160766602,
-6.29249095916748,
4.29661893844605,
-2.09479427337647,
-2.59619235992432,
10.7207851409912,
7.75627231597900,
14.5713348388672,
-15.3646993637085,
-7.46383333206177,
11.4402399063110,
-3.99211955070496,
16.1805553436279,
-7.12983131408691,
-14.9017410278320,
11.8812494277954,
-2.42547535896301,
-7.11111164093018,
-4.35227966308594,
11.2642250061035,
2.99096941947937,
-15.9365406036377,
7.41449832916260,
12.1566257476807,
-13.7486438751221,
-19.9542713165283,
6.93306446075439,
8.98659229278565,
-16.9407958984375,
8.66964149475098,
13.1153602600098,
-5.76974582672119,
5.48646974563599,
2.95691275596619,
15.0732927322388,
5.13567304611206,
4.53397417068481,
21.6384468078613,
5.58016109466553,
6.75671577453613,
4.47856044769287,
0.867714464664459,
7.36150264739990,
1.67710077762604,
-0.534055292606354,
2.02176547050476,
10.4380750656128,
-2.98575997352600,
-13.7627782821655,
15.8472614288330,
2.90397119522095,
-11.1273803710938,
5.66678953170776,
-15.2742624282837,
-1.36971354484558,
3.70828127861023,
2.57881951332092,
14.4415769577026,
-13.8910989761353,
0.811905980110169,
-9.83253383636475,
-1.02921509742737,
22.9530639648438,
-1.54686260223389,
12.0476360321045,
18.0840854644775,
4.50934553146362,
-5.57636737823486,
-0.194103986024857,
-9.94289684295654,
-6.14552259445190,
-6.55744123458862,
-14.5034389495850,
5.98371219635010,
-17.3547973632813,
-4.16895961761475,
15.9999752044678,
-11.1747922897339,
-5.10293102264404,
7.21103572845459,
5.53039932250977,
-2.65661334991455,
5.27058410644531,
8.46320629119873,
7.14212274551392,
0.886299312114716,
-14.2955951690674,
19.1024360656738,
3.67325139045715,
-22.0520095825195,
-6.41860103607178,
-9.28315639495850,
17.1225395202637,
-9.60204601287842,
-3.82313942909241,
19.5305671691895,
-25.2863121032715,
-9.72267246246338,
-4.58997106552124,
-11.7188262939453,
2.76228070259094,
13.3058376312256,
14.5326271057129,
-5.84730148315430,
-14.7656822204590,
-2.34135723114014,
7.94518661499023,
1.32360184192657,
2.80753874778748,
13.4967641830444,
10.3378343582153,
-16.7956027984619,
-4.05010938644409,
7.94688987731934,
-18.7400627136230,
-5.80440616607666,
-1.82379710674286,
-1.02290761470795,
0.924795687198639,
-6.63642406463623,
-15.8995189666748,
-8.56108951568604,
16.6026287078857,
-7.17978143692017,
-10.3467035293579,
-8.68994998931885,
-9.88752651214600,
4.18537807464600,
6.69096326828003,
2.69274258613586,
-18.3759288787842,
1.18928742408752,
15.7287616729736,
-7.19875955581665,
-2.05441784858704,
19.3694190979004,
-11.9823160171509,
-14.3442316055298,
12.3505401611328,
-14.3068370819092,
-10.6618719100952,
3.95377135276794,
-3.87812328338623,
-5.99961757659912,
14.4777278900146,
-0.353492408990860,
-19.3453140258789,
18.5092048645020,
1.86974251270294,
-6.89899969100952,
13.6047306060791,
2.05548381805420,
9.26614093780518,
2.69299411773682,
-9.63071441650391,
5.96953010559082,
15.2265367507935,
0.201623007655144,
-5.45465230941773,
-9.99402332305908,
3.11412525177002,
15.2315778732300,
-11.4220504760742,
10.8558816909790,
-5.92987346649170,
-15.8504323959351,
16.0280475616455,
-15.1325683593750,
3.87662100791931,
5.02519273757935,
-17.8863754272461,
11.9395771026611,
13.0629396438599,
-11.5049343109131,
-10.5742101669312,
-3.66894698143005,
0.461259931325913,
1.16137731075287,
-14.3324251174927,
12.1254644393921,
-1.91362762451172,
-10.7836074829102,
11.3750514984131,
-14.1814689636230,
-2.77769207954407,
-3.46967959403992,
4.02062463760376,
4.99368762969971,
-3.50054764747620,
0.614945352077484,
-15.1535778045654,
8.33222103118897,
14.5356636047363,
10.8612632751465,
4.52332639694214,
15.6529750823975,
8.74356460571289,
-13.0559539794922,
10.8601751327515,
2.55738067626953,
0.470121234655380,
-9.33493137359619,
4.38992357254028,
-3.20727944374084,
-14.6111297607422,
9.77425289154053,
-10.9697589874268,
-7.14014291763306,
-15.3321208953857,
-10.0770568847656,
11.5170335769653,
3.04981780052185,
-4.00864791870117,
-9.48377990722656,
-2.89324831962585,
18.4693622589111,
-3.03715610504150,
-4.84196329116821,
4.93816852569580,
-13.9725418090820,
13.7580718994141,
4.47402906417847,
3.60125803947449,
-4.85378789901733,
-23.4929714202881,
2.31351304054260,
-3.61944794654846,
-7.42050933837891,
9.71635532379150,
-7.25256681442261,
2.98348426818848,
10.9829721450806,
-11.9451847076416,
17.9975414276123,
-2.67916798591614,
-5.30362272262573,
8.94321918487549,
0.543842256069183,
8.66543006896973,
4.16712999343872,
13.2015895843506,
15.5082654953003,
4.15647602081299,
-2.17504072189331,
18.5953712463379,
-2.79161286354065,
2.51570296287537,
13.1219253540039,
-15.0004777908325,
-7.64564037322998,
-1.42359483242035,
2.86298203468323,
-10.8691673278809,
-10.4292793273926,
1.53230607509613,
5.76888942718506,
-1.10931265354157,
-4.77508354187012,
13.6258792877197,
4.92127752304077,
-5.19352912902832,
3.82182788848877,
8.02687358856201,
-2.49075794219971,
8.01173973083496,
4.17607593536377,
-8.54513072967529,
17.3651313781738,
0.478731423616409,
-13.8486385345459,
7.98186540603638,
14.3295030593872,
7.83969259262085,
-3.45025444030762,
6.33023405075073,
9.12532806396484,
-12.1088790893555,
-13.4548063278198,
-0.963169634342194,
-8.47940731048584,
1.40927875041962,
-1.31056988239288,
-14.8375549316406,
-0.389630317687988,
-6.74552679061890,
-2.72836542129517,
-6.17471599578857,
-12.1885938644409,
-1.23666691780090,
-12.4713315963745,
-4.81382417678833,
-5.85101079940796,
-3.95315647125244,
25.1233196258545,
-3.70604634284973,
-15.4220151901245,
14.5771131515503,
-1.11586070060730,
6.25171470642090,
2.42524361610413,
-15.2397670745850,
-9.29746627807617,
-16.6033382415772,
-5.41436910629273,
-13.9162082672119,
9.58430290222168,
2.35130381584168,
-13.6959867477417,
12.8839941024780,
-14.6714496612549,
12.6420087814331,
1.96156811714172,
-11.5898208618164,
22.2410907745361,
1.55988764762878,
5.90199804306030,
6.30316257476807,
9.04469203948975,
14.8873386383057,
2.29529786109924,
11.1565885543823,
11.2281332015991,
-3.71333742141724,
9.44561958312988,
15.0544910430908,
14.4698371887207,
0.897774338722229,
-9.90147781372070,
12.2980451583862,
7.09771442413330,
3.65569615364075,
-0.664995491504669,
-2.00504159927368,
12.3877267837524,
16.8758029937744,
-0.490803748369217,
-14.1288385391235,
-9.34495067596436,
-4.10147666931152,
11.4437980651855,
11.4496889114380,
-4.22844982147217,
-10.5161523818970,
7.99212789535523,
-1.02602052688599,
-13.4813890457153,
2.06742477416992,
-2.24335265159607,
2.83121633529663,
0.528813898563385,
-6.79536771774292,
-6.84109830856323,
4.26928997039795,
11.1444053649902,
-13.4602136611938,
-2.82553434371948,
9.80541324615479,
2.12311244010925,
-10.2036943435669,
-3.00853133201599,
5.82699775695801,
-16.2097434997559,
2.15648770332336,
19.0636558532715,
11.5756168365479,
-15.0561580657959,
-17.8889904022217,
1.72046756744385,
2.18963241577148,
18.9787788391113,
4.84666109085083,
-9.10584449768066,
-8.25858974456787,
0.826050639152527,
0.223563149571419,
-14.9188871383667,
10.1137161254883,
-10.4018640518188,
-18.0348434448242,
5.92243576049805,
-17.1140899658203,
-5.84712648391724,
-0.942220032215118,
-21.7300796508789,
-9.72916412353516,
-9.13018798828125,
-12.7930116653442,
2.96726059913635,
-3.48539566993713,
-8.28897380828857,
4.43920183181763,
1.99930357933044,
-9.38851547241211,
-7.29972553253174,
1.03865134716034,
3.42684412002563,
9.96374893188477,
-1.47156858444214,
-10.3291873931885,
9.53190135955811,
-0.257713496685028,
-16.2209720611572,
-4.73377323150635,
-5.56888484954834,
17.4525585174561,
3.07293701171875,
-16.4504966735840,
20.9201602935791,
8.17917823791504,
7.57022190093994,
5.67499208450317,
-9.73682785034180,
1.37104451656342,
-2.65865564346313,
-10.3303470611572,
-5.58706760406494,
-4.75008344650269,
-18.4282684326172,
-14.9405097961426,
4.74811124801636,
9.76279830932617,
-6.73740959167481,
-5.24950981140137,
9.43089294433594,
18.8296184539795,
0.618167757987976,
0.226276174187660,
11.0683164596558,
-13.0304632186890,
9.50494480133057,
13.7656354904175,
3.05149841308594,
-7.54927349090576,
-1.74822509288788,
29.2552719116211,
-9.77996730804443,
-4.60092401504517,
0.521298944950104,
-16.8471946716309,
3.81053924560547,
1.34756290912628,
4.19603824615479,
-5.57256841659546,
-4.34158897399902,
-2.95852327346802,
-10.2521562576294,
-8.47997379302979,
-4.26230239868164,
0.777846157550812,
-0.321977585554123,
15.9857015609741,
5.04163694381714,
-15.6162776947021,
-2.28500223159790,
8.47433757781982,
5.87041187286377,
16.5936794281006,
3.21923184394836,
-9.75627231597900,
-14.3114833831787,
-2.45077323913574,
17.3837203979492,
2.78194904327393,
9.99119758605957,
-11.6148347854614,
-17.5560169219971,
-5.00608158111572,
0.598314940929413,
-0.542393088340759,
-17.8817386627197,
2.80102300643921,
14.5387592315674,
9.74177074432373,
5.37954902648926,
14.7581052780151,
-3.13428068161011,
-9.93275451660156,
6.31521320343018,
-7.71506309509277,
-10.4804506301880,
-3.66732716560364,
-4.01443862915039,
-22.6006278991699,
-13.0657901763916,
-0.468873828649521,
-5.38479471206665,
-7.87983989715576,
-3.87705302238464,
6.02278661727905,
-14.2247076034546,
2.62369942665100,
2.68151640892029,
-5.02444744110107,
-4.50331592559814,
-13.7390003204346,
15.0099725723267,
8.22905158996582,
6.00241470336914,
11.1984052658081,
16.4483642578125,
-6.26652765274048,
2.01668930053711,
10.8875226974487,
-12.4427919387817,
-0.683354020118713,
-9.10700702667236,
10.7625274658203,
-10.9016561508179,
-9.38367557525635,
15.0269556045532,
-6.18128061294556,
-14.6435346603394,
-7.71684789657593,
2.76377153396606,
-11.5027427673340,
-0.513358592987061,
-5.00205802917481,
-8.55128574371338,
-12.9856281280518,
-11.0788021087646,
13.0642042160034,
-1.53834784030914,
-0.515877723693848,
-1.45037817955017,
1.02773964405060,
9.31696891784668,
-2.99124765396118,
5.20135688781738,
-1.34022021293640,
-9.37860202789307,
1.73207259178162,
0.392231374979019,
-5.62367820739746,
7.43250179290772,
2.66428971290588,
-15.3497104644775,
6.18619680404663,
-5.55827665328980,
-10.0966167449951,
11.3017177581787,
-18.2781314849854,
4.44812488555908,
8.89496803283691,
-25.2236156463623,
8.57238101959229,
5.90969705581665,
3.01573634147644,
-12.1820058822632,
4.32914972305298,
12.6482734680176,
-18.5440387725830,
13.7834854125977,
-9.24393367767334,
2.75513982772827,
1.76463019847870,
-13.8922882080078,
-9.92648601531982,
-7.00921726226807,
8.12637329101563,
-7.42727470397949,
-5.56471633911133,
-13.4729118347168,
9.61233711242676,
-10.8453245162964,
1.41092026233673,
2.20368576049805,
-20.1469478607178,
24.8114204406738,
-1.03763377666473,
11.0233078002930,
7.14627933502197,
-10.9356145858765,
5.29452991485596,
0.478690415620804,
4.93256282806397,
-8.36130142211914,
6.18539094924927,
7.66064786911011,
4.38745450973511,
8.14395809173584,
-0.201022386550903,
11.7246265411377,
-0.774272382259369,
-11.3871002197266,
2.63391160964966,
13.9538784027100,
5.87038707733154,
-5.30749702453613,
-4.08452320098877,
10.3934402465820,
6.58953952789307,
-2.09956288337708,
8.14958667755127,
-11.9306612014771,
-9.70180892944336,
17.3027915954590,
11.5910873413086,
-4.36236286163330,
-9.84329223632813,
3.41723275184631,
13.8209981918335,
-10.7073726654053,
0.154783621430397,
16.6939983367920,
-16.9452533721924,
3.07341766357422,
0.964140415191650,
-6.38871479034424,
2.73037719726563,
-22.1253242492676,
8.39183807373047,
-1.96543478965759,
-11.1584186553955,
0.686354994773865,
-3.00177574157715,
13.7714939117432,
-13.2152051925659,
9.41836833953857,
19.7016487121582,
-4.71853542327881,
0.594687581062317,
-9.94826889038086,
11.0317382812500,
5.24653387069702,
7.28536844253540,
1.02092003822327,
-13.4522666931152,
14.8550271987915,
8.56230449676514,
-5.59132337570190,
1.32905614376068,
1.74599182605743,
-25.8885955810547,
9.95198535919190,
-0.636754214763641,
-3.71522712707520,
8.49665832519531,
-18.5550193786621,
8.76062965393066,
-13.7832565307617,
11.1148681640625,
-4.92390441894531,
-11.2543659210205,
5.08325433731079,
-4.40541839599609,
19.9680957794189,
1.06059980392456,
-4.45308256149292,
-0.608428597450256,
15.2684946060181,
-2.03904604911804,
1.14522564411163,
7.64763212203980,
10.5258150100708,
4.08472681045532,
-9.54130172729492,
3.07381176948547,
-6.70701122283936,
12.0725784301758,
-8.15238857269287,
-1.42583179473877,
7.16194677352905,
-20.2166061401367,
4.52655744552612,
13.6177940368652,
6.26460552215576,
-6.42440986633301,
-1.96236097812653,
-3.43707680702209,
-7.66699981689453,
6.17506694793701,
-5.80379295349121,
-2.84858202934265,
-12.5326137542725,
-6.00326490402222,
20.8375415802002,
2.74026942253113,
5.74672555923462,
-4.15856695175171,
-1.23263490200043,
13.8602085113525,
-4.63936567306519,
-6.79918050765991,
1.45228135585785,
-0.223338365554810,
-19.4062061309814,
3.32435727119446,
-0.778049230575562,
-15.0435457229614,
20.4992179870605,
-1.36084902286530,
-12.8036069869995,
1.20373499393463,
-0.714227855205536,
-8.83776187896729,
-6.09387731552124,
17.2558116912842,
0.175023525953293,
-13.2315435409546,
-9.47945976257324,
9.35341167449951,
4.40458440780640,
-15.7020645141602,
8.33568000793457,
-1.74813365936279,
-13.5939931869507,
8.02303409576416,
0.752746641635895,
-15.7636890411377,
10.6147394180298,
-3.66670942306519,
-2.83081078529358,
8.42905235290527,
-16.7218208312988,
21.4410514831543,
11.1922683715820,
-15.1774291992188,
0.813959479331970,
7.16367864608765,
5.63329839706421,
6.81442689895630,
-5.17766141891480,
-11.9962291717529,
-4.10792636871338,
-18.6218051910400,
-1.17772746086121,
12.4196281433105,
7.17530870437622,
2.06803297996521,
-1.09778976440430,
1.19562470912933,
2.86692786216736,
11.7913808822632,
-4.07146024703980,
-1.66355073451996,
4.00092077255249,
-11.6694784164429,
13.2793817520142,
14.4351024627686,
3.95528674125671,
3.77485251426697,
0.726287782192230,
11.3287611007690,
-17.2514114379883,
1.66158711910248,
5.66137313842773,
-13.2494554519653,
-0.645135760307312,
-13.9465999603271,
1.97642982006073,
-2.06826376914978,
7.69320869445801,
-0.193779155611992,
-10.7201852798462,
3.84305477142334,
-8.25143814086914,
16.0336456298828,
11.6767206192017,
3.84674358367920,
-3.80574011802673,
-13.9865274429321,
3.87316966056824,
14.2519178390503,
2.78062844276428,
-7.68299722671509,
16.3278694152832,
-3.92920756340027,
-8.16404438018799,
19.8745059967041,
10.5993661880493,
-17.0135078430176,
-11.5570878982544,
14.8415870666504,
-14.0446214675903,
0.549165129661560,
15.6036796569824,
-4.97690916061401,
-12.9285125732422,
-2.09080719947815,
19.2437839508057,
10.3768148422241,
9.83218860626221,
3.06042575836182,
11.8945531845093,
14.6602497100830,
14.1966571807861,
-3.96037125587463,
-4.41946554183960,
0.507116377353668,
-7.93260431289673,
10.8404741287231,
2.38258385658264,
13.6977233886719,
0.688987076282501,
9.56145477294922,
6.76172876358032,
-11.3281288146973,
-2.80191659927368,
-16.3393554687500,
-6.74783802032471,
-10.8127136230469,
22.7601451873779,
0.306739240884781,
-15.5284976959229,
21.1589012145996,
-8.72752475738525,
10.5058450698853,
-5.25621986389160,
-0.491802692413330,
14.5102672576904,
-0.498369842767715,
16.1244812011719,
-9.73005008697510,
6.32857894897461,
-5.97241115570068,
-16.6271286010742,
13.5388860702515,
7.18867969512939,
-7.01135826110840,
-8.46527194976807,
12.4180850982666,
15.6671943664551,
0.622408211231232,
5.57255220413208,
13.5504617691040,
-11.4580154418945,
-13.7922172546387,
1.04516458511353,
-1.03297948837280,
-7.00995445251465,
-3.02339148521423,
-0.600792229175568,
1.09994709491730,
-3.55474925041199,
-12.1009330749512,
-6.95897340774536,
-6.19486761093140,
6.97705173492432,
10.7639217376709,
9.16511154174805,
8.19611454010010,
11.2818679809570,
12.7818861007690,
-1.80254101753235,
0.497679382562637,
11.1339941024780,
-2.39874672889709,
0.141300410032272,
18.5438995361328,
5.48683834075928,
-1.05251336097717,
5.54068708419800,
1.19009780883789,
-21.0975685119629,
2.77424001693726,
4.74189281463623,
-18.2863540649414,
11.9065265655518,
-12.4751234054565,
-11.3408699035645,
14.3046903610230,
3.29809641838074,
-3.43988347053528,
-13.5366897583008,
-9.41614532470703,
-2.00635695457459,
11.5155782699585,
-11.4248704910278,
-8.55550861358643,
17.4621658325195,
4.55207729339600,
4.00689125061035,
-7.85009479522705,
1.77085900306702,
8.50602626800537,
2.23359656333923,
11.7115297317505,
-0.227002546191216,
-10.7721538543701,
-12.8427705764771,
1.38814330101013,
-7.54678821563721,
-14.6243085861206,
10.9997062683105,
11.4011564254761,
3.25670409202576,
6.02790594100952,
9.33123207092285,
-7.11675453186035,
-0.0536885410547257,
3.16584658622742,
-1.80337405204773,
12.4571857452393,
-6.81064653396606,
9.13007068634033,
8.62425518035889,
-10.7262916564941,
14.4632854461670,
1.91948652267456,
-0.277435779571533,
0.539809823036194,
-14.3661994934082,
-6.58171987533569,
1.97790634632111,
8.39780521392822,
-0.365638345479965,
-13.8784847259521,
-2.91600728034973,
11.6675882339478,
-11.8000993728638,
9.95210266113281,
4.11969995498657,
-13.8756628036499,
10.3403072357178,
-9.14852714538574,
13.1162919998169,
-1.92573583126068,
-2.69105124473572,
8.30866432189941,
-10.4616975784302,
-4.70901012420654,
-1.78373277187347,
18.2263622283936,
-10.4992370605469,
-3.40257215499878,
18.5995273590088,
-7.55536127090454,
-6.98724985122681,
-6.53860521316528,
-14.7667312622070,
2.60888457298279,
0.561092555522919,
3.44232678413391,
11.6268739700317,
-14.4685535430908,
-8.14792442321777,
8.29515838623047,
10.4582691192627,
-2.48044657707214,
6.00418853759766,
6.03353738784790,
-12.0121583938599,
8.31047344207764,
7.56882572174072,
-1.20817184448242,
6.69751405715942,
-2.76144480705261,
-8.89453220367432,
13.3808279037476,
17.2055606842041,
-10.1105508804321,
-14.7115240097046,
8.30276298522949,
3.71625256538391,
4.43171262741089,
14.3717832565308,
8.89480590820313,
12.1071834564209,
7.88615846633911,
5.60394287109375,
-4.09735584259033,
5.60422945022583,
-5.76414537429810,
-6.04650783538818,
23.7772006988525,
-6.18358612060547,
-16.4450778961182,
-8.66361999511719,
-2.09574174880981,
4.57660102844238,
1.97597396373749,
-10.4837198257446,
-15.5591020584106,
-1.76396155357361,
-18.7482490539551,
10.0266885757446,
3.86129117012024,
-14.1002187728882,
16.6018028259277,
-4.37660837173462,
13.4767179489136,
16.9750194549561,
-8.76874351501465,
-3.75618982315063,
8.65848636627197,
-8.57310390472412,
-6.01041030883789,
12.5147600173950,
-12.6574020385742,
-1.81489372253418,
12.8609361648560,
3.31045126914978,
-4.34171104431152,
13.7912826538086,
3.67780494689941,
0.659437298774719,
4.47402524948120,
-20.5931873321533,
-1.69705665111542,
8.63898944854736,
-5.32576656341553,
-12.6602754592896,
-11.0770006179810,
-13.1143751144409,
7.70316457748413,
-6.41403675079346,
-13.8738927841187,
19.0773162841797,
0.903741180896759,
4.22006511688232,
14.1540660858154,
11.0694999694824,
11.2466220855713,
-13.0478496551514,
-11.3583049774170,
11.9404716491699,
1.48241436481476,
-2.41118741035461,
2.76930427551270,
-12.3991260528564,
-7.07537174224854,
-16.3161888122559,
-2.46065235137939,
13.5728921890259,
-18.6301269531250,
4.25361156463623,
3.62634539604187,
-2.26026678085327,
12.7831182479858,
-5.08231544494629,
-0.352847427129746,
-13.8504858016968,
-7.56887102127075,
4.30654525756836,
-2.38265371322632,
2.48432874679565,
-9.48580074310303,
5.33847618103027,
2.26496005058289,
-5.10286045074463,
12.9739589691162,
-1.18702292442322,
6.93916559219360,
-4.52792024612427,
-3.77836608886719,
17.6622428894043,
-0.848418474197388,
6.14435195922852,
-1.57494521141052,
-7.40130901336670,
-10.6943054199219,
-7.47540187835693,
11.2714653015137,
8.73961544036865,
5.45354318618774,
9.25389575958252,
12.1598863601685,
8.35356521606445,
1.51380825042725,
-4.37021732330322,
16.8267326354980,
-4.30764245986939,
-6.92706871032715,
12.8935689926147,
1.02213954925537,
6.60210704803467,
1.34360253810883,
9.87246608734131,
-6.17443990707398,
9.10684967041016,
14.2026166915894,
-1.50069618225098,
19.4121170043945,
-4.26626348495483,
-2.08827066421509,
7.33619403839111,
13.5415124893188,
7.27274465560913,
3.54309034347534,
0.0559295192360878,
-10.4255971908569,
17.7059974670410,
-3.33743143081665,
3.86344408988953,
6.16825437545776,
-7.71449136734009,
0.495854645967484,
-15.9373903274536,
4.60191488265991,
10.6833229064941,
1.02008616924286,
-2.84855532646179,
1.95340502262115,
-0.487840831279755,
13.8724536895752,
-2.17112565040588,
-8.48410034179688,
12.9616880416870,
-14.4692525863647,
16.0715293884277,
11.8501348495483,
-5.05098915100098,
-2.74764370918274,
-10.4964179992676,
5.46758031845093,
-8.67889022827148,
-11.9815616607666,
-2.84434914588928,
-8.61962985992432,
-18.0029869079590,
-8.81765365600586,
-11.4718246459961,
-6.48010683059692,
12.6888065338135,
-8.44581604003906,
-0.522065937519074,
17.4223041534424,
-6.71062183380127,
-9.52772998809815,
7.86700725555420,
-7.06833171844482,
-12.0232210159302,
4.20763969421387,
-6.67637109756470,
10.7153253555298,
-2.45592069625855,
-21.5680084228516,
9.00837421417236,
-12.2850198745728,
-11.5124721527100,
1.34292733669281,
0.372711718082428,
2.21345019340515,
-0.320124149322510,
10.5263404846191,
-10.7317466735840,
-7.14030265808106,
-0.0852114185690880,
6.51456975936890,
8.05042171478272,
-12.3626899719238,
11.4756336212158,
7.71447515487671,
12.7680444717407,
13.3046560287476,
-3.58520221710205,
13.2967443466187,
0.894922077655792,
-5.81144380569458,
-4.53378438949585,
-8.70451831817627,
-11.8104324340820,
11.8492336273193,
0.314905017614365,
-15.8788366317749,
-4.70532369613648,
-10.0715656280518,
12.4850139617920,
-15.7783346176147,
5.52781677246094,
6.53504896163940,
-9.35710334777832,
15.6052541732788,
-20.1759853363037,
10.9270067214966,
1.18999862670898,
-17.9319572448730,
13.0239429473877,
2.46298408508301,
6.71346426010132,
10.3850049972534,
-0.210399493575096,
-1.31163704395294,
15.4207916259766,
6.33792161941528,
-15.5164394378662,
-2.52922892570496,
8.40850830078125,
0.387925177812576,
-15.1006650924683,
-10.2033538818359,
8.94322109222412,
-8.66815471649170,
-8.42395210266113,
16.3662433624268,
-6.57894611358643,
-11.2145299911499,
14.3141479492188,
3.83258366584778,
6.87844991683960,
15.8383941650391,
8.44803142547607,
12.3757171630859,
5.70071840286255,
18.1221446990967,
0.108715265989304,
-8.24166011810303,
23.8793678283691,
10.0313930511475,
9.85764408111572,
-2.90879535675049,
-9.65310192108154,
2.73437643051147,
2.94620418548584,
15.7386369705200,
3.30390357971191,
7.64130830764771,
-8.10798072814941,
-5.44120550155640,
19.2188491821289,
-11.7892627716064,
7.29962682723999,
14.9086732864380,
-11.4114542007446,
-7.96764659881592,
-5.29620790481567,
-12.2225341796875,
-9.80076217651367,
-4.09044647216797,
11.2775774002075,
-4.61790418624878,
-16.0772895812988,
11.6125850677490,
-10.3969125747681,
-1.74642682075500,
-6.92615509033203,
-0.893892824649811,
9.36031913757324,
-6.60164785385132,
3.73657202720642,
-15.0439319610596,
-1.88126969337463,
10.5551471710205,
5.77378225326538,
-3.96806597709656,
3.60321998596191,
15.2608661651611,
2.53257679939270,
-7.57546281814575,
7.81377601623535,
5.04553842544556,
-13.9129438400269,
14.4900703430176,
-7.10630512237549,
-12.7281551361084,
9.91123962402344,
-11.7563161849976,
-4.73182868957520,
-1.02705180644989,
-12.1898832321167,
2.83993268013001,
-4.82621192932129,
-9.45471286773682,
7.25408649444580,
-11.0353355407715,
-11.8789358139038,
6.64584159851074,
9.33378982543945,
-7.70026636123657,
-19.0320358276367,
0.212033912539482,
8.96640396118164,
-3.27634549140930,
-15.5010833740234,
1.67470431327820,
-6.66629123687744,
-12.7931833267212,
12.4279966354370,
-6.57369804382324,
2.46465563774109,
1.04768764972687,
-8.57872390747070,
12.8037443161011,
5.12663412094116,
12.9414815902710,
-5.63042116165161,
-13.4960927963257,
-3.25135278701782,
0.850059568881989,
5.31062173843384,
-17.7165603637695,
4.06643104553223,
8.46233558654785,
8.55259990692139,
4.09808349609375,
-15.4935894012451,
0.267077326774597,
2.18488550186157,
7.03712892532349,
1.53150737285614,
3.75258183479309,
-9.35081768035889,
-2.70439028739929,
2.71083879470825,
-18.0917720794678,
-1.58555483818054,
-11.3625240325928,
-2.78137230873108,
-3.43628954887390,
-0.532094657421112,
16.6788177490234,
-14.5066699981689,
-17.3552684783936,
2.16126251220703,
11.8589639663696,
1.71788549423218,
11.3193130493164,
5.06808853149414,
-6.53804969787598,
14.1789503097534,
2.11391305923462,
5.67684459686279,
-1.04960656166077,
-6.19355106353760,
6.88596820831299,
7.14316844940186,
-11.3279781341553,
-2.67404651641846,
13.8031816482544,
-16.9676036834717,
7.56723690032959,
12.4425792694092,
-10.4620456695557,
-8.96198177337647,
-7.33463335037231,
12.5693063735962,
11.4362478256226,
0.167383670806885,
-1.61738908290863,
7.49672603607178,
12.7612457275391,
3.19251632690430,
-11.5457134246826,
-12.0060234069824,
8.35533046722412,
-4.57270574569702,
-13.5124206542969,
8.44027328491211,
-5.90609121322632,
-15.3930597305298,
-14.7790174484253,
-5.04672288894653,
8.40855026245117,
-14.6216583251953,
5.95415401458740,
18.7609672546387,
-0.581051051616669,
5.20874691009522,
4.43499898910523,
14.8158130645752,
3.59643745422363,
9.65670204162598,
2.66835069656372,
-9.74585056304932,
16.5832500457764,
3.90272831916809,
11.3035430908203,
-0.174154475331306,
1.90830123424530,
14.4682407379150,
-6.08135509490967,
0.960750043392181,
-2.20220971107483,
-3.01388430595398,
-15.1681079864502,
-0.941229760646820,
12.7969522476196,
-1.87731742858887,
2.13939690589905,
-4.61093664169312,
-4.09716558456421,
-8.24046230316162,
3.06720209121704,
14.7503261566162,
-9.22908115386963,
-9.95535850524902,
8.45219612121582,
6.88245820999146,
-13.1264677047730,
-12.5598974227905,
14.7678785324097,
0.268167018890381,
-15.5126914978027,
9.85108566284180,
-2.66498708724976,
2.21812844276428,
11.2758150100708,
-7.95464801788330,
8.97678184509277,
7.42069435119629,
7.03821420669556,
-1.26214349269867,
-2.74077749252319,
18.7821350097656,
-2.60253477096558,
11.6162900924683,
7.92783308029175,
-8.85243320465088,
12.9211006164551,
-11.1287822723389,
-15.6763620376587,
-7.18054342269898,
-11.1221380233765,
-11.7331676483154,
-12.2703523635864,
8.76590251922607,
3.89626646041870,
-0.186960548162460,
1.14144337177277,
-8.72398567199707,
-0.582658231258392,
1.40090560913086,
1.99565649032593,
-10.4684209823608,
-3.62940979003906,
19.1246871948242,
5.98375940322876,
5.73691463470459,
6.18672275543213,
-8.10184097290039,
5.13180494308472,
12.5598249435425,
-12.4011545181274,
-3.41500115394592,
16.2118530273438,
-1.90375447273254,
-19.4601554870605,
-0.768333017826080,
16.3412227630615,
-18.6500415802002,
-11.1755743026733,
8.84817028045654,
-15.7341003417969,
4.54690217971802,
19.2026615142822,
-6.35798406600952,
-13.0922899246216,
3.14263558387756,
13.4052705764771,
4.50402498245239,
9.78940486907959,
15.4542589187622,
0.599797368049622,
-5.56980562210083,
8.94028377532959,
12.8733930587769,
-5.92605829238892,
4.41021919250488,
14.1652784347534,
-10.3513231277466,
-0.427381426095963,
-3.38286542892456,
-12.3334064483643,
8.02093219757080,
-12.1592206954956,
-16.0060272216797,
-7.79566860198975,
-15.7042579650879,
-8.93447780609131,
7.25424528121948,
4.44127416610718,
6.23335456848145,
8.16137027740479,
-3.69512557983398,
1.21468329429626,
-9.06932163238525,
8.11106109619141,
3.80233621597290,
-3.70013070106506,
15.9114131927490,
-5.49834489822388,
-6.28960371017456,
11.9368133544922,
8.94310569763184,
-12.0432634353638,
-1.84292078018188,
-2.36310553550720,
-7.57056140899658,
1.56640243530273,
-14.4385585784912,
10.6375656127930,
0.464769750833511,
-14.8185272216797};
