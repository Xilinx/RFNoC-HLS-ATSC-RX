shortreal out[256] = '{0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
2.66733274356668e-10,
4.61779698923692e-08,
8.88920865804721e-08,
2.40675575469140e-07,
3.75603065094765e-07,
7.03452030847984e-07,
9.69933012129332e-07,
1.29138800275541e-06,
1.44344198815816e-06,
1.16488581625163e-06,
5.55104804789153e-07,
-1.50864423176245e-06,
-4.12428835261380e-06,
-9.97343886410818e-06,
-1.66061490745051e-05,
-2.93070279440144e-05,
-4.33042696386110e-05,
-6.28968482487835e-05,
-8.26158502604812e-05,
-0.000109618616988882,
-0.000135485097416677,
-0.000169940525665879,
-0.000196711524040438,
-0.000232703765504994,
-0.000269479904090986,
-0.000319680286338553,
-0.000365876738214865,
-0.000412882276577875,
-0.000463375705294311,
-0.000484685617266223,
-0.000518352142535150,
-0.000481719529489055,
-0.000460398208815604,
-0.000378229538910091,
-0.000304250832414255,
-0.000138650328153744,
3.90043060178869e-05,
0.000346178305335343,
0.000709121231921017,
0.00133546080905944,
0.00203764485195279,
0.000828407646622509,
-0.000164098266395740,
0.000443826109403744,
0.00152860209345818,
0.00253852317109704,
0.00246572657488287,
0.00145903252996504,
-0.00278176460415125,
-0.00930143520236015,
-0.0151211181655526,
-0.0211840625852346,
-0.0274639334529638,
-0.0331572517752647,
-0.0382524840533733,
-0.0402852371335030,
-0.0426312424242497,
-0.0488962978124619,
-0.0527118891477585,
-0.0558072961866856,
-0.0595176331698895,
-0.0636265948414803,
-0.0682977437973023,
-0.0723522379994392,
-0.0786263942718506,
-0.0834880322217941,
-0.0900844484567642,
-0.0977268517017365,
-0.102426938712597,
-0.106446087360382,
-0.110056966543198,
-0.113005034625530,
-0.112995333969593,
-0.115802332758904,
-0.120785333216190,
-0.124023377895355,
-0.129985094070435,
-0.138116985559464,
-0.145112141966820,
-0.149007260799408,
-0.152734398841858,
-0.155624285340309,
-0.157868370413780,
-0.162615567445755,
-0.164934813976288,
-0.165648058056831,
-0.166938826441765,
-0.166304692625999,
-0.165646821260452,
-0.166397407650948,
-0.165914252400398,
-0.165702477097511,
-0.168807461857796,
-0.173451632261276,
-0.180884554982185,
-0.191604703664780,
-0.205968424677849,
-0.222640424966812,
-0.237902969121933,
-0.252401411533356,
-0.267516911029816,
-0.283818393945694,
-0.301323086023331,
-0.323074132204056,
-0.344285577535629,
-0.366065919399262,
-0.391435056924820,
-0.413394212722778,
-0.436231315135956,
-0.461046218872070,
-0.487918585538864,
-0.515781342983246,
-0.542690634727478,
-0.572834849357605,
-0.602167546749115,
-0.628717839717865,
-0.654793381690979,
-0.681293725967407,
-0.711295187473297,
-0.741962134838104,
-0.770132780075073,
-0.800409078598023,
-0.831766486167908,
-0.861421883106232,
-0.891208231449127,
-0.923237681388855,
-0.957089722156525,
-0.989833295345306,
-1.02549278736115,
-1.05915129184723,
-1.09429097175598,
-1.12863922119141,
-1.16699731349945,
-1.19983541965485,
-1.24054110050201,
-1.27346599102020,
-1.30639815330505,
-1.34320008754730,
-1.35967159271240,
-1.41375851631165,
-1.40902137756348,
-1.48928344249725,
-1.44385445117950,
-1.56168282032013,
-1.53146159648895,
-1.66402149200439,
-1.59063935279846,
-1.77560651302338,
-1.66132295131683,
-1.97566211223602,
-1.74351978302002,
-1.93009102344513,
-1.77221107482910,
-2.10655736923218,
-2.07735800743103,
-2.08543753623962,
-2.67423486709595,
-2.04501700401306,
-3.45785474777222,
-2.10116052627563,
-3.40740656852722,
-2.32184433937073,
-4.01396083831787,
-2.75939559936523,
-4.74696207046509,
-3.58684921264648,
-7.06039142608643,
-4.03296995162964,
28.5958690643311,
-6.46929311752319,
-29.2790966033936,
-10.8618860244751,
-1.85944569110870,
14.6394586563110,
12.1251249313355,
49.8559417724609,
34.0829582214356,
-14.8897504806519,
0.546998322010040,
0.0616941004991531,
-13.1817846298218,
-13.4242677688599,
-53.9235954284668,
1.41867196559906,
60.5001068115234,
-43.9936714172363,
-15.6954030990601,
6.12152004241943,
2.51854372024536,
5.14021348953247,
-14.2292461395264,
32.1670761108398,
-27.3752059936523,
24.0887718200684,
12.7488117218018,
-52.5718345642090,
-15.6252298355103,
-11.2332286834717,
-15.4616622924805,
-53.0448799133301,
41.2601470947266,
30.7026271820068,
-33.3981590270996,
39.4755363464356,
30.3536262512207,
-23.6638984680176,
-55.7390747070313,
-7.99319791793823,
-18.9758110046387,
-15.9265842437744,
35.2927474975586,
-45.1014823913574,
-31.7794551849365,
3.67967939376831,
-37.1234207153320,
-6.27180528640747,
16.9350051879883,
-26.1258907318115,
-1.74089634418488,
47.6758651733398,
18.6767349243164,
38.8855247497559,
46.8841285705566,
52.5687522888184,
30.8023815155029,
-29.5765094757080,
-19.1707916259766,
3.15768241882324,
12.3086957931519,
12.5174455642700,
61.7739105224609,
-15.8419904708862,
2.05365490913391,
50.8995513916016,
-62.4646110534668};
