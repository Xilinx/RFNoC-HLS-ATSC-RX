shortreal in[32768] = '{0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
-1.00000000000000,1.00000000000000,
2.00000000000000,-1.00000000000000,
-3.00000000000000,1.00000000000000,
4.00000000000000,-2.00000000000000,
-7.00000000000000,2.00000000000000,
9.00000000000000,-3.00000000000000,
-13.0000000000000,4.00000000000000,
18.0000000000000,-5.00000000000000,
-26.0000000000000,7.00000000000000,
36.0000000000000,-9.00000000000000,
-53.0000000000000,15.0000000000000,
87.0000000000000,-27.0000000000000,
-243.000000000000,78.0000000000000,
-534.000000000000,321.000000000000,
-436.000000000000,-100.000000000000,
3.00000000000000,627.000000000000,
452.000000000000,-536.000000000000,
-256.000000000000,-957.000000000000,
100.000000000000,61.0000000000000,
183.000000000000,108.000000000000,
21.0000000000000,-780.000000000000,
280.000000000000,-1292.00000000000,
916.000000000000,-107.000000000000,
-54.0000000000000,-122.000000000000,
165.000000000000,-139.000000000000,
201.000000000000,631.000000000000,
-693.000000000000,-483.000000000000,
-85.0000000000000,-858.000000000000,
-268.000000000000,24.0000000000000,
926.000000000000,-324.000000000000,
1170.00000000000,-200.000000000000,
-369.000000000000,835.000000000000,
-174.000000000000,887.000000000000,
-21.0000000000000,819.000000000000,
59.0000000000000,-410.000000000000,
390.000000000000,-675.000000000000,
986.000000000000,240.000000000000,
-626.000000000000,-41.0000000000000,
-425.000000000000,665.000000000000,
117.000000000000,-1303.00000000000,
-860.000000000000,-96.0000000000000,
1030.00000000000,702.000000000000,
117.000000000000,-1260.00000000000,
47.0000000000000,-397.000000000000,
-202.000000000000,-599.000000000000,
-153.000000000000,856.000000000000,
-18.0000000000000,790.000000000000,
-1071.00000000000,-951.000000000000,
752.000000000000,-835.000000000000,
-396.000000000000,-437.000000000000,
-228.000000000000,-287.000000000000,
1066.00000000000,-351.000000000000,
729.000000000000,143.000000000000,
162.000000000000,-934.000000000000,
136.000000000000,-847.000000000000,
966.000000000000,-132.000000000000,
200.000000000000,409.000000000000,
665.000000000000,546.000000000000,
206.000000000000,228.000000000000,
-791.000000000000,109.000000000000,
242.000000000000,-1065.00000000000,
346.000000000000,549.000000000000,
-335.000000000000,847.000000000000,
-126.000000000000,-180.000000000000,
1328.00000000000,-321.000000000000,
566.000000000000,-113.000000000000,
-590.000000000000,465.000000000000,
-518.000000000000,-852.000000000000,
-434.000000000000,319.000000000000,
18.0000000000000,518.000000000000,
-109.000000000000,-229.000000000000,
746.000000000000,678.000000000000,
-345.000000000000,655.000000000000,
-1011.00000000000,216.000000000000,
942.000000000000,-646.000000000000,
407.000000000000,417.000000000000,
-618.000000000000,220.000000000000,
-1470.00000000000,489.000000000000,
-541.000000000000,-625.000000000000,
288.000000000000,-1029.00000000000,
-305.000000000000,904.000000000000,
-505.000000000000,-690.000000000000,
-1152.00000000000,-90.0000000000000,
123.000000000000,-273.000000000000,
981.000000000000,-295.000000000000,
480.000000000000,-378.000000000000,
22.0000000000000,-496.000000000000,
-487.000000000000,336.000000000000,
388.000000000000,-616.000000000000,
432.000000000000,388.000000000000,
-459.000000000000,-36.0000000000000,
81.0000000000000,567.000000000000,
489.000000000000,727.000000000000,
-819.000000000000,-892.000000000000,
757.000000000000,-612.000000000000,
1615.00000000000,-239.000000000000,
167.000000000000,105.000000000000,
418.000000000000,-1046.00000000000,
-409.000000000000,24.0000000000000,
296.000000000000,1090.00000000000,
154.000000000000,856.000000000000,
-789.000000000000,277.000000000000,
-115.000000000000,-1478.00000000000,
179.000000000000,-104.000000000000,
44.0000000000000,-183.000000000000,
-270.000000000000,283.000000000000,
1081.00000000000,233.000000000000,
-41.0000000000000,91.0000000000000,
-1001.00000000000,534.000000000000,
-682.000000000000,-1228.00000000000,
-747.000000000000,117.000000000000,
-578.000000000000,-59.0000000000000,
-450.000000000000,-1178.00000000000,
545.000000000000,-1102.00000000000,
-9.00000000000000,-561.000000000000,
-632.000000000000,561.000000000000,
-994.000000000000,-814.000000000000,
1124.00000000000,-412.000000000000,
625.000000000000,592.000000000000,
-758.000000000000,-800.000000000000,
655.000000000000,-302.000000000000,
-1017.00000000000,-174.000000000000,
320.000000000000,-469.000000000000,
868.000000000000,-70.0000000000000,
200.000000000000,-338.000000000000,
626.000000000000,-808.000000000000,
-216.000000000000,-275.000000000000,
207.000000000000,-371.000000000000,
-478.000000000000,-589.000000000000,
-465.000000000000,-450.000000000000,
581.000000000000,-467.000000000000,
987.000000000000,-71.0000000000000,
218.000000000000,-448.000000000000,
-531.000000000000,741.000000000000,
-686.000000000000,193.000000000000,
-706.000000000000,-641.000000000000,
507.000000000000,490.000000000000,
107.000000000000,697.000000000000,
-1193.00000000000,529.000000000000,
-313.000000000000,-723.000000000000,
-523.000000000000,-361.000000000000,
-566.000000000000,425.000000000000,
370.000000000000,-183.000000000000,
483.000000000000,-415.000000000000,
711.000000000000,393.000000000000,
-255.000000000000,706.000000000000,
-1712.00000000000,-547.000000000000,
-366.000000000000,-223.000000000000,
-217.000000000000,419.000000000000,
-698.000000000000,-745.000000000000,
1529.00000000000,-354.000000000000,
716.000000000000,299.000000000000,
-153.000000000000,335.000000000000,
-618.000000000000,459.000000000000,
48.0000000000000,611.000000000000,
445.000000000000,156.000000000000,
-567.000000000000,-694.000000000000,
922.000000000000,146.000000000000,
-411.000000000000,603.000000000000,
343.000000000000,486.000000000000,
842.000000000000,5.00000000000000,
-490.000000000000,1121.00000000000,
247.000000000000,810.000000000000,
-639.000000000000,-860.000000000000,
761.000000000000,-482.000000000000,
918.000000000000,20.0000000000000,
-122.000000000000,-382.000000000000,
446.000000000000,-764.000000000000,
-279.000000000000,152.000000000000,
-283.000000000000,-842.000000000000,
30.0000000000000,599.000000000000,
-696.000000000000,872.000000000000,
-889.000000000000,-1252.00000000000,
201.000000000000,800.000000000000,
-574.000000000000,199.000000000000,
72.0000000000000,-518.000000000000,
1223.00000000000,877.000000000000,
298.000000000000,549.000000000000,
586.000000000000,973.000000000000,
201.000000000000,862.000000000000,
-33.0000000000000,-759.000000000000,
-151.000000000000,-369.000000000000,
519.000000000000,-21.0000000000000,
1292.00000000000,-163.000000000000,
167.000000000000,764.000000000000,
-166.000000000000,301.000000000000,
0.00000000000000,448.000000000000,
381.000000000000,788.000000000000,
405.000000000000,181.000000000000,
-705.000000000000,347.000000000000,
-448.000000000000,-1410.00000000000,
44.0000000000000,-677.000000000000,
80.0000000000000,596.000000000000,
-618.000000000000,-668.000000000000,
-328.000000000000,-923.000000000000,
776.000000000000,125.000000000000,
28.0000000000000,1154.00000000000,
-7.00000000000000,-197.000000000000,
1032.00000000000,-142.000000000000,
-149.000000000000,423.000000000000,
-588.000000000000,-783.000000000000,
947.000000000000,-234.000000000000,
-914.000000000000,502.000000000000,
-630.000000000000,102.000000000000,
-101.000000000000,-172.000000000000,
-918.000000000000,9.00000000000000,
857.000000000000,135.000000000000,
634.000000000000,-266.000000000000,
161.000000000000,1100.00000000000,
-216.000000000000,551.000000000000,
-321.000000000000,-1142.00000000000,
32.0000000000000,-552.000000000000,
523.000000000000,350.000000000000,
412.000000000000,830.000000000000,
-585.000000000000,1245.00000000000,
300.000000000000,-1.00000000000000,
-495.000000000000,-1130.00000000000,
463.000000000000,-316.000000000000,
1838.00000000000,-229.000000000000,
-597.000000000000,689.000000000000,
-720.000000000000,44.0000000000000,
97.0000000000000,-132.000000000000,
31.0000000000000,315.000000000000,
-703.000000000000,-96.0000000000000,
-892.000000000000,-71.0000000000000,
951.000000000000,-1112.00000000000,
1271.00000000000,659.000000000000,
885.000000000000,659.000000000000,
506.000000000000,-300.000000000000,
-53.0000000000000,-698.000000000000,
-34.0000000000000,-1474.00000000000,
1003.00000000000,-234.000000000000,
710.000000000000,-282.000000000000,
257.000000000000,442.000000000000,
-23.0000000000000,863.000000000000,
-1013.00000000000,-488.000000000000,
747.000000000000,-652.000000000000,
1114.00000000000,-66.0000000000000,
375.000000000000,-473.000000000000,
181.000000000000,-673.000000000000,
-766.000000000000,742.000000000000,
247.000000000000,-437.000000000000,
594.000000000000,-626.000000000000,
-430.000000000000,779.000000000000,
-337.000000000000,-75.0000000000000,
407.000000000000,-889.000000000000,
35.0000000000000,-686.000000000000,
-40.0000000000000,134.000000000000,
-244.000000000000,670.000000000000,
-246.000000000000,797.000000000000,
-596.000000000000,748.000000000000,
-890.000000000000,-272.000000000000,
955.000000000000,251.000000000000,
-62.0000000000000,423.000000000000,
-295.000000000000,-220.000000000000,
1062.00000000000,-150.000000000000,
244.000000000000,-395.000000000000,
517.000000000000,383.000000000000,
-346.000000000000,217.000000000000,
-268.000000000000,-1221.00000000000,
366.000000000000,-623.000000000000,
-525.000000000000,943.000000000000,
-599.000000000000,126.000000000000,
537.000000000000,-434.000000000000,
288.000000000000,-176.000000000000,
-1092.00000000000,-247.000000000000,
329.000000000000,1051.00000000000,
174.000000000000,426.000000000000,
717.000000000000,-60.0000000000000,
395.000000000000,125.000000000000,
-1023.00000000000,-673.000000000000,
495.000000000000,181.000000000000,
352.000000000000,221.000000000000,
-582.000000000000,471.000000000000,
-1220.00000000000,-361.000000000000,
344.000000000000,-731.000000000000,
71.0000000000000,790.000000000000,
-184.000000000000,54.0000000000000,
976.000000000000,-796.000000000000,
-769.000000000000,-296.000000000000,
695.000000000000,115.000000000000,
249.000000000000,-480.000000000000,
-1012.00000000000,550.000000000000,
111.000000000000,895.000000000000,
-264.000000000000,-517.000000000000,
-507.000000000000,104.000000000000,
-131.000000000000,348.000000000000,
-328.000000000000,-336.000000000000,
-865.000000000000,-210.000000000000,
894.000000000000,708.000000000000,
-321.000000000000,-41.0000000000000,
-468.000000000000,-29.0000000000000,
1133.00000000000,246.000000000000,
-679.000000000000,68.0000000000000,
-446.000000000000,863.000000000000,
-1103.00000000000,-534.000000000000,
-288.000000000000,-283.000000000000,
334.000000000000,88.0000000000000,
-608.000000000000,-766.000000000000,
30.0000000000000,574.000000000000,
-476.000000000000,-238.000000000000,
-154.000000000000,-951.000000000000,
-384.000000000000,334.000000000000,
-553.000000000000,261.000000000000,
-423.000000000000,-1239.00000000000,
651.000000000000,-693.000000000000,
666.000000000000,743.000000000000,
-1067.00000000000,810.000000000000,
106.000000000000,-185.000000000000,
540.000000000000,-394.000000000000,
354.000000000000,432.000000000000,
443.000000000000,318.000000000000,
-80.0000000000000,1105.00000000000,
-437.000000000000,345.000000000000,
-557.000000000000,-38.0000000000000,
-57.0000000000000,-150.000000000000,
-831.000000000000,-883.000000000000,
-165.000000000000,947.000000000000,
-470.000000000000,249.000000000000,
91.0000000000000,-368.000000000000,
832.000000000000,-75.0000000000000,
-444.000000000000,-802.000000000000,
413.000000000000,319.000000000000,
-643.000000000000,-182.000000000000,
-244.000000000000,-784.000000000000,
331.000000000000,-685.000000000000,
615.000000000000,-339.000000000000,
790.000000000000,102.000000000000,
-192.000000000000,382.000000000000,
32.0000000000000,1054.00000000000,
-985.000000000000,-192.000000000000,
-122.000000000000,-304.000000000000,
-476.000000000000,420.000000000000,
-441.000000000000,283.000000000000,
174.000000000000,617.000000000000,
-1110.00000000000,-6.00000000000000,
-173.000000000000,-675.000000000000,
433.000000000000,474.000000000000,
-800.000000000000,634.000000000000,
-479.000000000000,-201.000000000000,
-658.000000000000,-257.000000000000,
-608.000000000000,-4.00000000000000,
-390.000000000000,96.0000000000000,
259.000000000000,-1438.00000000000,
958.000000000000,316.000000000000,
-917.000000000000,689.000000000000,
-805.000000000000,-777.000000000000,
-404.000000000000,-505.000000000000,
395.000000000000,-1313.00000000000,
567.000000000000,158.000000000000,
140.000000000000,-383.000000000000,
542.000000000000,-50.0000000000000,
-492.000000000000,956.000000000000,
-645.000000000000,-224.000000000000,
-22.0000000000000,808.000000000000,
612.000000000000,-202.000000000000,
741.000000000000,-441.000000000000,
-95.0000000000000,-95.0000000000000,
-1201.00000000000,-159.000000000000,
312.000000000000,679.000000000000,
222.000000000000,39.0000000000000,
-748.000000000000,-248.000000000000,
-223.000000000000,-35.0000000000000,
-122.000000000000,111.000000000000,
610.000000000000,-754.000000000000,
203.000000000000,-105.000000000000,
481.000000000000,1100.00000000000,
605.000000000000,66.0000000000000,
882.000000000000,282.000000000000,
-111.000000000000,670.000000000000,
-1513.00000000000,615.000000000000,
-155.000000000000,-1015.00000000000,
-30.0000000000000,-1330.00000000000,
96.0000000000000,-72.0000000000000,
-186.000000000000,-1120.00000000000,
-586.000000000000,-1007.00000000000,
917.000000000000,-230.000000000000,
659.000000000000,-406.000000000000,
-320.000000000000,451.000000000000,
371.000000000000,706.000000000000,
160.000000000000,-488.000000000000,
128.000000000000,-32.0000000000000,
-225.000000000000,200.000000000000,
-1471.00000000000,-744.000000000000,
187.000000000000,-326.000000000000,
223.000000000000,543.000000000000,
-737.000000000000,-540.000000000000,
571.000000000000,-535.000000000000,
86.0000000000000,-196.000000000000,
920.000000000000,-66.0000000000000,
110.000000000000,288.000000000000,
-378.000000000000,539.000000000000,
1169.00000000000,-212.000000000000,
-264.000000000000,258.000000000000,
990.000000000000,474.000000000000,
516.000000000000,-566.000000000000,
-408.000000000000,657.000000000000,
-19.0000000000000,65.0000000000000,
-993.000000000000,-527.000000000000,
-410.000000000000,-289.000000000000,
494.000000000000,80.0000000000000,
721.000000000000,-428.000000000000,
-474.000000000000,-733.000000000000,
-464.000000000000,329.000000000000,
-192.000000000000,-467.000000000000,
1010.00000000000,-57.0000000000000,
405.000000000000,-491.000000000000,
-872.000000000000,-44.0000000000000,
443.000000000000,687.000000000000,
-318.000000000000,-965.000000000000,
822.000000000000,-143.000000000000,
121.000000000000,172.000000000000,
-566.000000000000,882.000000000000,
-40.0000000000000,1002.00000000000,
-433.000000000000,-559.000000000000,
1326.00000000000,9.00000000000000,
-64.0000000000000,-157.000000000000,
-69.0000000000000,-731.000000000000,
-218.000000000000,365.000000000000,
-1267.00000000000,272.000000000000,
125.000000000000,-1439.00000000000,
451.000000000000,975.000000000000,
160.000000000000,997.000000000000,
-535.000000000000,-139.000000000000,
743.000000000000,641.000000000000,
151.000000000000,-303.000000000000,
-390.000000000000,948.000000000000,
818.000000000000,-295.000000000000,
-247.000000000000,193.000000000000,
-125.000000000000,1228.00000000000,
-544.000000000000,480.000000000000,
-150.000000000000,477.000000000000,
663.000000000000,-403.000000000000,
1426.00000000000,222.000000000000,
712.000000000000,-584.000000000000,
-426.000000000000,-910.000000000000,
270.000000000000,-1021.00000000000,
-577.000000000000,-909.000000000000,
-45.0000000000000,-536.000000000000,
-277.000000000000,-977.000000000000,
611.000000000000,252.000000000000,
1643.00000000000,412.000000000000,
-591.000000000000,1301.00000000000,
-517.000000000000,865.000000000000,
39.0000000000000,146.000000000000,
328.000000000000,955.000000000000,
-31.0000000000000,560.000000000000,
-329.000000000000,-62.0000000000000,
-823.000000000000,-1114.00000000000,
538.000000000000,-244.000000000000,
1238.00000000000,-264.000000000000,
-533.000000000000,-169.000000000000,
-73.0000000000000,806.000000000000,
-603.000000000000,-343.000000000000,
577.000000000000,135.000000000000,
6.00000000000000,436.000000000000,
-1667.00000000000,162.000000000000,
-303.000000000000,-901.000000000000,
-627.000000000000,-691.000000000000,
1207.00000000000,-16.0000000000000,
-154.000000000000,-21.0000000000000,
-1206.00000000000,449.000000000000,
801.000000000000,-557.000000000000,
-229.000000000000,1051.00000000000,
-604.000000000000,425.000000000000,
-900.000000000000,89.0000000000000,
269.000000000000,-503.000000000000,
528.000000000000,-417.000000000000,
48.0000000000000,1137.00000000000,
680.000000000000,-871.000000000000,
75.0000000000000,580.000000000000,
-255.000000000000,305.000000000000,
-394.000000000000,136.000000000000,
85.0000000000000,449.000000000000,
-986.000000000000,-282.000000000000,
-608.000000000000,392.000000000000,
-154.000000000000,8.00000000000000,
-330.000000000000,745.000000000000,
345.000000000000,-916.000000000000,
-299.000000000000,-1166.00000000000,
455.000000000000,-650.000000000000,
-466.000000000000,-1138.00000000000,
-485.000000000000,457.000000000000,
-528.000000000000,-298.000000000000,
205.000000000000,-306.000000000000,
1103.00000000000,-620.000000000000,
-146.000000000000,-744.000000000000,
870.000000000000,-241.000000000000,
-224.000000000000,414.000000000000,
-46.0000000000000,683.000000000000,
56.0000000000000,-1157.00000000000,
383.000000000000,-488.000000000000,
1762.00000000000,132.000000000000,
-141.000000000000,910.000000000000,
-122.000000000000,51.0000000000000,
372.000000000000,-224.000000000000,
-343.000000000000,405.000000000000,
-923.000000000000,-506.000000000000,
-1294.00000000000,157.000000000000,
-1014.00000000000,-379.000000000000,
-958.000000000000,-127.000000000000,
-154.000000000000,-830.000000000000,
411.000000000000,-236.000000000000,
1101.00000000000,949.000000000000,
-417.000000000000,-137.000000000000,
-71.0000000000000,618.000000000000,
915.000000000000,-492.000000000000,
-499.000000000000,812.000000000000,
41.0000000000000,972.000000000000,
-1485.00000000000,-600.000000000000,
-290.000000000000,-789.000000000000,
1347.00000000000,-579.000000000000,
615.000000000000,991.000000000000,
1333.00000000000,-85.0000000000000,
500.000000000000,-216.000000000000,
326.000000000000,-565.000000000000,
986.000000000000,-337.000000000000,
941.000000000000,780.000000000000,
-273.000000000000,589.000000000000,
-575.000000000000,100.000000000000,
-151.000000000000,-859.000000000000,
-589.000000000000,175.000000000000,
-610.000000000000,-490.000000000000,
-501.000000000000,-162.000000000000,
916.000000000000,387.000000000000,
308.000000000000,-332.000000000000,
306.000000000000,480.000000000000,
-51.0000000000000,-1322.00000000000,
-197.000000000000,-105.000000000000,
966.000000000000,690.000000000000,
144.000000000000,-674.000000000000,
1122.00000000000,421.000000000000,
-412.000000000000,-167.000000000000,
113.000000000000,-635.000000000000,
992.000000000000,-186.000000000000,
-182.000000000000,778.000000000000,
1408.00000000000,505.000000000000,
308.000000000000,341.000000000000,
-359.000000000000,-36.0000000000000,
721.000000000000,-243.000000000000,
554.000000000000,420.000000000000,
600.000000000000,335.000000000000,
800.000000000000,300.000000000000,
481.000000000000,-462.000000000000,
-509.000000000000,925.000000000000,
-299.000000000000,495.000000000000,
27.0000000000000,339.000000000000,
-116.000000000000,1693.00000000000,
-344.000000000000,15.0000000000000,
-225.000000000000,16.0000000000000,
751.000000000000,218.000000000000,
-253.000000000000,559.000000000000,
-769.000000000000,805.000000000000,
635.000000000000,-242.000000000000,
352.000000000000,-86.0000000000000,
-1106.00000000000,-148.000000000000,
-213.000000000000,-265.000000000000,
146.000000000000,-113.000000000000,
-175.000000000000,-667.000000000000,
384.000000000000,-790.000000000000,
-438.000000000000,-470.000000000000,
520.000000000000,-843.000000000000,
1042.00000000000,126.000000000000,
-87.0000000000000,738.000000000000,
683.000000000000,-322.000000000000,
453.000000000000,476.000000000000,
-1179.00000000000,744.000000000000,
-508.000000000000,-789.000000000000,
536.000000000000,-547.000000000000,
-713.000000000000,-135.000000000000,
-599.000000000000,759.000000000000,
-318.000000000000,716.000000000000,
-4.00000000000000,-540.000000000000,
665.000000000000,353.000000000000,
-403.000000000000,1503.00000000000,
142.000000000000,730.000000000000,
-470.000000000000,-122.000000000000,
-723.000000000000,657.000000000000,
101.000000000000,682.000000000000,
-276.000000000000,323.000000000000,
-707.000000000000,407.000000000000,
-961.000000000000,-816.000000000000,
-110.000000000000,-45.0000000000000,
98.0000000000000,248.000000000000,
368.000000000000,-649.000000000000,
-230.000000000000,550.000000000000,
-798.000000000000,644.000000000000,
173.000000000000,-420.000000000000,
311.000000000000,-512.000000000000,
-36.0000000000000,85.0000000000000,
89.0000000000000,401.000000000000,
-241.000000000000,-86.0000000000000,
-803.000000000000,-698.000000000000,
-653.000000000000,-176.000000000000,
-936.000000000000,-73.0000000000000,
-241.000000000000,-1016.00000000000,
1361.00000000000,142.000000000000,
802.000000000000,938.000000000000,
-203.000000000000,397.000000000000,
-345.000000000000,554.000000000000,
167.000000000000,-185.000000000000,
796.000000000000,-36.0000000000000,
609.000000000000,83.0000000000000,
-477.000000000000,-148.000000000000,
284.000000000000,273.000000000000,
460.000000000000,-482.000000000000,
-111.000000000000,189.000000000000,
-46.0000000000000,36.0000000000000,
-287.000000000000,-55.0000000000000,
334.000000000000,478.000000000000,
-427.000000000000,107.000000000000,
10.0000000000000,669.000000000000,
-22.0000000000000,857.000000000000,
-1283.00000000000,52.0000000000000,
-732.000000000000,-390.000000000000,
379.000000000000,310.000000000000,
400.000000000000,308.000000000000,
-727.000000000000,-193.000000000000,
-1142.00000000000,-420.000000000000,
-254.000000000000,383.000000000000,
-93.0000000000000,250.000000000000,
-11.0000000000000,-603.000000000000,
94.0000000000000,-213.000000000000,
366.000000000000,-299.000000000000,
859.000000000000,-723.000000000000,
-634.000000000000,-616.000000000000,
-71.0000000000000,866.000000000000,
-94.0000000000000,749.000000000000,
29.0000000000000,-232.000000000000,
632.000000000000,-772.000000000000,
81.0000000000000,-388.000000000000,
534.000000000000,1297.00000000000,
-841.000000000000,564.000000000000,
-526.000000000000,153.000000000000,
647.000000000000,188.000000000000,
261.000000000000,-33.0000000000000,
-222.000000000000,65.0000000000000,
-1065.00000000000,305.000000000000,
-711.000000000000,-591.000000000000,
-400.000000000000,-1422.00000000000,
1034.00000000000,-313.000000000000,
632.000000000000,798.000000000000,
-508.000000000000,1185.00000000000,
510.000000000000,-361.000000000000,
568.000000000000,391.000000000000,
743.000000000000,67.0000000000000,
91.0000000000000,-241.000000000000,
87.0000000000000,807.000000000000,
-128.000000000000,-529.000000000000,
-581.000000000000,966.000000000000,
-314.000000000000,631.000000000000,
-460.000000000000,-1205.00000000000,
-155.000000000000,-333.000000000000,
-108.000000000000,364.000000000000,
675.000000000000,481.000000000000,
-311.000000000000,-722.000000000000,
473.000000000000,86.0000000000000,
88.0000000000000,338.000000000000,
-357.000000000000,-677.000000000000,
1296.00000000000,-170.000000000000,
-910.000000000000,123.000000000000,
-822.000000000000,486.000000000000,
-312.000000000000,520.000000000000,
-61.0000000000000,677.000000000000,
515.000000000000,150.000000000000,
117.000000000000,751.000000000000,
722.000000000000,68.0000000000000,
136.000000000000,-1110.00000000000,
58.0000000000000,-277.000000000000,
-66.0000000000000,-1413.00000000000,
537.000000000000,-121.000000000000,
523.000000000000,1509.00000000000,
-9.00000000000000,-345.000000000000,
177.000000000000,74.0000000000000,
758.000000000000,465.000000000000,
-47.0000000000000,-44.0000000000000,
-946.000000000000,321.000000000000,
491.000000000000,-135.000000000000,
-58.0000000000000,-117.000000000000,
-611.000000000000,213.000000000000,
555.000000000000,671.000000000000,
-85.0000000000000,405.000000000000,
-469.000000000000,-463.000000000000,
350.000000000000,289.000000000000,
122.000000000000,1552.00000000000,
-786.000000000000,-151.000000000000,
-154.000000000000,-1411.00000000000,
-159.000000000000,86.0000000000000,
-583.000000000000,135.000000000000,
1334.00000000000,-506.000000000000,
754.000000000000,198.000000000000,
-546.000000000000,58.0000000000000,
-160.000000000000,-905.000000000000,
-57.0000000000000,310.000000000000,
61.0000000000000,176.000000000000,
-580.000000000000,755.000000000000,
386.000000000000,154.000000000000,
18.0000000000000,-261.000000000000,
-693.000000000000,1183.00000000000,
-817.000000000000,-126.000000000000,
-891.000000000000,292.000000000000,
783.000000000000,-701.000000000000,
166.000000000000,178.000000000000,
517.000000000000,886.000000000000,
-16.0000000000000,-478.000000000000,
-438.000000000000,-9.00000000000000,
-310.000000000000,-451.000000000000,
-470.000000000000,798.000000000000,
1087.00000000000,-312.000000000000,
895.000000000000,134.000000000000,
225.000000000000,1393.00000000000,
-1375.00000000000,-102.000000000000,
-1069.00000000000,71.0000000000000,
-269.000000000000,-355.000000000000,
99.0000000000000,36.0000000000000,
-232.000000000000,-626.000000000000,
-516.000000000000,-489.000000000000,
292.000000000000,862.000000000000,
-956.000000000000,-429.000000000000,
814.000000000000,-857.000000000000,
956.000000000000,236.000000000000,
62.0000000000000,613.000000000000,
564.000000000000,340.000000000000,
-1150.00000000000,449.000000000000,
-580.000000000000,-637.000000000000,
209.000000000000,342.000000000000,
238.000000000000,712.000000000000,
265.000000000000,-1573.00000000000,
-257.000000000000,-701.000000000000,
784.000000000000,-178.000000000000,
579.000000000000,626.000000000000,
-209.000000000000,898.000000000000,
-98.0000000000000,770.000000000000,
242.000000000000,-300.000000000000,
-208.000000000000,-559.000000000000,
230.000000000000,460.000000000000,
281.000000000000,-1399.00000000000,
-322.000000000000,792.000000000000,
600.000000000000,308.000000000000,
-645.000000000000,-1235.00000000000,
635.000000000000,886.000000000000,
-315.000000000000,157.000000000000,
-1702.00000000000,228.000000000000,
-271.000000000000,-500.000000000000,
-114.000000000000,152.000000000000,
1181.00000000000,-233.000000000000,
69.0000000000000,-241.000000000000,
212.000000000000,465.000000000000,
494.000000000000,285.000000000000,
-420.000000000000,836.000000000000,
-1021.00000000000,-906.000000000000,
-72.0000000000000,-717.000000000000,
1276.00000000000,-735.000000000000,
-562.000000000000,-306.000000000000,
-37.0000000000000,-2.00000000000000,
387.000000000000,-1743.00000000000,
-549.000000000000,-450.000000000000,
30.0000000000000,140.000000000000,
-234.000000000000,-517.000000000000,
-299.000000000000,-42.0000000000000,
1053.00000000000,357.000000000000,
968.000000000000,743.000000000000,
-426.000000000000,779.000000000000,
-44.0000000000000,-585.000000000000,
-74.0000000000000,-737.000000000000,
4.00000000000000,457.000000000000,
231.000000000000,334.000000000000,
-893.000000000000,131.000000000000,
-66.0000000000000,-36.0000000000000,
573.000000000000,404.000000000000,
-408.000000000000,232.000000000000,
93.0000000000000,-154.000000000000,
58.0000000000000,868.000000000000,
-512.000000000000,309.000000000000,
-358.000000000000,479.000000000000,
310.000000000000,-509.000000000000,
-342.000000000000,-851.000000000000,
92.0000000000000,-471.000000000000,
1010.00000000000,-758.000000000000,
-485.000000000000,1091.00000000000,
317.000000000000,-458.000000000000,
119.000000000000,-252.000000000000,
-162.000000000000,-264.000000000000,
717.000000000000,-1097.00000000000,
767.000000000000,724.000000000000,
-367.000000000000,170.000000000000,
-197.000000000000,855.000000000000,
374.000000000000,677.000000000000,
-934.000000000000,294.000000000000,
-52.0000000000000,482.000000000000,
-428.000000000000,538.000000000000,
-1192.00000000000,287.000000000000,
-1151.00000000000,-483.000000000000,
-637.000000000000,316.000000000000,
749.000000000000,350.000000000000,
-396.000000000000,485.000000000000,
-488.000000000000,-112.000000000000,
865.000000000000,-15.0000000000000,
1131.00000000000,-68.0000000000000,
96.0000000000000,-467.000000000000,
-958.000000000000,183.000000000000,
-360.000000000000,-1399.00000000000,
-132.000000000000,-1276.00000000000,
-23.0000000000000,-491.000000000000,
69.0000000000000,-419.000000000000,
245.000000000000,513.000000000000,
567.000000000000,455.000000000000,
951.000000000000,207.000000000000,
231.000000000000,-862.000000000000,
-109.000000000000,-919.000000000000,
108.000000000000,-404.000000000000,
-301.000000000000,-42.0000000000000,
1021.00000000000,636.000000000000,
303.000000000000,-153.000000000000,
430.000000000000,645.000000000000,
-59.0000000000000,476.000000000000,
-308.000000000000,-789.000000000000,
1145.00000000000,442.000000000000,
19.0000000000000,130.000000000000,
674.000000000000,-726.000000000000,
539.000000000000,-236.000000000000,
-622.000000000000,521.000000000000,
-289.000000000000,86.0000000000000,
-15.0000000000000,-434.000000000000,
668.000000000000,432.000000000000,
-184.000000000000,747.000000000000,
-748.000000000000,-486.000000000000,
1102.00000000000,-630.000000000000,
973.000000000000,525.000000000000,
-332.000000000000,730.000000000000,
53.0000000000000,320.000000000000,
385.000000000000,59.0000000000000,
843.000000000000,322.000000000000,
174.000000000000,74.0000000000000,
-1361.00000000000,666.000000000000,
-727.000000000000,-272.000000000000,
177.000000000000,-1164.00000000000,
-750.000000000000,113.000000000000,
-402.000000000000,-672.000000000000,
35.0000000000000,165.000000000000,
-467.000000000000,1495.00000000000,
-720.000000000000,-33.0000000000000,
-896.000000000000,208.000000000000,
-898.000000000000,-495.000000000000,
635.000000000000,-1038.00000000000,
247.000000000000,135.000000000000,
-365.000000000000,-422.000000000000,
326.000000000000,691.000000000000,
-67.0000000000000,591.000000000000,
1002.00000000000,428.000000000000,
-561.000000000000,221.000000000000,
-153.000000000000,-603.000000000000,
1233.00000000000,370.000000000000,
35.0000000000000,-512.000000000000,
-231.000000000000,-265.000000000000,
-871.000000000000,179.000000000000,
463.000000000000,28.0000000000000,
-684.000000000000,649.000000000000,
-1212.00000000000,458.000000000000,
239.000000000000,-570.000000000000,
-1258.00000000000,25.0000000000000,
-204.000000000000,-358.000000000000,
838.000000000000,-1255.00000000000,
76.0000000000000,-704.000000000000,
277.000000000000,-516.000000000000,
-473.000000000000,253.000000000000,
155.000000000000,-396.000000000000,
1488.00000000000,193.000000000000,
412.000000000000,1285.00000000000,
-152.000000000000,702.000000000000,
203.000000000000,421.000000000000,
-1173.00000000000,-349.000000000000,
-534.000000000000,28.0000000000000,
758.000000000000,772.000000000000,
-1382.00000000000,392.000000000000,
-510.000000000000,-375.000000000000,
505.000000000000,-49.0000000000000,
-680.000000000000,-381.000000000000,
558.000000000000,-313.000000000000,
372.000000000000,-485.000000000000,
-88.0000000000000,-716.000000000000,
948.000000000000,692.000000000000,
1007.00000000000,-138.000000000000,
332.000000000000,761.000000000000,
-133.000000000000,1318.00000000000,
299.000000000000,-37.0000000000000,
675.000000000000,490.000000000000,
1219.00000000000,309.000000000000,
49.0000000000000,688.000000000000,
-699.000000000000,504.000000000000,
-755.000000000000,361.000000000000,
-347.000000000000,561.000000000000,
-414.000000000000,691.000000000000,
-930.000000000000,734.000000000000,
417.000000000000,-434.000000000000,
317.000000000000,-26.0000000000000,
-381.000000000000,-997.000000000000,
-123.000000000000,-894.000000000000,
537.000000000000,110.000000000000,
-318.000000000000,-1073.00000000000,
-39.0000000000000,511.000000000000,
-14.0000000000000,876.000000000000,
-973.000000000000,-203.000000000000,
320.000000000000,-215.000000000000,
335.000000000000,809.000000000000,
894.000000000000,-255.000000000000,
-27.0000000000000,-308.000000000000,
-45.0000000000000,1309.00000000000,
389.000000000000,-993.000000000000,
-695.000000000000,-891.000000000000,
1092.00000000000,-463.000000000000,
97.0000000000000,92.0000000000000,
-364.000000000000,-418.000000000000,
168.000000000000,-1097.00000000000,
-180.000000000000,-80.0000000000000,
84.0000000000000,-860.000000000000,
-68.0000000000000,1273.00000000000,
125.000000000000,305.000000000000,
-216.000000000000,-578.000000000000,
364.000000000000,1048.00000000000,
-534.000000000000,-677.000000000000,
-711.000000000000,-701.000000000000,
-156.000000000000,-298.000000000000,
-78.0000000000000,-1312.00000000000,
712.000000000000,-391.000000000000,
7.00000000000000,1353.00000000000,
-150.000000000000,406.000000000000,
61.0000000000000,-830.000000000000,
-13.0000000000000,-48.0000000000000,
-406.000000000000,-950.000000000000,
637.000000000000,-358.000000000000,
255.000000000000,1063.00000000000,
-194.000000000000,-225.000000000000,
691.000000000000,-591.000000000000,
-50.0000000000000,-577.000000000000,
-30.0000000000000,2.00000000000000,
-466.000000000000,-534.000000000000,
171.000000000000,-1135.00000000000,
-231.000000000000,363.000000000000,
-559.000000000000,-328.000000000000,
1105.00000000000,-742.000000000000,
347.000000000000,698.000000000000,
197.000000000000,533.000000000000,
534.000000000000,-503.000000000000,
559.000000000000,701.000000000000,
395.000000000000,817.000000000000,
-242.000000000000,-484.000000000000,
1084.00000000000,-410.000000000000,
749.000000000000,392.000000000000,
-723.000000000000,683.000000000000,
307.000000000000,-215.000000000000,
-76.0000000000000,-494.000000000000,
-339.000000000000,357.000000000000,
501.000000000000,304.000000000000,
-45.0000000000000,-914.000000000000,
306.000000000000,-22.0000000000000,
597.000000000000,-708.000000000000,
-93.0000000000000,-878.000000000000,
-121.000000000000,494.000000000000,
-306.000000000000,-415.000000000000,
-1305.00000000000,-47.0000000000000,
540.000000000000,-449.000000000000,
932.000000000000,-93.0000000000000,
-279.000000000000,-18.0000000000000,
435.000000000000,-1199.00000000000,
418.000000000000,436.000000000000,
398.000000000000,742.000000000000,
98.0000000000000,181.000000000000,
639.000000000000,-110.000000000000,
699.000000000000,95.0000000000000,
-97.0000000000000,377.000000000000,
-135.000000000000,316.000000000000,
-725.000000000000,517.000000000000,
-739.000000000000,-183.000000000000,
107.000000000000,28.0000000000000,
17.0000000000000,872.000000000000,
-372.000000000000,543.000000000000,
492.000000000000,-407.000000000000,
180.000000000000,211.000000000000,
300.000000000000,497.000000000000,
408.000000000000,-743.000000000000,
-21.0000000000000,53.0000000000000,
645.000000000000,271.000000000000,
-342.000000000000,861.000000000000,
-658.000000000000,1044.00000000000,
-535.000000000000,-538.000000000000,
435.000000000000,-261.000000000000,
562.000000000000,-509.000000000000,
-200.000000000000,903.000000000000,
-280.000000000000,795.000000000000,
-1243.00000000000,58.0000000000000,
40.0000000000000,-49.0000000000000,
-891.000000000000,-755.000000000000,
101.000000000000,1014.00000000000,
548.000000000000,-809.000000000000,
-557.000000000000,-771.000000000000,
178.000000000000,-81.0000000000000,
-1210.00000000000,-634.000000000000,
444.000000000000,426.000000000000,
-84.0000000000000,304.000000000000,
67.0000000000000,-89.0000000000000,
639.000000000000,-317.000000000000,
-314.000000000000,1573.00000000000,
480.000000000000,538.000000000000,
-374.000000000000,876.000000000000,
453.000000000000,-7.00000000000000,
-117.000000000000,-966.000000000000,
-290.000000000000,1253.00000000000,
437.000000000000,424.000000000000,
-766.000000000000,744.000000000000,
-780.000000000000,78.0000000000000,
-886.000000000000,-384.000000000000,
-196.000000000000,113.000000000000,
579.000000000000,-69.0000000000000,
458.000000000000,706.000000000000,
-145.000000000000,976.000000000000,
-794.000000000000,934.000000000000,
-918.000000000000,-165.000000000000,
219.000000000000,24.0000000000000,
197.000000000000,581.000000000000,
-161.000000000000,-136.000000000000,
1397.00000000000,555.000000000000,
-291.000000000000,-261.000000000000,
-410.000000000000,118.000000000000,
-21.0000000000000,754.000000000000,
39.0000000000000,-282.000000000000,
1240.00000000000,156.000000000000,
349.000000000000,-303.000000000000,
335.000000000000,53.0000000000000,
-1351.00000000000,-131.000000000000,
580.000000000000,-461.000000000000,
971.000000000000,-104.000000000000,
-1340.00000000000,687.000000000000,
953.000000000000,-235.000000000000,
-374.000000000000,35.0000000000000,
-107.000000000000,1392.00000000000,
659.000000000000,-1028.00000000000,
-800.000000000000,-511.000000000000,
482.000000000000,403.000000000000,
-343.000000000000,476.000000000000,
-1208.00000000000,-101.000000000000,
-177.000000000000,-91.0000000000000,
317.000000000000,-268.000000000000,
-246.000000000000,-1525.00000000000,
1206.00000000000,-99.0000000000000,
161.000000000000,-301.000000000000,
-539.000000000000,565.000000000000,
853.000000000000,429.000000000000,
-714.000000000000,-367.000000000000,
802.000000000000,888.000000000000,
608.000000000000,3.00000000000000,
-537.000000000000,572.000000000000,
-594.000000000000,317.000000000000,
-1290.00000000000,-571.000000000000,
-7.00000000000000,-471.000000000000,
47.0000000000000,393.000000000000,
-239.000000000000,905.000000000000,
-754.000000000000,198.000000000000,
-135.000000000000,41.0000000000000,
355.000000000000,164.000000000000,
-2.00000000000000,1096.00000000000,
825.000000000000,4.00000000000000,
708.000000000000,-107.000000000000,
1202.00000000000,-28.0000000000000,
52.0000000000000,-465.000000000000,
288.000000000000,731.000000000000,
-57.0000000000000,-687.000000000000,
-1099.00000000000,609.000000000000,
410.000000000000,-317.000000000000,
45.0000000000000,-993.000000000000,
977.000000000000,572.000000000000,
1257.00000000000,-239.000000000000,
906.000000000000,1145.00000000000,
-1017.00000000000,-3.00000000000000,
-18.0000000000000,-276.000000000000,
999.000000000000,70.0000000000000,
-1424.00000000000,-373.000000000000,
-530.000000000000,176.000000000000,
-537.000000000000,-1073.00000000000,
1278.00000000000,-20.0000000000000,
680.000000000000,129.000000000000,
-430.000000000000,898.000000000000,
-92.0000000000000,1142.00000000000,
-232.000000000000,-720.000000000000,
888.000000000000,978.000000000000,
-865.000000000000,860.000000000000,
-483.000000000000,-686.000000000000,
-219.000000000000,-397.000000000000,
-409.000000000000,198.000000000000,
-257.000000000000,-582.000000000000,
175.000000000000,148.000000000000,
1030.00000000000,133.000000000000,
-352.000000000000,-1038.00000000000,
-525.000000000000,555.000000000000,
-994.000000000000,-754.000000000000,
308.000000000000,-818.000000000000,
325.000000000000,78.0000000000000,
-342.000000000000,-1008.00000000000,
640.000000000000,364.000000000000,
-150.000000000000,325.000000000000,
1440.00000000000,-229.000000000000,
1072.00000000000,570.000000000000,
-666.000000000000,463.000000000000,
-17.0000000000000,189.000000000000,
160.000000000000,627.000000000000,
116.000000000000,-874.000000000000,
-57.0000000000000,-286.000000000000,
110.000000000000,1564.00000000000,
-867.000000000000,-506.000000000000,
-636.000000000000,-191.000000000000,
-548.000000000000,120.000000000000,
-946.000000000000,75.0000000000000,
267.000000000000,1228.00000000000,
-438.000000000000,437.000000000000,
-546.000000000000,290.000000000000,
76.0000000000000,420.000000000000,
830.000000000000,-46.0000000000000,
961.000000000000,-139.000000000000,
-40.0000000000000,1158.00000000000,
-237.000000000000,-526.000000000000,
-122.000000000000,-1048.00000000000,
1394.00000000000,113.000000000000,
561.000000000000,-304.000000000000,
496.000000000000,642.000000000000,
689.000000000000,102.000000000000,
-1513.00000000000,289.000000000000,
-274.000000000000,435.000000000000,
75.0000000000000,258.000000000000,
-257.000000000000,-175.000000000000,
-318.000000000000,-298.000000000000,
-785.000000000000,-60.0000000000000,
111.000000000000,-846.000000000000,
-865.000000000000,497.000000000000,
-441.000000000000,-854.000000000000,
641.000000000000,-41.0000000000000,
907.000000000000,866.000000000000,
-76.0000000000000,-589.000000000000,
546.000000000000,708.000000000000,
1162.00000000000,-363.000000000000,
184.000000000000,-537.000000000000,
-151.000000000000,312.000000000000,
-376.000000000000,811.000000000000,
71.0000000000000,1119.00000000000,
-1208.00000000000,-498.000000000000,
461.000000000000,-734.000000000000,
1077.00000000000,-542.000000000000,
669.000000000000,1008.00000000000,
330.000000000000,340.000000000000,
-593.000000000000,-647.000000000000,
591.000000000000,702.000000000000,
-1251.00000000000,-201.000000000000,
-604.000000000000,940.000000000000,
-510.000000000000,28.0000000000000,
-552.000000000000,-1368.00000000000,
803.000000000000,-321.000000000000,
-478.000000000000,-121.000000000000,
-117.000000000000,-76.0000000000000,
180.000000000000,-728.000000000000,
410.000000000000,-335.000000000000,
-504.000000000000,526.000000000000,
-788.000000000000,600.000000000000,
947.000000000000,-89.0000000000000,
543.000000000000,241.000000000000,
-195.000000000000,487.000000000000,
-114.000000000000,780.000000000000,
-1044.00000000000,558.000000000000,
-1353.00000000000,-937.000000000000,
68.0000000000000,-711.000000000000,
-53.0000000000000,-404.000000000000,
17.0000000000000,-778.000000000000,
1724.00000000000,-128.000000000000,
964.000000000000,464.000000000000,
-226.000000000000,-558.000000000000,
443.000000000000,-489.000000000000,
311.000000000000,-224.000000000000,
162.000000000000,-23.0000000000000,
-426.000000000000,988.000000000000,
-104.000000000000,-293.000000000000,
620.000000000000,680.000000000000,
-412.000000000000,2065.00000000000,
-550.000000000000,-52.0000000000000,
-480.000000000000,-1070.00000000000,
117.000000000000,-9.00000000000000,
525.000000000000,741.000000000000,
-215.000000000000,-260.000000000000,
-618.000000000000,-612.000000000000,
-166.000000000000,11.0000000000000,
475.000000000000,164.000000000000,
-120.000000000000,-373.000000000000,
-169.000000000000,-313.000000000000,
263.000000000000,936.000000000000,
-76.0000000000000,136.000000000000,
-695.000000000000,-853.000000000000,
-155.000000000000,-288.000000000000,
53.0000000000000,486.000000000000,
-616.000000000000,-380.000000000000,
422.000000000000,-527.000000000000,
-118.000000000000,332.000000000000,
-1002.00000000000,-47.0000000000000,
-362.000000000000,817.000000000000,
-722.000000000000,611.000000000000,
-168.000000000000,77.0000000000000,
520.000000000000,-132.000000000000,
721.000000000000,-316.000000000000,
-195.000000000000,589.000000000000,
5.00000000000000,625.000000000000,
158.000000000000,83.0000000000000,
-140.000000000000,-381.000000000000,
918.000000000000,21.0000000000000,
-135.000000000000,-594.000000000000,
-239.000000000000,58.0000000000000,
-207.000000000000,684.000000000000,
-90.0000000000000,-671.000000000000,
90.0000000000000,846.000000000000,
46.0000000000000,1042.00000000000,
282.000000000000,564.000000000000,
-765.000000000000,165.000000000000,
-822.000000000000,-416.000000000000,
-550.000000000000,781.000000000000,
142.000000000000,328.000000000000,
-637.000000000000,780.000000000000,
86.0000000000000,173.000000000000,
565.000000000000,38.0000000000000,
-1253.00000000000,641.000000000000,
-839.000000000000,-567.000000000000,
-178.000000000000,609.000000000000,
198.000000000000,-648.000000000000,
-95.0000000000000,-1272.00000000000,
932.000000000000,299.000000000000,
387.000000000000,760.000000000000,
-1130.00000000000,966.000000000000,
-927.000000000000,-794.000000000000,
-297.000000000000,-969.000000000000,
665.000000000000,-456.000000000000,
722.000000000000,-127.000000000000,
423.000000000000,1256.00000000000,
-963.000000000000,770.000000000000,
-753.000000000000,277.000000000000,
-313.000000000000,770.000000000000,
-1011.00000000000,408.000000000000,
-1334.00000000000,-703.000000000000,
127.000000000000,37.0000000000000,
421.000000000000,414.000000000000,
-899.000000000000,-111.000000000000,
852.000000000000,389.000000000000,
-146.000000000000,-920.000000000000,
292.000000000000,-423.000000000000,
1623.00000000000,-95.0000000000000,
-284.000000000000,-412.000000000000,
214.000000000000,-37.0000000000000,
-845.000000000000,-67.0000000000000,
-179.000000000000,189.000000000000,
783.000000000000,-437.000000000000,
658.000000000000,1076.00000000000,
1063.00000000000,-22.0000000000000,
82.0000000000000,58.0000000000000,
756.000000000000,1155.00000000000,
-274.000000000000,-275.000000000000,
60.0000000000000,-705.000000000000,
210.000000000000,-935.000000000000,
95.0000000000000,-203.000000000000,
1023.00000000000,-249.000000000000,
-100.000000000000,1633.00000000000,
-36.0000000000000,1120.00000000000,
-787.000000000000,405.000000000000,
-78.0000000000000,408.000000000000,
-257.000000000000,-1291.00000000000,
-844.000000000000,257.000000000000,
546.000000000000,507.000000000000,
305.000000000000,298.000000000000,
775.000000000000,-152.000000000000,
69.0000000000000,310.000000000000,
-698.000000000000,716.000000000000,
-736.000000000000,107.000000000000,
-179.000000000000,1426.00000000000,
-520.000000000000,162.000000000000,
-170.000000000000,-240.000000000000,
1736.00000000000,-60.0000000000000,
-336.000000000000,111.000000000000,
-21.0000000000000,170.000000000000,
597.000000000000,-230.000000000000,
-809.000000000000,472.000000000000,
-663.000000000000,-523.000000000000,
-1190.00000000000,-166.000000000000,
-893.000000000000,-27.0000000000000,
215.000000000000,-509.000000000000,
-266.000000000000,215.000000000000,
-225.000000000000,311.000000000000,
870.000000000000,817.000000000000,
-631.000000000000,-19.0000000000000,
-332.000000000000,-760.000000000000,
675.000000000000,-419.000000000000,
-24.0000000000000,-1082.00000000000,
437.000000000000,-166.000000000000,
-40.0000000000000,984.000000000000,
-8.00000000000000,183.000000000000,
531.000000000000,217.000000000000,
316.000000000000,229.000000000000,
149.000000000000,-716.000000000000,
47.0000000000000,-54.0000000000000,
690.000000000000,-475.000000000000,
-493.000000000000,-344.000000000000,
-358.000000000000,1071.00000000000,
-286.000000000000,-921.000000000000,
-1055.00000000000,-313.000000000000,
204.000000000000,-1035.00000000000,
589.000000000000,-841.000000000000,
1107.00000000000,953.000000000000,
-748.000000000000,255.000000000000,
324.000000000000,397.000000000000,
536.000000000000,-794.000000000000,
-518.000000000000,-687.000000000000,
1032.00000000000,-1294.00000000000,
-839.000000000000,-352.000000000000,
-42.0000000000000,-596.000000000000,
-584.000000000000,-927.000000000000,
-501.000000000000,677.000000000000,
1006.00000000000,-94.0000000000000,
-503.000000000000,1276.00000000000,
559.000000000000,-339.000000000000,
911.000000000000,-394.000000000000,
290.000000000000,851.000000000000,
-1179.00000000000,-25.0000000000000,
-321.000000000000,-1024.00000000000,
526.000000000000,-1100.00000000000,
-699.000000000000,891.000000000000,
-470.000000000000,-518.000000000000,
-839.000000000000,-160.000000000000,
-207.000000000000,31.0000000000000,
-1131.00000000000,-159.000000000000,
-352.000000000000,-102.000000000000,
437.000000000000,-1270.00000000000,
859.000000000000,844.000000000000,
1095.00000000000,-370.000000000000,
-210.000000000000,-630.000000000000,
1044.00000000000,-595.000000000000,
-335.000000000000,-185.000000000000,
113.000000000000,1341.00000000000,
415.000000000000,160.000000000000,
-367.000000000000,1665.00000000000,
-471.000000000000,395.000000000000,
-977.000000000000,-1113.00000000000,
1058.00000000000,-519.000000000000,
109.000000000000,-308.000000000000,
-130.000000000000,296.000000000000,
733.000000000000,82.0000000000000,
-17.0000000000000,650.000000000000,
-312.000000000000,603.000000000000,
11.0000000000000,150.000000000000,
-255.000000000000,-820.000000000000,
-539.000000000000,-393.000000000000,
214.000000000000,706.000000000000,
-424.000000000000,771.000000000000,
401.000000000000,619.000000000000,
724.000000000000,453.000000000000,
-404.000000000000,979.000000000000,
735.000000000000,-24.0000000000000,
726.000000000000,-357.000000000000,
-149.000000000000,730.000000000000,
-141.000000000000,-363.000000000000,
-345.000000000000,-778.000000000000,
-189.000000000000,290.000000000000,
575.000000000000,-305.000000000000,
-305.000000000000,-312.000000000000,
-151.000000000000,1294.00000000000,
-6.00000000000000,769.000000000000,
-1406.00000000000,-311.000000000000,
82.0000000000000,339.000000000000,
-67.0000000000000,-900.000000000000,
-560.000000000000,-172.000000000000,
500.000000000000,793.000000000000,
50.0000000000000,-51.0000000000000,
188.000000000000,1307.00000000000,
-387.000000000000,675.000000000000,
926.000000000000,135.000000000000,
239.000000000000,114.000000000000,
-856.000000000000,337.000000000000,
140.000000000000,-633.000000000000,
-391.000000000000,-983.000000000000,
641.000000000000,-803.000000000000,
243.000000000000,-1290.00000000000,
539.000000000000,273.000000000000,
-146.000000000000,42.0000000000000,
-248.000000000000,503.000000000000,
1109.00000000000,121.000000000000,
-550.000000000000,349.000000000000,
394.000000000000,514.000000000000,
523.000000000000,-348.000000000000,
505.000000000000,191.000000000000,
349.000000000000,-605.000000000000,
-450.000000000000,956.000000000000,
-368.000000000000,707.000000000000,
-1701.00000000000,-62.0000000000000,
38.0000000000000,-657.000000000000,
974.000000000000,-444.000000000000,
384.000000000000,1643.00000000000,
-1164.00000000000,-244.000000000000,
-1315.00000000000,-220.000000000000,
-173.000000000000,-1196.00000000000,
394.000000000000,-1241.00000000000,
1340.00000000000,912.000000000000,
695.000000000000,359.000000000000,
991.000000000000,819.000000000000,
-721.000000000000,456.000000000000,
-622.000000000000,133.000000000000,
151.000000000000,-514.000000000000,
-745.000000000000,-872.000000000000,
343.000000000000,-869.000000000000,
-152.000000000000,-460.000000000000,
329.000000000000,488.000000000000,
-367.000000000000,-102.000000000000,
-11.0000000000000,-4.00000000000000,
1315.00000000000,62.0000000000000,
-394.000000000000,1354.00000000000,
157.000000000000,415.000000000000,
-586.000000000000,-31.0000000000000,
-1021.00000000000,395.000000000000,
32.0000000000000,-1251.00000000000,
333.000000000000,-1047.00000000000,
614.000000000000,-901.000000000000,
-304.000000000000,631.000000000000,
-339.000000000000,-353.000000000000,
-861.000000000000,100.000000000000,
700.000000000000,849.000000000000,
-193.000000000000,-1152.00000000000,
-445.000000000000,451.000000000000,
1424.00000000000,15.0000000000000,
110.000000000000,796.000000000000,
-124.000000000000,1286.00000000000,
-480.000000000000,-732.000000000000,
-281.000000000000,-429.000000000000,
125.000000000000,71.0000000000000,
495.000000000000,66.0000000000000,
701.000000000000,-404.000000000000,
871.000000000000,281.000000000000,
-19.0000000000000,667.000000000000,
-438.000000000000,-109.000000000000,
729.000000000000,-654.000000000000,
466.000000000000,-1093.00000000000,
408.000000000000,-220.000000000000,
-48.0000000000000,715.000000000000,
59.0000000000000,-729.000000000000,
288.000000000000,-784.000000000000,
72.0000000000000,487.000000000000,
284.000000000000,215.000000000000,
476.000000000000,-274.000000000000,
112.000000000000,91.0000000000000,
-1245.00000000000,-275.000000000000,
-1015.00000000000,-124.000000000000,
-43.0000000000000,-269.000000000000,
284.000000000000,-537.000000000000,
927.000000000000,-307.000000000000,
318.000000000000,-1112.00000000000,
378.000000000000,-497.000000000000,
534.000000000000,-618.000000000000,
682.000000000000,39.0000000000000,
272.000000000000,139.000000000000,
80.0000000000000,-681.000000000000,
802.000000000000,-21.0000000000000,
-418.000000000000,-426.000000000000,
986.000000000000,426.000000000000,
149.000000000000,187.000000000000,
-681.000000000000,-20.0000000000000,
134.000000000000,301.000000000000,
-1541.00000000000,376.000000000000,
257.000000000000,-618.000000000000,
531.000000000000,-128.000000000000,
536.000000000000,981.000000000000,
1068.00000000000,-330.000000000000,
-565.000000000000,647.000000000000,
-1017.00000000000,-421.000000000000,
-1417.00000000000,-460.000000000000,
-271.000000000000,467.000000000000,
-28.0000000000000,259.000000000000,
418.000000000000,757.000000000000,
319.000000000000,-340.000000000000,
-458.000000000000,242.000000000000,
-465.000000000000,-302.000000000000,
-527.000000000000,-343.000000000000,
973.000000000000,-275.000000000000,
706.000000000000,-237.000000000000,
260.000000000000,1015.00000000000,
-540.000000000000,645.000000000000,
-714.000000000000,1101.00000000000,
-270.000000000000,859.000000000000,
-326.000000000000,334.000000000000,
1123.00000000000,-58.0000000000000,
-237.000000000000,-239.000000000000,
-718.000000000000,-369.000000000000,
12.0000000000000,-53.0000000000000,
-951.000000000000,934.000000000000,
-717.000000000000,-249.000000000000,
270.000000000000,55.0000000000000,
99.0000000000000,1099.00000000000,
-898.000000000000,547.000000000000,
-1040.00000000000,-73.0000000000000,
-874.000000000000,-601.000000000000,
-634.000000000000,-1026.00000000000,
446.000000000000,-853.000000000000,
261.000000000000,391.000000000000,
-355.000000000000,932.000000000000,
-294.000000000000,-59.0000000000000,
528.000000000000,-1178.00000000000,
35.0000000000000,241.000000000000,
-120.000000000000,683.000000000000,
920.000000000000,-495.000000000000,
549.000000000000,1068.00000000000,
-532.000000000000,445.000000000000,
-1026.00000000000,-843.000000000000,
-586.000000000000,-252.000000000000,
-902.000000000000,-237.000000000000,
-730.000000000000,96.0000000000000,
-348.000000000000,-934.000000000000,
430.000000000000,-417.000000000000,
1236.00000000000,-159.000000000000,
369.000000000000,-504.000000000000,
1576.00000000000,115.000000000000,
70.0000000000000,-639.000000000000,
-1124.00000000000,164.000000000000,
-895.000000000000,-696.000000000000,
-693.000000000000,-805.000000000000,
961.000000000000,-147.000000000000,
456.000000000000,659.000000000000,
1300.00000000000,386.000000000000,
133.000000000000,-204.000000000000,
336.000000000000,915.000000000000,
820.000000000000,-701.000000000000,
-410.000000000000,-266.000000000000,
709.000000000000,428.000000000000,
-889.000000000000,335.000000000000,
2.00000000000000,-505.000000000000,
552.000000000000,453.000000000000,
-528.000000000000,341.000000000000,
332.000000000000,-1886.00000000000,
-314.000000000000,519.000000000000,
104.000000000000,487.000000000000,
-651.000000000000,298.000000000000,
-1149.00000000000,684.000000000000,
-23.0000000000000,-260.000000000000,
893.000000000000,519.000000000000,
18.0000000000000,-359.000000000000,
-211.000000000000,-603.000000000000,
66.0000000000000,-1061.00000000000,
309.000000000000,-1079.00000000000,
919.000000000000,-602.000000000000,
-192.000000000000,-1176.00000000000,
218.000000000000,17.0000000000000,
-661.000000000000,-62.0000000000000,
63.0000000000000,113.000000000000,
1089.00000000000,900.000000000000,
-469.000000000000,466.000000000000,
217.000000000000,-775.000000000000,
211.000000000000,-1235.00000000000,
-65.0000000000000,-192.000000000000,
-53.0000000000000,-537.000000000000,
410.000000000000,-769.000000000000,
151.000000000000,-536.000000000000,
-1009.00000000000,-244.000000000000,
95.0000000000000,-51.0000000000000,
165.000000000000,681.000000000000,
-933.000000000000,417.000000000000,
-590.000000000000,-945.000000000000,
352.000000000000,-23.0000000000000,
632.000000000000,49.0000000000000,
419.000000000000,4.00000000000000,
272.000000000000,-496.000000000000,
-720.000000000000,-528.000000000000,
604.000000000000,602.000000000000,
548.000000000000,411.000000000000,
354.000000000000,883.000000000000,
834.000000000000,96.0000000000000,
64.0000000000000,299.000000000000,
696.000000000000,300.000000000000,
-135.000000000000,-266.000000000000,
-669.000000000000,198.000000000000,
-1022.00000000000,-182.000000000000,
-948.000000000000,-272.000000000000,
147.000000000000,-1237.00000000000,
930.000000000000,-261.000000000000,
367.000000000000,848.000000000000,
-596.000000000000,-580.000000000000,
105.000000000000,83.0000000000000,
603.000000000000,428.000000000000,
-396.000000000000,-221.000000000000,
-600.000000000000,528.000000000000,
935.000000000000,168.000000000000,
-24.0000000000000,-730.000000000000,
40.0000000000000,-207.000000000000,
1562.00000000000,249.000000000000,
-736.000000000000,147.000000000000,
-603.000000000000,258.000000000000,
364.000000000000,-1574.00000000000,
70.0000000000000,-283.000000000000,
941.000000000000,1227.00000000000,
82.0000000000000,186.000000000000,
-446.000000000000,779.000000000000,
-657.000000000000,-13.0000000000000,
98.0000000000000,-337.000000000000,
256.000000000000,403.000000000000,
-511.000000000000,399.000000000000,
-44.0000000000000,-869.000000000000,
-157.000000000000,190.000000000000,
931.000000000000,673.000000000000,
441.000000000000,-948.000000000000,
103.000000000000,-816.000000000000,
1181.00000000000,-369.000000000000,
821.000000000000,211.000000000000,
45.0000000000000,-356.000000000000,
-748.000000000000,-577.000000000000,
605.000000000000,-900.000000000000,
-30.0000000000000,-650.000000000000,
-734.000000000000,-308.000000000000,
841.000000000000,-126.000000000000,
-494.000000000000,773.000000000000,
-599.000000000000,582.000000000000,
-498.000000000000,562.000000000000,
-420.000000000000,-604.000000000000,
249.000000000000,-430.000000000000,
-493.000000000000,-384.000000000000,
-22.0000000000000,-17.0000000000000,
-364.000000000000,718.000000000000,
-475.000000000000,-453.000000000000,
453.000000000000,762.000000000000,
695.000000000000,457.000000000000,
-257.000000000000,-184.000000000000,
-453.000000000000,1190.00000000000,
43.0000000000000,373.000000000000,
-139.000000000000,-39.0000000000000,
-681.000000000000,12.0000000000000,
205.000000000000,-1127.00000000000,
274.000000000000,-141.000000000000,
190.000000000000,921.000000000000,
868.000000000000,872.000000000000,
-186.000000000000,-940.000000000000,
503.000000000000,-76.0000000000000,
-535.000000000000,394.000000000000,
-217.000000000000,-663.000000000000,
326.000000000000,803.000000000000,
-1107.00000000000,-329.000000000000,
1057.00000000000,-127.000000000000,
471.000000000000,-168.000000000000,
724.000000000000,-420.000000000000,
462.000000000000,-379.000000000000,
-769.000000000000,545.000000000000,
-257.000000000000,653.000000000000,
-1795.00000000000,-600.000000000000,
187.000000000000,-362.000000000000,
279.000000000000,-1357.00000000000,
-735.000000000000,149.000000000000,
-220.000000000000,-26.0000000000000,
-513.000000000000,-298.000000000000,
896.000000000000,-110.000000000000,
214.000000000000,-823.000000000000,
586.000000000000,-313.000000000000,
593.000000000000,327.000000000000,
-761.000000000000,746.000000000000,
-615.000000000000,-116.000000000000,
-824.000000000000,345.000000000000,
-334.000000000000,-1020.00000000000,
-838.000000000000,-681.000000000000,
130.000000000000,-291.000000000000,
-95.0000000000000,-884.000000000000,
-107.000000000000,1397.00000000000,
-54.0000000000000,268.000000000000,
-1339.00000000000,146.000000000000,
-591.000000000000,-421.000000000000,
-1012.00000000000,-607.000000000000,
376.000000000000,414.000000000000,
601.000000000000,-420.000000000000,
-67.0000000000000,100.000000000000,
698.000000000000,-124.000000000000,
650.000000000000,443.000000000000,
350.000000000000,462.000000000000,
-194.000000000000,-271.000000000000,
1364.00000000000,294.000000000000,
702.000000000000,742.000000000000,
-1442.00000000000,232.000000000000,
-489.000000000000,146.000000000000,
-225.000000000000,811.000000000000,
-772.000000000000,584.000000000000,
-345.000000000000,142.000000000000,
-483.000000000000,-125.000000000000,
-700.000000000000,251.000000000000,
-468.000000000000,-381.000000000000,
-605.000000000000,-418.000000000000,
-548.000000000000,465.000000000000,
-464.000000000000,-1134.00000000000,
-667.000000000000,-260.000000000000,
-27.0000000000000,561.000000000000,
110.000000000000,-1155.00000000000,
666.000000000000,593.000000000000,
176.000000000000,903.000000000000,
349.000000000000,-654.000000000000,
3.00000000000000,-1311.00000000000,
-516.000000000000,-26.0000000000000,
783.000000000000,305.000000000000,
-543.000000000000,-407.000000000000,
-366.000000000000,787.000000000000,
-1224.00000000000,-371.000000000000,
-1144.00000000000,224.000000000000,
760.000000000000,646.000000000000,
-728.000000000000,691.000000000000,
-771.000000000000,541.000000000000,
-586.000000000000,-1247.00000000000,
-103.000000000000,102.000000000000,
116.000000000000,227.000000000000,
361.000000000000,-313.000000000000,
529.000000000000,802.000000000000,
-860.000000000000,451.000000000000,
-275.000000000000,-695.000000000000,
943.000000000000,-548.000000000000,
-98.0000000000000,-494.000000000000,
-1273.00000000000,-417.000000000000,
-524.000000000000,374.000000000000,
-618.000000000000,206.000000000000,
-311.000000000000,586.000000000000,
512.000000000000,-487.000000000000,
712.000000000000,-597.000000000000,
803.000000000000,1003.00000000000,
-1041.00000000000,-462.000000000000,
-423.000000000000,425.000000000000,
64.0000000000000,458.000000000000,
-929.000000000000,-712.000000000000,
-837.000000000000,-274.000000000000,
-53.0000000000000,-1140.00000000000,
1118.00000000000,109.000000000000,
-916.000000000000,155.000000000000,
-243.000000000000,-811.000000000000,
1217.00000000000,260.000000000000,
-546.000000000000,287.000000000000,
371.000000000000,-1084.00000000000,
-53.0000000000000,-374.000000000000,
-531.000000000000,-217.000000000000,
754.000000000000,-303.000000000000,
-330.000000000000,578.000000000000,
225.000000000000,412.000000000000,
222.000000000000,77.0000000000000,
-620.000000000000,-463.000000000000,
795.000000000000,-570.000000000000,
-168.000000000000,-325.000000000000,
-561.000000000000,340.000000000000,
339.000000000000,745.000000000000,
-988.000000000000,-521.000000000000,
202.000000000000,-67.0000000000000,
-210.000000000000,676.000000000000,
-501.000000000000,-504.000000000000,
1565.00000000000,207.000000000000,
506.000000000000,-2.00000000000000,
236.000000000000,317.000000000000,
-150.000000000000,1252.00000000000,
-1430.00000000000,131.000000000000,
-682.000000000000,48.0000000000000,
598.000000000000,421.000000000000,
-92.0000000000000,906.000000000000,
-295.000000000000,-12.0000000000000,
782.000000000000,324.000000000000,
-561.000000000000,-28.0000000000000,
-247.000000000000,-736.000000000000,
833.000000000000,265.000000000000,
177.000000000000,187.000000000000,
-177.000000000000,-432.000000000000,
12.0000000000000,-845.000000000000,
847.000000000000,-326.000000000000,
164.000000000000,293.000000000000,
-426.000000000000,686.000000000000,
14.0000000000000,-713.000000000000,
-20.0000000000000,-579.000000000000,
-9.00000000000000,712.000000000000,
-410.000000000000,-205.000000000000,
556.000000000000,-406.000000000000,
73.0000000000000,136.000000000000,
-465.000000000000,1017.00000000000,
417.000000000000,381.000000000000,
-843.000000000000,-449.000000000000,
-389.000000000000,44.0000000000000,
487.000000000000,179.000000000000,
-373.000000000000,-363.000000000000,
-527.000000000000,-1158.00000000000,
697.000000000000,-567.000000000000,
856.000000000000,188.000000000000,
-206.000000000000,1253.00000000000,
447.000000000000,276.000000000000,
193.000000000000,-329.000000000000,
-361.000000000000,1080.00000000000,
-190.000000000000,195.000000000000,
-255.000000000000,95.0000000000000,
207.000000000000,659.000000000000,
-51.0000000000000,-542.000000000000,
-456.000000000000,-463.000000000000,
-662.000000000000,124.000000000000,
120.000000000000,-1079.00000000000,
802.000000000000,-8.00000000000000,
659.000000000000,824.000000000000,
135.000000000000,-953.000000000000,
-631.000000000000,-218.000000000000,
128.000000000000,-256.000000000000,
248.000000000000,168.000000000000,
24.0000000000000,1251.00000000000,
-723.000000000000,388.000000000000,
-946.000000000000,-487.000000000000,
734.000000000000,-183.000000000000,
15.0000000000000,261.000000000000,
156.000000000000,-863.000000000000,
-302.000000000000,-183.000000000000,
-273.000000000000,-298.000000000000,
633.000000000000,-1004.00000000000,
-637.000000000000,-199.000000000000,
-178.000000000000,-479.000000000000,
746.000000000000,-103.000000000000,
1013.00000000000,-11.0000000000000,
615.000000000000,326.000000000000,
1034.00000000000,158.000000000000,
487.000000000000,108.000000000000,
-408.000000000000,1159.00000000000,
423.000000000000,188.000000000000,
625.000000000000,562.000000000000,
-781.000000000000,763.000000000000,
-292.000000000000,-763.000000000000,
886.000000000000,58.0000000000000,
-458.000000000000,346.000000000000,
-162.000000000000,534.000000000000,
530.000000000000,393.000000000000,
546.000000000000,201.000000000000,
226.000000000000,967.000000000000,
-346.000000000000,314.000000000000,
35.0000000000000,-28.0000000000000,
356.000000000000,-342.000000000000,
11.0000000000000,-597.000000000000,
-1048.00000000000,-456.000000000000,
112.000000000000,-295.000000000000,
1556.00000000000,326.000000000000,
-112.000000000000,984.000000000000,
-1052.00000000000,-129.000000000000,
-704.000000000000,-774.000000000000,
78.0000000000000,616.000000000000,
-15.0000000000000,722.000000000000,
-15.0000000000000,489.000000000000,
429.000000000000,-1106.00000000000,
143.000000000000,-447.000000000000,
893.000000000000,1058.00000000000,
7.00000000000000,62.0000000000000,
102.000000000000,351.000000000000,
894.000000000000,500.000000000000,
-434.000000000000,940.000000000000,
-246.000000000000,631.000000000000,
74.0000000000000,31.0000000000000,
-272.000000000000,155.000000000000,
-1087.00000000000,-76.0000000000000,
-586.000000000000,-618.000000000000,
-127.000000000000,-1540.00000000000,
886.000000000000,149.000000000000,
628.000000000000,-228.000000000000,
72.0000000000000,-9.00000000000000,
989.000000000000,518.000000000000,
360.000000000000,-1266.00000000000,
500.000000000000,625.000000000000,
-540.000000000000,263.000000000000,
533.000000000000,375.000000000000,
643.000000000000,264.000000000000,
-469.000000000000,-29.0000000000000,
734.000000000000,662.000000000000,
-507.000000000000,-181.000000000000,
74.0000000000000,519.000000000000,
-778.000000000000,-601.000000000000,
-483.000000000000,-503.000000000000,
1141.00000000000,35.0000000000000,
-431.000000000000,-165.000000000000,
591.000000000000,229.000000000000,
-32.0000000000000,647.000000000000,
-428.000000000000,157.000000000000,
1272.00000000000,-54.0000000000000,
-166.000000000000,243.000000000000,
-208.000000000000,-166.000000000000,
271.000000000000,187.000000000000,
358.000000000000,-130.000000000000,
-213.000000000000,1309.00000000000,
-460.000000000000,1191.00000000000,
-721.000000000000,689.000000000000,
-1075.00000000000,275.000000000000,
909.000000000000,-851.000000000000,
728.000000000000,-174.000000000000,
760.000000000000,-437.000000000000,
379.000000000000,790.000000000000,
-748.000000000000,120.000000000000,
-729.000000000000,-492.000000000000,
114.000000000000,875.000000000000,
-430.000000000000,-609.000000000000,
-976.000000000000,52.0000000000000,
1222.00000000000,-381.000000000000,
176.000000000000,363.000000000000,
-147.000000000000,1126.00000000000,
-1061.00000000000,-1003.00000000000,
137.000000000000,564.000000000000,
764.000000000000,-222.000000000000,
-1331.00000000000,402.000000000000,
-107.000000000000,433.000000000000,
-1151.00000000000,-450.000000000000,
594.000000000000,350.000000000000,
242.000000000000,120.000000000000,
-596.000000000000,-14.0000000000000,
419.000000000000,-1550.00000000000,
-932.000000000000,370.000000000000,
142.000000000000,189.000000000000,
-452.000000000000,-736.000000000000,
97.0000000000000,-706.000000000000,
833.000000000000,-1096.00000000000,
-6.00000000000000,-157.000000000000,
-199.000000000000,173.000000000000,
-547.000000000000,443.000000000000,
-68.0000000000000,-449.000000000000,
793.000000000000,-168.000000000000,
412.000000000000,508.000000000000,
-386.000000000000,47.0000000000000,
450.000000000000,515.000000000000,
336.000000000000,221.000000000000,
547.000000000000,-139.000000000000,
80.0000000000000,-308.000000000000,
-1028.00000000000,47.0000000000000,
-500.000000000000,335.000000000000,
-428.000000000000,182.000000000000,
1118.00000000000,544.000000000000,
369.000000000000,-792.000000000000,
-148.000000000000,-677.000000000000,
553.000000000000,-774.000000000000,
-455.000000000000,181.000000000000,
688.000000000000,781.000000000000,
-860.000000000000,-483.000000000000,
-775.000000000000,-242.000000000000,
774.000000000000,-850.000000000000,
656.000000000000,265.000000000000,
697.000000000000,-933.000000000000,
303.000000000000,-376.000000000000,
89.0000000000000,808.000000000000,
-1054.00000000000,-986.000000000000,
417.000000000000,279.000000000000,
318.000000000000,703.000000000000,
-416.000000000000,562.000000000000,
-435.000000000000,-504.000000000000,
-325.000000000000,-62.0000000000000,
1390.00000000000,242.000000000000,
-492.000000000000,79.0000000000000,
-150.000000000000,43.0000000000000,
-395.000000000000,-1122.00000000000,
-201.000000000000,342.000000000000,
1248.00000000000,308.000000000000,
-1065.00000000000,353.000000000000,
553.000000000000,-369.000000000000,
-179.000000000000,-315.000000000000,
-1145.00000000000,-94.0000000000000,
430.000000000000,-379.000000000000,
-956.000000000000,730.000000000000,
-797.000000000000,-899.000000000000,
24.0000000000000,-1002.00000000000,
-342.000000000000,-365.000000000000,
535.000000000000,-230.000000000000,
775.000000000000,-399.000000000000,
-140.000000000000,-979.000000000000,
718.000000000000,184.000000000000,
-866.000000000000,-187.000000000000,
-1044.00000000000,-158.000000000000,
792.000000000000,-359.000000000000,
-303.000000000000,-953.000000000000,
746.000000000000,615.000000000000,
91.0000000000000,414.000000000000,
-561.000000000000,118.000000000000,
644.000000000000,-176.000000000000,
-483.000000000000,-601.000000000000,
-519.000000000000,-34.0000000000000,
-391.000000000000,996.000000000000,
-505.000000000000,862.000000000000,
35.0000000000000,16.0000000000000,
345.000000000000,-591.000000000000,
418.000000000000,-280.000000000000,
921.000000000000,567.000000000000,
1070.00000000000,-54.0000000000000,
-763.000000000000,368.000000000000,
-559.000000000000,-620.000000000000,
-329.000000000000,-668.000000000000,
-952.000000000000,455.000000000000,
-297.000000000000,-21.0000000000000,
-755.000000000000,729.000000000000,
221.000000000000,644.000000000000,
715.000000000000,-87.0000000000000,
-159.000000000000,-788.000000000000,
-771.000000000000,-569.000000000000,
9.00000000000000,-319.000000000000,
-269.000000000000,-779.000000000000,
-529.000000000000,409.000000000000,
181.000000000000,-322.000000000000,
-1116.00000000000,-23.0000000000000,
904.000000000000,40.0000000000000,
656.000000000000,-72.0000000000000,
102.000000000000,1214.00000000000,
489.000000000000,-452.000000000000,
-160.000000000000,934.000000000000,
186.000000000000,40.0000000000000,
-1471.00000000000,-687.000000000000,
-721.000000000000,210.000000000000,
-35.0000000000000,-1055.00000000000,
751.000000000000,392.000000000000,
458.000000000000,-213.000000000000,
797.000000000000,262.000000000000,
457.000000000000,690.000000000000,
-1592.00000000000,153.000000000000,
-601.000000000000,-497.000000000000,
-1380.00000000000,-619.000000000000,
182.000000000000,617.000000000000,
648.000000000000,303.000000000000,
-680.000000000000,1239.00000000000,
-256.000000000000,-727.000000000000,
24.0000000000000,-780.000000000000,
819.000000000000,639.000000000000,
-767.000000000000,-888.000000000000,
-78.0000000000000,-963.000000000000,
999.000000000000,-224.000000000000,
-296.000000000000,522.000000000000,
-409.000000000000,-1150.00000000000,
304.000000000000,-662.000000000000,
-31.0000000000000,589.000000000000,
-761.000000000000,-268.000000000000,
674.000000000000,436.000000000000,
-327.000000000000,1119.00000000000,
-250.000000000000,851.000000000000,
1049.00000000000,114.000000000000,
-365.000000000000,124.000000000000,
992.000000000000,-631.000000000000,
744.000000000000,-17.0000000000000,
801.000000000000,-107.000000000000,
323.000000000000,46.0000000000000,
-1267.00000000000,-9.00000000000000,
957.000000000000,-776.000000000000,
-89.0000000000000,1154.00000000000,
-1000.00000000000,9.00000000000000,
-351.000000000000,-768.000000000000,
82.0000000000000,-535.000000000000,
449.000000000000,-792.000000000000,
-54.0000000000000,-488.000000000000,
387.000000000000,-551.000000000000,
488.000000000000,699.000000000000,
-197.000000000000,-111.000000000000,
354.000000000000,-381.000000000000,
1467.00000000000,592.000000000000,
-427.000000000000,-66.0000000000000,
-876.000000000000,103.000000000000,
-600.000000000000,-752.000000000000,
-412.000000000000,-348.000000000000,
407.000000000000,-29.0000000000000,
-53.0000000000000,-93.0000000000000,
472.000000000000,890.000000000000,
-429.000000000000,-681.000000000000,
-3.00000000000000,-900.000000000000,
481.000000000000,-912.000000000000,
28.0000000000000,-1164.00000000000,
1431.00000000000,-397.000000000000,
457.000000000000,368.000000000000,
-948.000000000000,35.0000000000000,
-431.000000000000,-161.000000000000,
1190.00000000000,292.000000000000,
398.000000000000,-147.000000000000,
-877.000000000000,109.000000000000,
643.000000000000,-468.000000000000,
-487.000000000000,-195.000000000000,
-1191.00000000000,150.000000000000,
495.000000000000,-238.000000000000,
-158.000000000000,381.000000000000,
-334.000000000000,366.000000000000,
1295.00000000000,483.000000000000,
295.000000000000,-77.0000000000000,
97.0000000000000,-1020.00000000000,
1151.00000000000,73.0000000000000,
67.0000000000000,752.000000000000,
-374.000000000000,197.000000000000,
-353.000000000000,49.0000000000000,
-833.000000000000,311.000000000000,
-575.000000000000,296.000000000000,
406.000000000000,-639.000000000000,
427.000000000000,-347.000000000000,
110.000000000000,798.000000000000,
-126.000000000000,371.000000000000,
-781.000000000000,417.000000000000,
-807.000000000000,708.000000000000,
103.000000000000,116.000000000000,
376.000000000000,752.000000000000,
986.000000000000,375.000000000000,
456.000000000000,-503.000000000000,
141.000000000000,-343.000000000000,
-270.000000000000,-1020.00000000000,
-505.000000000000,-70.0000000000000,
308.000000000000,-375.000000000000,
506.000000000000,173.000000000000,
447.000000000000,1228.00000000000,
-822.000000000000,1046.00000000000,
241.000000000000,737.000000000000,
-167.000000000000,-427.000000000000,
-1278.00000000000,-266.000000000000,
330.000000000000,-1497.00000000000,
-369.000000000000,-891.000000000000,
-468.000000000000,547.000000000000,
-342.000000000000,186.000000000000,
-524.000000000000,601.000000000000,
-132.000000000000,700.000000000000,
773.000000000000,546.000000000000,
555.000000000000,691.000000000000,
-74.0000000000000,587.000000000000,
750.000000000000,-401.000000000000,
-403.000000000000,459.000000000000,
10.0000000000000,-386.000000000000,
197.000000000000,-1210.00000000000,
-464.000000000000,1118.00000000000,
-85.0000000000000,-385.000000000000,
-249.000000000000,-97.0000000000000,
-203.000000000000,294.000000000000,
-1554.00000000000,-682.000000000000,
173.000000000000,-862.000000000000,
699.000000000000,-912.000000000000,
541.000000000000,1031.00000000000,
1102.00000000000,-167.000000000000,
-136.000000000000,-63.0000000000000,
-76.0000000000000,61.0000000000000,
-1050.00000000000,-774.000000000000,
-496.000000000000,154.000000000000,
-139.000000000000,241.000000000000,
339.000000000000,197.000000000000,
492.000000000000,-532.000000000000,
-5.00000000000000,-107.000000000000,
657.000000000000,-186.000000000000,
-832.000000000000,807.000000000000,
259.000000000000,39.0000000000000,
431.000000000000,-920.000000000000,
-65.0000000000000,1038.00000000000,
581.000000000000,-768.000000000000,
565.000000000000,555.000000000000,
412.000000000000,555.000000000000,
64.0000000000000,-1032.00000000000,
466.000000000000,521.000000000000,
165.000000000000,-329.000000000000,
237.000000000000,518.000000000000,
-1072.00000000000,-516.000000000000,
252.000000000000,-121.000000000000,
272.000000000000,623.000000000000,
-306.000000000000,-638.000000000000,
1254.00000000000,-66.0000000000000,
42.0000000000000,-1135.00000000000,
825.000000000000,-230.000000000000,
-300.000000000000,399.000000000000,
-1240.00000000000,-713.000000000000,
596.000000000000,-472.000000000000,
546.000000000000,41.0000000000000,
152.000000000000,2.00000000000000,
-344.000000000000,1188.00000000000,
152.000000000000,1302.00000000000,
158.000000000000,-806.000000000000,
44.0000000000000,651.000000000000,
212.000000000000,564.000000000000,
-271.000000000000,949.000000000000,
-268.000000000000,869.000000000000,
-1436.00000000000,-805.000000000000,
-36.0000000000000,-351.000000000000,
-51.0000000000000,-1429.00000000000,
-64.0000000000000,308.000000000000,
377.000000000000,-415.000000000000,
-301.000000000000,-447.000000000000,
668.000000000000,556.000000000000,
-378.000000000000,-1191.00000000000,
763.000000000000,91.0000000000000,
-763.000000000000,-207.000000000000,
-1072.00000000000,-407.000000000000,
633.000000000000,-1334.00000000000,
-615.000000000000,200.000000000000,
1282.00000000000,792.000000000000,
871.000000000000,184.000000000000,
458.000000000000,1271.00000000000,
232.000000000000,-561.000000000000,
158.000000000000,-956.000000000000,
1288.00000000000,-82.0000000000000,
-393.000000000000,266.000000000000,
-519.000000000000,-828.000000000000,
-187.000000000000,-330.000000000000,
682.000000000000,406.000000000000,
539.000000000000,338.000000000000,
-788.000000000000,331.000000000000,
-289.000000000000,-1330.00000000000,
-627.000000000000,-222.000000000000,
-493.000000000000,645.000000000000,
333.000000000000,231.000000000000,
852.000000000000,-74.0000000000000,
-177.000000000000,105.000000000000,
-523.000000000000,217.000000000000,
-538.000000000000,-1122.00000000000,
-195.000000000000,134.000000000000,
597.000000000000,-302.000000000000,
-731.000000000000,-795.000000000000,
-19.0000000000000,745.000000000000,
-1047.00000000000,-214.000000000000,
-694.000000000000,-321.000000000000,
530.000000000000,-58.0000000000000,
-575.000000000000,535.000000000000,
489.000000000000,-872.000000000000,
285.000000000000,-1069.00000000000,
389.000000000000,574.000000000000,
-7.00000000000000,106.000000000000,
-214.000000000000,124.000000000000,
151.000000000000,-1213.00000000000,
736.000000000000,-438.000000000000,
1400.00000000000,535.000000000000,
-835.000000000000,667.000000000000,
-108.000000000000,190.000000000000,
572.000000000000,-312.000000000000,
763.000000000000,1018.00000000000,
474.000000000000,-262.000000000000,
-302.000000000000,-595.000000000000,
653.000000000000,-353.000000000000,
560.000000000000,321.000000000000,
372.000000000000,416.000000000000,
-845.000000000000,302.000000000000,
-166.000000000000,1212.00000000000,
-381.000000000000,-271.000000000000,
-1401.00000000000,53.0000000000000,
-216.000000000000,-487.000000000000,
230.000000000000,-856.000000000000,
572.000000000000,678.000000000000,
713.000000000000,31.0000000000000,
434.000000000000,668.000000000000,
-59.0000000000000,1017.00000000000,
122.000000000000,-427.000000000000,
193.000000000000,-281.000000000000,
-26.0000000000000,319.000000000000,
-464.000000000000,30.0000000000000,
-295.000000000000,-148.000000000000,
561.000000000000,-312.000000000000,
-27.0000000000000,-700.000000000000,
295.000000000000,490.000000000000,
146.000000000000,864.000000000000,
222.000000000000,966.000000000000,
422.000000000000,255.000000000000,
-1209.00000000000,-272.000000000000,
55.0000000000000,334.000000000000,
-49.0000000000000,-960.000000000000,
-1152.00000000000,-487.000000000000,
-233.000000000000,-546.000000000000,
-369.000000000000,33.0000000000000,
-393.000000000000,382.000000000000,
-533.000000000000,-751.000000000000,
972.000000000000,-172.000000000000,
595.000000000000,-758.000000000000,
138.000000000000,-356.000000000000,
1323.00000000000,-20.0000000000000,
835.000000000000,562.000000000000,
612.000000000000,-105.000000000000,
-336.000000000000,-211.000000000000,
-36.0000000000000,1384.00000000000,
71.0000000000000,207.000000000000,
113.000000000000,-110.000000000000,
-35.0000000000000,631.000000000000,
-506.000000000000,906.000000000000,
360.000000000000,-417.000000000000,
-150.000000000000,331.000000000000,
-685.000000000000,1437.00000000000,
-1185.00000000000,-927.000000000000,
-67.0000000000000,204.000000000000,
853.000000000000,1138.00000000000,
-347.000000000000,-483.000000000000,
-110.000000000000,-290.000000000000,
1012.00000000000,263.000000000000,
171.000000000000,298.000000000000,
-816.000000000000,1034.00000000000,
80.0000000000000,452.000000000000,
311.000000000000,99.0000000000000,
90.0000000000000,357.000000000000,
677.000000000000,309.000000000000,
-262.000000000000,688.000000000000,
-1180.00000000000,523.000000000000,
-96.0000000000000,224.000000000000,
-38.0000000000000,-143.000000000000,
-437.000000000000,-898.000000000000,
323.000000000000,93.0000000000000,
156.000000000000,-465.000000000000,
341.000000000000,-447.000000000000,
738.000000000000,1049.00000000000,
-1020.00000000000,-773.000000000000,
-293.000000000000,-282.000000000000,
-378.000000000000,855.000000000000,
-704.000000000000,1193.00000000000,
-159.000000000000,-89.0000000000000,
-799.000000000000,-654.000000000000,
1402.00000000000,359.000000000000,
183.000000000000,77.0000000000000,
-924.000000000000,561.000000000000,
-369.000000000000,-261.000000000000,
-737.000000000000,756.000000000000,
378.000000000000,579.000000000000,
-358.000000000000,-482.000000000000,
-288.000000000000,557.000000000000,
198.000000000000,355.000000000000,
53.0000000000000,-801.000000000000,
55.0000000000000,-122.000000000000,
-185.000000000000,1000.00000000000,
509.000000000000,-786.000000000000,
176.000000000000,-887.000000000000,
-315.000000000000,-28.0000000000000,
258.000000000000,-41.0000000000000,
999.000000000000,-130.000000000000,
577.000000000000,-595.000000000000,
556.000000000000,40.0000000000000,
330.000000000000,-512.000000000000,
251.000000000000,-435.000000000000,
806.000000000000,222.000000000000,
-258.000000000000,-345.000000000000,
42.0000000000000,204.000000000000,
-265.000000000000,-648.000000000000,
30.0000000000000,-861.000000000000,
1491.00000000000,107.000000000000,
-301.000000000000,410.000000000000,
-980.000000000000,-343.000000000000,
239.000000000000,-335.000000000000,
1135.00000000000,391.000000000000,
263.000000000000,-216.000000000000,
-477.000000000000,472.000000000000,
-188.000000000000,695.000000000000,
15.0000000000000,773.000000000000,
311.000000000000,341.000000000000,
-1153.00000000000,413.000000000000,
125.000000000000,-48.0000000000000,
157.000000000000,-722.000000000000,
-581.000000000000,356.000000000000,
1241.00000000000,-241.000000000000,
-577.000000000000,838.000000000000,
-300.000000000000,734.000000000000,
-675.000000000000,-102.000000000000,
-738.000000000000,557.000000000000,
275.000000000000,379.000000000000,
178.000000000000,-580.000000000000,
929.000000000000,-630.000000000000,
-371.000000000000,719.000000000000,
-132.000000000000,-1442.00000000000,
1025.00000000000,-332.000000000000,
895.000000000000,940.000000000000,
-579.000000000000,-868.000000000000,
882.000000000000,405.000000000000,
649.000000000000,-78.0000000000000,
-1078.00000000000,1033.00000000000,
581.000000000000,396.000000000000,
-663.000000000000,-546.000000000000,
782.000000000000,408.000000000000,
253.000000000000,-1181.00000000000,
-653.000000000000,-246.000000000000,
183.000000000000,246.000000000000,
-817.000000000000,1518.00000000000,
161.000000000000,334.000000000000,
-309.000000000000,-324.000000000000,
1326.00000000000,290.000000000000,
-124.000000000000,-676.000000000000,
-673.000000000000,28.0000000000000,
928.000000000000,-523.000000000000,
-1004.00000000000,439.000000000000,
-572.000000000000,-159.000000000000,
-624.000000000000,257.000000000000,
-655.000000000000,1123.00000000000,
-882.000000000000,-187.000000000000,
-1120.00000000000,105.000000000000,
-80.0000000000000,98.0000000000000,
258.000000000000,-101.000000000000,
107.000000000000,230.000000000000,
-318.000000000000,327.000000000000,
589.000000000000,-363.000000000000,
-182.000000000000,956.000000000000,
-577.000000000000,404.000000000000,
-313.000000000000,-538.000000000000,
-48.0000000000000,989.000000000000,
544.000000000000,-613.000000000000,
-761.000000000000,238.000000000000,
683.000000000000,683.000000000000,
-293.000000000000,-963.000000000000,
-1166.00000000000,65.0000000000000,
678.000000000000,-419.000000000000,
-276.000000000000,-121.000000000000,
-676.000000000000,-445.000000000000,
505.000000000000,-410.000000000000,
1048.00000000000,-172.000000000000,
-156.000000000000,-284.000000000000,
603.000000000000,1071.00000000000,
234.000000000000,-173.000000000000,
534.000000000000,73.0000000000000,
788.000000000000,-212.000000000000,
-469.000000000000,-149.000000000000,
397.000000000000,-76.0000000000000,
297.000000000000,-1049.00000000000,
1120.00000000000,612.000000000000,
147.000000000000,252.000000000000,
-349.000000000000,357.000000000000,
-427.000000000000,-492.000000000000,
-1305.00000000000,-411.000000000000,
751.000000000000,-327.000000000000,
441.000000000000,-83.0000000000000,
855.000000000000,903.000000000000,
15.0000000000000,-754.000000000000,
-591.000000000000,1068.00000000000,
-186.000000000000,439.000000000000,
-1039.00000000000,-270.000000000000,
601.000000000000,292.000000000000,
-288.000000000000,-262.000000000000,
-606.000000000000,550.000000000000,
346.000000000000,205.000000000000,
312.000000000000,495.000000000000,
-904.000000000000,139.000000000000,
-640.000000000000,670.000000000000,
622.000000000000,350.000000000000,
-373.000000000000,656.000000000000,
760.000000000000,833.000000000000,
21.0000000000000,-1051.00000000000,
505.000000000000,562.000000000000,
858.000000000000,528.000000000000,
-899.000000000000,799.000000000000,
-114.000000000000,54.0000000000000,
-162.000000000000,-1430.00000000000,
331.000000000000,-541.000000000000,
-37.0000000000000,-1153.00000000000,
-166.000000000000,262.000000000000,
-293.000000000000,-678.000000000000,
-206.000000000000,-265.000000000000,
-360.000000000000,242.000000000000,
-383.000000000000,-819.000000000000,
529.000000000000,575.000000000000,
-1000.00000000000,-492.000000000000,
145.000000000000,-495.000000000000,
312.000000000000,-607.000000000000,
-112.000000000000,-569.000000000000,
1268.00000000000,210.000000000000,
422.000000000000,-173.000000000000,
1146.00000000000,378.000000000000,
835.000000000000,706.000000000000,
-1080.00000000000,55.0000000000000,
-688.000000000000,64.0000000000000,
48.0000000000000,808.000000000000,
406.000000000000,-543.000000000000,
1164.00000000000,148.000000000000,
-35.0000000000000,1431.00000000000,
-420.000000000000,2.00000000000000,
664.000000000000,471.000000000000,
-918.000000000000,1249.00000000000,
-778.000000000000,897.000000000000,
-229.000000000000,-111.000000000000,
-791.000000000000,-498.000000000000,
627.000000000000,-857.000000000000,
172.000000000000,-1283.00000000000,
-156.000000000000,280.000000000000,
-736.000000000000,-333.000000000000,
-1168.00000000000,-541.000000000000,
93.0000000000000,-1151.00000000000,
317.000000000000,-623.000000000000,
455.000000000000,1494.00000000000,
-401.000000000000,443.000000000000,
-247.000000000000,69.0000000000000,
168.000000000000,290.000000000000,
39.0000000000000,-256.000000000000,
-675.000000000000,-1004.00000000000,
-902.000000000000,228.000000000000,
1016.00000000000,116.000000000000,
258.000000000000,201.000000000000,
-453.000000000000,899.000000000000,
-684.000000000000,-560.000000000000,
-547.000000000000,705.000000000000,
-683.000000000000,35.0000000000000,
-695.000000000000,68.0000000000000,
672.000000000000,92.0000000000000,
-212.000000000000,-1058.00000000000,
275.000000000000,1134.00000000000,
436.000000000000,-353.000000000000,
196.000000000000,-144.000000000000,
222.000000000000,-20.0000000000000,
-15.0000000000000,45.0000000000000,
64.0000000000000,1227.00000000000,
104.000000000000,-19.0000000000000,
461.000000000000,479.000000000000,
-1325.00000000000,-473.000000000000,
112.000000000000,-158.000000000000,
1152.00000000000,-426.000000000000,
475.000000000000,-209.000000000000,
303.000000000000,940.000000000000,
-1345.00000000000,344.000000000000,
-54.0000000000000,-33.0000000000000,
-446.000000000000,-436.000000000000,
-293.000000000000,1115.00000000000,
757.000000000000,-476.000000000000,
7.00000000000000,284.000000000000,
445.000000000000,1295.00000000000,
-170.000000000000,-244.000000000000,
365.000000000000,-437.000000000000,
-279.000000000000,-894.000000000000,
-303.000000000000,-250.000000000000,
616.000000000000,37.0000000000000,
-417.000000000000,1206.00000000000,
-301.000000000000,674.000000000000,
-546.000000000000,381.000000000000,
513.000000000000,456.000000000000,
536.000000000000,-932.000000000000,
195.000000000000,-411.000000000000,
123.000000000000,469.000000000000,
-964.000000000000,-110.000000000000,
168.000000000000,-938.000000000000,
250.000000000000,112.000000000000,
9.00000000000000,-8.00000000000000,
-726.000000000000,290.000000000000,
-450.000000000000,348.000000000000,
1070.00000000000,-853.000000000000,
548.000000000000,474.000000000000,
850.000000000000,556.000000000000,
128.000000000000,335.000000000000,
-601.000000000000,478.000000000000,
-106.000000000000,113.000000000000,
-74.0000000000000,42.0000000000000,
-795.000000000000,102.000000000000,
-43.0000000000000,801.000000000000,
818.000000000000,84.0000000000000,
-1039.00000000000,-539.000000000000,
-895.000000000000,-89.0000000000000,
153.000000000000,273.000000000000,
322.000000000000,99.0000000000000,
665.000000000000,370.000000000000,
472.000000000000,248.000000000000,
382.000000000000,-1379.00000000000,
805.000000000000,-297.000000000000,
1527.00000000000,-110.000000000000,
-442.000000000000,-543.000000000000,
297.000000000000,525.000000000000,
912.000000000000,-153.000000000000,
-1348.00000000000,562.000000000000,
-775.000000000000,-559.000000000000,
-744.000000000000,-365.000000000000,
5.00000000000000,961.000000000000,
285.000000000000,-899.000000000000,
403.000000000000,-421.000000000000,
76.0000000000000,749.000000000000,
-908.000000000000,-169.000000000000,
-249.000000000000,180.000000000000,
-805.000000000000,770.000000000000,
-506.000000000000,-625.000000000000,
-300.000000000000,-421.000000000000,
-732.000000000000,-493.000000000000,
-465.000000000000,140.000000000000,
-353.000000000000,1190.00000000000,
-382.000000000000,500.000000000000,
-931.000000000000,665.000000000000,
-291.000000000000,-447.000000000000,
606.000000000000,-953.000000000000,
324.000000000000,-156.000000000000,
-480.000000000000,-830.000000000000,
622.000000000000,-463.000000000000,
1122.00000000000,-44.0000000000000,
-648.000000000000,705.000000000000,
7.00000000000000,1210.00000000000,
-833.000000000000,627.000000000000,
-1080.00000000000,-126.000000000000,
610.000000000000,-300.000000000000,
783.000000000000,40.0000000000000,
1039.00000000000,440.000000000000,
610.000000000000,254.000000000000,
394.000000000000,-318.000000000000,
-374.000000000000,365.000000000000,
-414.000000000000,-169.000000000000,
12.0000000000000,-61.0000000000000,
-193.000000000000,864.000000000000,
-592.000000000000,852.000000000000,
-1090.00000000000,557.000000000000,
318.000000000000,-1075.00000000000,
-562.000000000000,-180.000000000000,
-174.000000000000,-837.000000000000,
415.000000000000,-1526.00000000000,
-542.000000000000,805.000000000000,
-56.0000000000000,-372.000000000000,
337.000000000000,320.000000000000,
962.000000000000,538.000000000000,
136.000000000000,-817.000000000000,
242.000000000000,-12.0000000000000,
-285.000000000000,-555.000000000000,
374.000000000000,7.00000000000000,
236.000000000000,-318.000000000000,
-460.000000000000,376.000000000000,
728.000000000000,213.000000000000,
-929.000000000000,-404.000000000000,
-581.000000000000,145.000000000000,
-18.0000000000000,195.000000000000,
433.000000000000,679.000000000000,
624.000000000000,-149.000000000000,
-480.000000000000,951.000000000000,
-956.000000000000,-34.0000000000000,
-729.000000000000,-1021.00000000000,
560.000000000000,-502.000000000000,
-549.000000000000,-1025.00000000000,
132.000000000000,998.000000000000,
273.000000000000,-384.000000000000,
-253.000000000000,-525.000000000000,
523.000000000000,-538.000000000000,
28.0000000000000,-627.000000000000,
295.000000000000,1123.00000000000,
-307.000000000000,160.000000000000,
-258.000000000000,617.000000000000,
-86.0000000000000,335.000000000000,
404.000000000000,-291.000000000000,
1051.00000000000,53.0000000000000,
915.000000000000,108.000000000000,
443.000000000000,748.000000000000,
-192.000000000000,799.000000000000,
115.000000000000,-122.000000000000,
-607.000000000000,152.000000000000,
-571.000000000000,780.000000000000,
209.000000000000,233.000000000000,
-666.000000000000,898.000000000000,
-808.000000000000,1046.00000000000,
-125.000000000000,-247.000000000000,
-40.0000000000000,-951.000000000000,
-146.000000000000,-334.000000000000,
-56.0000000000000,774.000000000000,
-192.000000000000,608.000000000000,
-341.000000000000,1029.00000000000,
55.0000000000000,-418.000000000000,
436.000000000000,-1402.00000000000,
811.000000000000,-3.00000000000000,
-70.0000000000000,-1082.00000000000,
-138.000000000000,335.000000000000,
-368.000000000000,255.000000000000,
-12.0000000000000,-665.000000000000,
399.000000000000,567.000000000000,
63.0000000000000,-83.0000000000000,
755.000000000000,519.000000000000,
-570.000000000000,-248.000000000000,
-545.000000000000,-193.000000000000,
-172.000000000000,-450.000000000000,
-448.000000000000,-1123.00000000000,
-53.0000000000000,286.000000000000,
100.000000000000,659.000000000000,
497.000000000000,420.000000000000,
-588.000000000000,302.000000000000,
-774.000000000000,-570.000000000000,
200.000000000000,-1045.00000000000,
-579.000000000000,107.000000000000,
-552.000000000000,-200.000000000000,
-347.000000000000,-612.000000000000,
-217.000000000000,281.000000000000,
99.0000000000000,126.000000000000,
285.000000000000,-146.000000000000,
932.000000000000,-396.000000000000,
1148.00000000000,471.000000000000,
911.000000000000,112.000000000000,
530.000000000000,421.000000000000,
-247.000000000000,437.000000000000,
-809.000000000000,-1171.00000000000,
200.000000000000,445.000000000000,
-707.000000000000,-359.000000000000,
-349.000000000000,-451.000000000000,
-28.0000000000000,702.000000000000,
-1657.00000000000,204.000000000000,
722.000000000000,29.0000000000000,
-53.0000000000000,-1139.00000000000,
-419.000000000000,-555.000000000000,
1045.00000000000,-1356.00000000000,
528.000000000000,-672.000000000000,
777.000000000000,546.000000000000,
-1182.00000000000,633.000000000000,
324.000000000000,42.0000000000000,
629.000000000000,-13.0000000000000,
-484.000000000000,1065.00000000000,
926.000000000000,130.000000000000,
464.000000000000,253.000000000000,
-26.0000000000000,-1396.00000000000,
-70.0000000000000,-108.000000000000,
177.000000000000,839.000000000000,
-1136.00000000000,-652.000000000000,
74.0000000000000,805.000000000000,
-581.000000000000,-224.000000000000,
-1179.00000000000,-949.000000000000,
1063.00000000000,-372.000000000000,
-985.000000000000,-62.0000000000000,
422.000000000000,-591.000000000000,
287.000000000000,262.000000000000,
-833.000000000000,357.000000000000,
723.000000000000,-735.000000000000,
-374.000000000000,1063.00000000000,
-232.000000000000,748.000000000000,
-283.000000000000,847.000000000000,
-463.000000000000,1160.00000000000,
476.000000000000,78.0000000000000,
-65.0000000000000,37.0000000000000,
-338.000000000000,-841.000000000000,
673.000000000000,-999.000000000000,
-587.000000000000,-628.000000000000,
-588.000000000000,-4.00000000000000,
-581.000000000000,52.0000000000000,
-1350.00000000000,-840.000000000000,
371.000000000000,785.000000000000,
-186.000000000000,744.000000000000,
-932.000000000000,-695.000000000000,
2.00000000000000,152.000000000000,
705.000000000000,402.000000000000,
937.000000000000,110.000000000000,
919.000000000000,492.000000000000,
637.000000000000,213.000000000000,
246.000000000000,26.0000000000000,
311.000000000000,774.000000000000,
21.0000000000000,523.000000000000,
-227.000000000000,289.000000000000,
-592.000000000000,340.000000000000,
-186.000000000000,367.000000000000,
-76.0000000000000,926.000000000000,
-419.000000000000,92.0000000000000,
-235.000000000000,687.000000000000,
-517.000000000000,1157.00000000000,
-57.0000000000000,34.0000000000000,
-70.0000000000000,-129.000000000000,
111.000000000000,-955.000000000000,
135.000000000000,-443.000000000000,
14.0000000000000,187.000000000000,
438.000000000000,228.000000000000,
-509.000000000000,417.000000000000,
-70.0000000000000,-297.000000000000,
526.000000000000,134.000000000000,
-578.000000000000,711.000000000000,
-24.0000000000000,-681.000000000000,
238.000000000000,-461.000000000000,
367.000000000000,604.000000000000,
550.000000000000,-166.000000000000,
-605.000000000000,415.000000000000,
-316.000000000000,-838.000000000000,
-584.000000000000,-627.000000000000,
268.000000000000,550.000000000000,
-68.0000000000000,-276.000000000000,
-314.000000000000,491.000000000000,
413.000000000000,-55.0000000000000,
-840.000000000000,-595.000000000000,
173.000000000000,-342.000000000000,
-241.000000000000,141.000000000000,
153.000000000000,-520.000000000000,
762.000000000000,-1065.00000000000,
-347.000000000000,388.000000000000,
-304.000000000000,526.000000000000,
-226.000000000000,118.000000000000,
-290.000000000000,-452.000000000000,
-632.000000000000,-668.000000000000,
-103.000000000000,-467.000000000000,
306.000000000000,-305.000000000000,
-694.000000000000,-156.000000000000,
-666.000000000000,-1075.00000000000,
778.000000000000,-95.0000000000000,
-10.0000000000000,144.000000000000,
30.0000000000000,-1102.00000000000,
1132.00000000000,90.0000000000000,
-31.0000000000000,686.000000000000,
125.000000000000,13.0000000000000,
113.000000000000,273.000000000000,
-478.000000000000,111.000000000000,
275.000000000000,-894.000000000000,
87.0000000000000,-143.000000000000,
32.0000000000000,587.000000000000,
-611.000000000000,706.000000000000,
163.000000000000,355.000000000000,
307.000000000000,-193.000000000000,
-441.000000000000,728.000000000000,
1045.00000000000,172.000000000000,
613.000000000000,243.000000000000,
876.000000000000,573.000000000000,
-15.0000000000000,505.000000000000,
-509.000000000000,224.000000000000,
586.000000000000,-372.000000000000,
71.0000000000000,1388.00000000000,
-982.000000000000,54.0000000000000,
-1550.00000000000,-563.000000000000,
502.000000000000,145.000000000000,
-87.0000000000000,-218.000000000000,
254.000000000000,331.000000000000,
134.000000000000,416.000000000000,
-853.000000000000,395.000000000000,
454.000000000000,225.000000000000,
-870.000000000000,788.000000000000,
-990.000000000000,-994.000000000000,
190.000000000000,-903.000000000000,
1027.00000000000,890.000000000000,
101.000000000000,-483.000000000000,
-419.000000000000,408.000000000000,
-243.000000000000,956.000000000000,
-1247.00000000000,35.0000000000000,
-700.000000000000,-877.000000000000,
-570.000000000000,-825.000000000000,
513.000000000000,-742.000000000000,
29.0000000000000,-1103.00000000000,
-433.000000000000,588.000000000000,
509.000000000000,-313.000000000000,
739.000000000000,524.000000000000,
571.000000000000,778.000000000000,
-321.000000000000,-395.000000000000,
887.000000000000,473.000000000000,
310.000000000000,-819.000000000000,
593.000000000000,327.000000000000,
922.000000000000,803.000000000000,
-483.000000000000,756.000000000000,
-91.0000000000000,545.000000000000,
213.000000000000,22.0000000000000,
332.000000000000,738.000000000000,
-379.000000000000,276.000000000000,
-466.000000000000,-325.000000000000,
-270.000000000000,-1036.00000000000,
-250.000000000000,-23.0000000000000,
388.000000000000,1087.00000000000,
389.000000000000,101.000000000000,
121.000000000000,334.000000000000,
-451.000000000000,769.000000000000,
-508.000000000000,-831.000000000000,
564.000000000000,-541.000000000000,
801.000000000000,-516.000000000000,
813.000000000000,-490.000000000000,
50.0000000000000,1224.00000000000,
-844.000000000000,-182.000000000000,
-762.000000000000,-45.0000000000000,
-73.0000000000000,1032.00000000000,
387.000000000000,-84.0000000000000,
15.0000000000000,244.000000000000,
648.000000000000,603.000000000000,
335.000000000000,-347.000000000000,
320.000000000000,-713.000000000000,
68.0000000000000,28.0000000000000,
266.000000000000,357.000000000000,
1235.00000000000,418.000000000000,
30.0000000000000,264.000000000000,
-996.000000000000,-333.000000000000,
-911.000000000000,868.000000000000,
458.000000000000,-15.0000000000000,
674.000000000000,-855.000000000000,
953.000000000000,890.000000000000,
76.0000000000000,564.000000000000,
-1174.00000000000,-94.0000000000000,
719.000000000000,-507.000000000000,
84.0000000000000,53.0000000000000,
-244.000000000000,127.000000000000,
-572.000000000000,-56.0000000000000,
-491.000000000000,451.000000000000,
-910.000000000000,-684.000000000000,
-974.000000000000,-1098.00000000000,
1374.00000000000,-493.000000000000,
308.000000000000,1040.00000000000,
-120.000000000000,696.000000000000,
-238.000000000000,726.000000000000,
-483.000000000000,824.000000000000,
14.0000000000000,-941.000000000000,
583.000000000000,-175.000000000000,
102.000000000000,-753.000000000000,
-649.000000000000,-604.000000000000,
700.000000000000,-2.00000000000000,
158.000000000000,-109.000000000000,
366.000000000000,436.000000000000,
62.0000000000000,-963.000000000000,
636.000000000000,671.000000000000,
847.000000000000,85.0000000000000,
-770.000000000000,-832.000000000000,
577.000000000000,153.000000000000,
-309.000000000000,-301.000000000000,
-254.000000000000,-291.000000000000,
446.000000000000,-740.000000000000,
950.000000000000,-255.000000000000,
781.000000000000,-231.000000000000,
-1010.00000000000,641.000000000000,
123.000000000000,-844.000000000000,
47.0000000000000,-820.000000000000,
1062.00000000000,699.000000000000,
539.000000000000,-709.000000000000,
-218.000000000000,-684.000000000000,
510.000000000000,111.000000000000,
-754.000000000000,-112.000000000000,
759.000000000000,-385.000000000000,
-299.000000000000,920.000000000000,
-404.000000000000,-686.000000000000,
1082.00000000000,-1301.00000000000,
718.000000000000,1112.00000000000,
677.000000000000,346.000000000000,
412.000000000000,797.000000000000,
889.000000000000,555.000000000000,
-185.000000000000,1052.00000000000,
-707.000000000000,831.000000000000,
-397.000000000000,-1357.00000000000,
1361.00000000000,600.000000000000,
758.000000000000,-397.000000000000,
7.00000000000000,-1047.00000000000,
1187.00000000000,-912.000000000000,
-131.000000000000,-459.000000000000,
610.000000000000,222.000000000000,
173.000000000000,-1089.00000000000,
764.000000000000,923.000000000000,
-393.000000000000,525.000000000000,
-1567.00000000000,-659.000000000000,
1367.00000000000,111.000000000000,
-133.000000000000,170.000000000000,
291.000000000000,-198.000000000000,
448.000000000000,688.000000000000,
-950.000000000000,-5.00000000000000,
222.000000000000,-964.000000000000,
-671.000000000000,943.000000000000,
-266.000000000000,334.000000000000,
234.000000000000,488.000000000000,
-779.000000000000,37.0000000000000,
-322.000000000000,-818.000000000000,
525.000000000000,904.000000000000,
-437.000000000000,-145.000000000000,
455.000000000000,250.000000000000,
355.000000000000,158.000000000000,
68.0000000000000,-527.000000000000,
1059.00000000000,1081.00000000000,
100.000000000000,619.000000000000,
509.000000000000,-36.0000000000000,
-164.000000000000,-577.000000000000,
-548.000000000000,-315.000000000000,
368.000000000000,-469.000000000000,
250.000000000000,-33.0000000000000,
428.000000000000,859.000000000000,
-1311.00000000000,367.000000000000,
-175.000000000000,-736.000000000000,
405.000000000000,-954.000000000000,
-486.000000000000,897.000000000000,
792.000000000000,-568.000000000000,
-34.0000000000000,-201.000000000000,
575.000000000000,824.000000000000,
-141.000000000000,-263.000000000000,
-509.000000000000,-258.000000000000,
872.000000000000,-184.000000000000,
587.000000000000,-533.000000000000,
1000.00000000000,-633.000000000000,
455.000000000000,61.0000000000000,
58.0000000000000,-144.000000000000,
490.000000000000,-430.000000000000,
27.0000000000000,-385.000000000000,
-87.0000000000000,98.0000000000000,
504.000000000000,538.000000000000,
-65.0000000000000,713.000000000000,
-383.000000000000,575.000000000000,
-933.000000000000,-379.000000000000,
-933.000000000000,-315.000000000000,
-54.0000000000000,270.000000000000,
414.000000000000,183.000000000000,
497.000000000000,811.000000000000,
-378.000000000000,288.000000000000,
-363.000000000000,-2.00000000000000,
-25.0000000000000,228.000000000000,
-1228.00000000000,-919.000000000000,
-607.000000000000,-251.000000000000,
274.000000000000,517.000000000000,
-22.0000000000000,-193.000000000000,
-145.000000000000,358.000000000000,
-237.000000000000,524.000000000000,
141.000000000000,-73.0000000000000,
-1118.00000000000,-42.0000000000000,
52.0000000000000,-1023.00000000000,
485.000000000000,195.000000000000,
-127.000000000000,301.000000000000,
865.000000000000,-442.000000000000,
-891.000000000000,121.000000000000,
521.000000000000,-371.000000000000,
1026.00000000000,414.000000000000,
741.000000000000,-342.000000000000,
501.000000000000,870.000000000000,
-603.000000000000,1475.00000000000,
-298.000000000000,397.000000000000,
-1270.00000000000,856.000000000000,
999.000000000000,295.000000000000,
645.000000000000,-122.000000000000,
-791.000000000000,15.0000000000000,
45.0000000000000,305.000000000000,
436.000000000000,-963.000000000000,
212.000000000000,-542.000000000000,
-1003.00000000000,454.000000000000,
-588.000000000000,318.000000000000,
-800.000000000000,620.000000000000,
-377.000000000000,220.000000000000,
545.000000000000,559.000000000000,
474.000000000000,-482.000000000000,
248.000000000000,111.000000000000,
-337.000000000000,983.000000000000,
333.000000000000,93.0000000000000,
-245.000000000000,213.000000000000,
-546.000000000000,-523.000000000000,
-56.0000000000000,-632.000000000000,
-928.000000000000,70.0000000000000,
-103.000000000000,47.0000000000000,
1034.00000000000,1072.00000000000,
-560.000000000000,157.000000000000,
-957.000000000000,-562.000000000000,
-69.0000000000000,804.000000000000,
224.000000000000,-273.000000000000,
125.000000000000,-99.0000000000000,
-743.000000000000,408.000000000000,
-260.000000000000,-665.000000000000,
-205.000000000000,-345.000000000000,
-979.000000000000,-69.0000000000000,
-309.000000000000,-1126.00000000000,
721.000000000000,-815.000000000000,
900.000000000000,1029.00000000000,
524.000000000000,727.000000000000,
202.000000000000,-290.000000000000,
720.000000000000,777.000000000000,
366.000000000000,31.0000000000000,
-927.000000000000,-238.000000000000,
-185.000000000000,575.000000000000,
-518.000000000000,-162.000000000000,
-995.000000000000,225.000000000000,
-166.000000000000,-589.000000000000,
52.0000000000000,-1134.00000000000,
205.000000000000,-286.000000000000,
71.0000000000000,-300.000000000000,
-931.000000000000,142.000000000000,
-189.000000000000,129.000000000000,
370.000000000000,-30.0000000000000,
467.000000000000,748.000000000000,
1094.00000000000,765.000000000000,
-677.000000000000,657.000000000000,
-775.000000000000,-785.000000000000,
-315.000000000000,-574.000000000000,
-3.00000000000000,895.000000000000,
-649.000000000000,-823.000000000000,
30.0000000000000,-749.000000000000,
900.000000000000,15.0000000000000,
-161.000000000000,1233.00000000000,
496.000000000000,276.000000000000,
-1203.00000000000,-990.000000000000,
-126.000000000000,-454.000000000000,
785.000000000000,-615.000000000000,
-323.000000000000,221.000000000000,
393.000000000000,399.000000000000,
-523.000000000000,820.000000000000,
-1044.00000000000,-436.000000000000,
-639.000000000000,-893.000000000000,
815.000000000000,224.000000000000,
-147.000000000000,464.000000000000,
-640.000000000000,419.000000000000,
-130.000000000000,-1453.00000000000,
-594.000000000000,399.000000000000,
-272.000000000000,180.000000000000,
-473.000000000000,-1057.00000000000,
403.000000000000,775.000000000000,
-840.000000000000,617.000000000000,
155.000000000000,649.000000000000,
604.000000000000,-233.000000000000,
-836.000000000000,722.000000000000,
541.000000000000,311.000000000000,
-863.000000000000,24.0000000000000,
-1108.00000000000,160.000000000000,
-491.000000000000,-1538.00000000000,
149.000000000000,-128.000000000000,
840.000000000000,-90.0000000000000,
372.000000000000,448.000000000000,
-139.000000000000,518.000000000000,
248.000000000000,-126.000000000000,
778.000000000000,744.000000000000,
-1063.00000000000,415.000000000000,
100.000000000000,-760.000000000000,
1019.00000000000,-14.0000000000000,
-80.0000000000000,1403.00000000000,
9.00000000000000,-63.0000000000000,
-1050.00000000000,-214.000000000000,
-433.000000000000,421.000000000000,
-542.000000000000,510.000000000000,
-1231.00000000000,662.000000000000,
-664.000000000000,-415.000000000000,
-655.000000000000,-554.000000000000,
-149.000000000000,-1250.00000000000,
520.000000000000,-871.000000000000,
372.000000000000,422.000000000000,
-547.000000000000,249.000000000000,
368.000000000000,3.00000000000000,
376.000000000000,492.000000000000,
460.000000000000,898.000000000000,
950.000000000000,86.0000000000000,
-507.000000000000,813.000000000000,
486.000000000000,518.000000000000,
-489.000000000000,-146.000000000000,
-1296.00000000000,557.000000000000,
-198.000000000000,316.000000000000,
-131.000000000000,107.000000000000,
-311.000000000000,298.000000000000,
-769.000000000000,1412.00000000000,
137.000000000000,170.000000000000,
-266.000000000000,-114.000000000000,
-471.000000000000,589.000000000000,
11.0000000000000,-860.000000000000,
-111.000000000000,593.000000000000,
172.000000000000,822.000000000000,
257.000000000000,-488.000000000000,
-34.0000000000000,618.000000000000,
-468.000000000000,676.000000000000,
833.000000000000,-225.000000000000,
427.000000000000,256.000000000000,
-22.0000000000000,76.0000000000000,
268.000000000000,-607.000000000000,
-1307.00000000000,-217.000000000000,
-535.000000000000,-373.000000000000,
-367.000000000000,318.000000000000,
-1043.00000000000,133.000000000000,
549.000000000000,-336.000000000000,
618.000000000000,701.000000000000,
-572.000000000000,1029.00000000000,
-86.0000000000000,562.000000000000,
-382.000000000000,19.0000000000000,
-1038.00000000000,-184.000000000000,
336.000000000000,-392.000000000000,
-430.000000000000,-129.000000000000,
-978.000000000000,-218.000000000000,
-349.000000000000,-291.000000000000,
-626.000000000000,205.000000000000,
1019.00000000000,-121.000000000000,
131.000000000000,567.000000000000,
-276.000000000000,847.000000000000,
695.000000000000,272.000000000000,
-202.000000000000,924.000000000000,
-737.000000000000,702.000000000000,
-559.000000000000,-286.000000000000,
54.0000000000000,-994.000000000000,
67.0000000000000,-108.000000000000,
-128.000000000000,-353.000000000000,
469.000000000000,-1297.00000000000,
301.000000000000,452.000000000000,
-576.000000000000,-338.000000000000,
-208.000000000000,-1299.00000000000,
-128.000000000000,151.000000000000,
536.000000000000,285.000000000000,
-200.000000000000,770.000000000000,
-872.000000000000,817.000000000000,
-337.000000000000,178.000000000000,
-766.000000000000,53.0000000000000,
467.000000000000,553.000000000000,
342.000000000000,517.000000000000,
-351.000000000000,378.000000000000,
699.000000000000,556.000000000000,
386.000000000000,-288.000000000000,
-30.0000000000000,-294.000000000000,
124.000000000000,50.0000000000000,
498.000000000000,-122.000000000000,
383.000000000000,-127.000000000000,
-929.000000000000,1081.00000000000,
393.000000000000,203.000000000000,
419.000000000000,-541.000000000000,
-388.000000000000,498.000000000000,
323.000000000000,-749.000000000000,
367.000000000000,-369.000000000000,
421.000000000000,-193.000000000000,
-167.000000000000,-407.000000000000,
-92.0000000000000,-476.000000000000,
-109.000000000000,-1083.00000000000,
812.000000000000,-496.000000000000,
580.000000000000,-237.000000000000,
223.000000000000,863.000000000000,
718.000000000000,432.000000000000,
187.000000000000,-828.000000000000,
927.000000000000,-132.000000000000,
831.000000000000,397.000000000000,
642.000000000000,-462.000000000000,
151.000000000000,-295.000000000000,
-682.000000000000,152.000000000000,
216.000000000000,-940.000000000000,
443.000000000000,-75.0000000000000,
-49.0000000000000,14.0000000000000,
-373.000000000000,-297.000000000000,
33.0000000000000,107.000000000000,
-355.000000000000,-705.000000000000,
-522.000000000000,600.000000000000,
281.000000000000,191.000000000000,
-121.000000000000,-877.000000000000,
-204.000000000000,332.000000000000,
769.000000000000,70.0000000000000,
152.000000000000,-84.0000000000000,
-486.000000000000,355.000000000000,
487.000000000000,220.000000000000,
305.000000000000,-626.000000000000,
801.000000000000,-4.00000000000000,
-36.0000000000000,813.000000000000,
-1472.00000000000,888.000000000000,
762.000000000000,297.000000000000,
-421.000000000000,-407.000000000000,
-573.000000000000,387.000000000000,
508.000000000000,-528.000000000000,
-790.000000000000,395.000000000000,
1068.00000000000,-29.0000000000000,
-762.000000000000,-385.000000000000,
-728.000000000000,346.000000000000,
-219.000000000000,-652.000000000000,
-994.000000000000,-399.000000000000,
-193.000000000000,-536.000000000000,
-654.000000000000,1083.00000000000,
602.000000000000,-3.00000000000000,
-540.000000000000,-251.000000000000,
377.000000000000,697.000000000000,
-21.0000000000000,-469.000000000000,
-85.0000000000000,-10.0000000000000,
630.000000000000,-477.000000000000,
-963.000000000000,987.000000000000,
-603.000000000000,-12.0000000000000,
-944.000000000000,-778.000000000000,
83.0000000000000,-644.000000000000,
81.0000000000000,-1309.00000000000,
26.0000000000000,707.000000000000,
-537.000000000000,-732.000000000000,
-166.000000000000,269.000000000000,
300.000000000000,206.000000000000,
-1434.00000000000,-116.000000000000,
627.000000000000,980.000000000000,
617.000000000000,-289.000000000000,
80.0000000000000,1146.00000000000,
-653.000000000000,110.000000000000,
-1337.00000000000,-700.000000000000,
89.0000000000000,-414.000000000000,
-278.000000000000,415.000000000000,
361.000000000000,-208.000000000000,
-22.0000000000000,-217.000000000000,
772.000000000000,994.000000000000,
-232.000000000000,-807.000000000000,
-1091.00000000000,556.000000000000,
438.000000000000,-420.000000000000,
-909.000000000000,-1414.00000000000,
131.000000000000,123.000000000000,
-398.000000000000,47.0000000000000,
-32.0000000000000,-463.000000000000,
1233.00000000000,138.000000000000,
-453.000000000000,877.000000000000,
-659.000000000000,-120.000000000000,
-460.000000000000,-480.000000000000,
425.000000000000,-331.000000000000,
-289.000000000000,-49.0000000000000,
-867.000000000000,-453.000000000000,
-396.000000000000,146.000000000000,
-67.0000000000000,1176.00000000000,
23.0000000000000,-539.000000000000,
-142.000000000000,-158.000000000000,
355.000000000000,-714.000000000000,
64.0000000000000,-970.000000000000,
497.000000000000,113.000000000000,
226.000000000000,-1318.00000000000,
330.000000000000,653.000000000000,
530.000000000000,706.000000000000,
120.000000000000,-465.000000000000,
-195.000000000000,1337.00000000000,
-334.000000000000,441.000000000000,
378.000000000000,-524.000000000000,
-254.000000000000,106.000000000000,
-751.000000000000,-284.000000000000,
-887.000000000000,-864.000000000000,
-989.000000000000,-43.0000000000000,
-40.0000000000000,289.000000000000,
364.000000000000,216.000000000000,
1143.00000000000,-111.000000000000,
855.000000000000,717.000000000000,
31.0000000000000,931.000000000000,
-614.000000000000,-505.000000000000,
-887.000000000000,-728.000000000000,
582.000000000000,-1078.00000000000,
-647.000000000000,-662.000000000000,
353.000000000000,-591.000000000000,
1129.00000000000,-252.000000000000,
19.0000000000000,1113.00000000000,
652.000000000000,593.000000000000,
-447.000000000000,905.000000000000,
-107.000000000000,-415.000000000000,
517.000000000000,-812.000000000000,
-156.000000000000,936.000000000000,
-626.000000000000,443.000000000000,
509.000000000000,330.000000000000,
516.000000000000,-70.0000000000000,
-486.000000000000,-273.000000000000,
79.0000000000000,-675.000000000000,
177.000000000000,-1235.00000000000,
15.0000000000000,-321.000000000000,
-311.000000000000,55.0000000000000,
488.000000000000,-362.000000000000,
644.000000000000,810.000000000000,
-377.000000000000,180.000000000000,
327.000000000000,-1103.00000000000,
467.000000000000,-823.000000000000,
86.0000000000000,-52.0000000000000,
643.000000000000,775.000000000000,
151.000000000000,-186.000000000000,
583.000000000000,587.000000000000,
672.000000000000,399.000000000000,
783.000000000000,116.000000000000,
670.000000000000,336.000000000000,
147.000000000000,-70.0000000000000,
620.000000000000,418.000000000000,
106.000000000000,-688.000000000000,
287.000000000000,337.000000000000,
744.000000000000,212.000000000000,
311.000000000000,-803.000000000000,
1022.00000000000,714.000000000000,
1025.00000000000,483.000000000000,
-663.000000000000,80.0000000000000,
-1106.00000000000,68.0000000000000,
-490.000000000000,-1148.00000000000,
395.000000000000,390.000000000000,
428.000000000000,771.000000000000,
-300.000000000000,-211.000000000000,
575.000000000000,868.000000000000,
-1073.00000000000,677.000000000000,
-209.000000000000,-134.000000000000,
541.000000000000,53.0000000000000,
-919.000000000000,1157.00000000000,
894.000000000000,-113.000000000000,
391.000000000000,403.000000000000,
-478.000000000000,243.000000000000,
-1.00000000000000,-985.000000000000,
331.000000000000,964.000000000000,
-449.000000000000,-97.0000000000000,
-158.000000000000,-894.000000000000,
621.000000000000,-666.000000000000,
337.000000000000,-375.000000000000,
863.000000000000,-325.000000000000,
1024.00000000000,443.000000000000,
478.000000000000,981.000000000000,
-814.000000000000,-779.000000000000,
-761.000000000000,495.000000000000,
-387.000000000000,1156.00000000000,
-65.0000000000000,-62.0000000000000,
276.000000000000,611.000000000000,
-1109.00000000000,645.000000000000,
422.000000000000,-615.000000000000,
520.000000000000,233.000000000000,
-860.000000000000,225.000000000000,
263.000000000000,-1862.00000000000,
703.000000000000,-11.0000000000000,
568.000000000000,399.000000000000,
-407.000000000000,-171.000000000000,
624.000000000000,493.000000000000,
58.0000000000000,432.000000000000,
-1066.00000000000,1290.00000000000,
-293.000000000000,-953.000000000000,
-129.000000000000,-737.000000000000,
864.000000000000,-499.000000000000,
301.000000000000,-862.000000000000,
1069.00000000000,567.000000000000,
182.000000000000,-558.000000000000,
253.000000000000,248.000000000000,
720.000000000000,456.000000000000,
-675.000000000000,329.000000000000,
268.000000000000,327.000000000000,
-998.000000000000,-215.000000000000,
-819.000000000000,-194.000000000000,
19.0000000000000,66.0000000000000,
430.000000000000,-525.000000000000,
959.000000000000,-1436.00000000000,
886.000000000000,943.000000000000,
171.000000000000,155.000000000000,
-1238.00000000000,-188.000000000000,
652.000000000000,82.0000000000000,
-71.0000000000000,-1301.00000000000,
-79.0000000000000,-640.000000000000,
1262.00000000000,-1020.00000000000,
-179.000000000000,905.000000000000,
-460.000000000000,1388.00000000000,
-588.000000000000,561.000000000000,
-190.000000000000,947.000000000000,
-668.000000000000,-413.000000000000,
207.000000000000,-288.000000000000,
868.000000000000,-568.000000000000,
-198.000000000000,548.000000000000,
-248.000000000000,636.000000000000,
-72.0000000000000,-342.000000000000,
76.0000000000000,72.0000000000000,
411.000000000000,277.000000000000,
786.000000000000,111.000000000000,
-409.000000000000,-401.000000000000,
-679.000000000000,1060.00000000000,
-873.000000000000,-107.000000000000,
-1070.00000000000,-1531.00000000000,
585.000000000000,-523.000000000000,
1255.00000000000,494.000000000000,
283.000000000000,1117.00000000000,
-463.000000000000,-569.000000000000,
481.000000000000,459.000000000000,
-748.000000000000,197.000000000000,
-1062.00000000000,-336.000000000000,
226.000000000000,95.0000000000000,
-368.000000000000,-216.000000000000,
394.000000000000,1169.00000000000,
311.000000000000,-269.000000000000,
85.0000000000000,494.000000000000,
601.000000000000,446.000000000000,
387.000000000000,-705.000000000000,
459.000000000000,0.00000000000000,
-562.000000000000,62.0000000000000,
-951.000000000000,-58.0000000000000,
-664.000000000000,-1034.00000000000,
771.000000000000,348.000000000000,
683.000000000000,1002.00000000000,
-895.000000000000,893.000000000000,
-323.000000000000,1029.00000000000,
-1122.00000000000,463.000000000000,
-1131.00000000000,-850.000000000000,
-543.000000000000,-1451.00000000000,
-441.000000000000,-236.000000000000,
61.0000000000000,-271.000000000000,
-314.000000000000,390.000000000000,
-709.000000000000,361.000000000000,
-947.000000000000,-874.000000000000,
-1052.00000000000,-590.000000000000,
676.000000000000,-220.000000000000,
397.000000000000,-94.0000000000000,
-815.000000000000,-798.000000000000,
473.000000000000,-616.000000000000,
-216.000000000000,691.000000000000,
302.000000000000,411.000000000000,
873.000000000000,652.000000000000,
418.000000000000,578.000000000000,
626.000000000000,105.000000000000,
6.00000000000000,-200.000000000000,
185.000000000000,-16.0000000000000,
-352.000000000000,498.000000000000,
-216.000000000000,439.000000000000,
-507.000000000000,1049.00000000000,
-957.000000000000,502.000000000000,
-453.000000000000,-605.000000000000,
-1027.00000000000,-535.000000000000,
-754.000000000000,5.00000000000000,
52.0000000000000,608.000000000000,
-393.000000000000,128.000000000000,
-850.000000000000,-549.000000000000,
353.000000000000,141.000000000000,
845.000000000000,299.000000000000,
-81.0000000000000,-352.000000000000,
69.0000000000000,765.000000000000,
342.000000000000,-466.000000000000,
-91.0000000000000,-759.000000000000,
-391.000000000000,769.000000000000,
-728.000000000000,-311.000000000000,
-232.000000000000,521.000000000000,
-1062.00000000000,-120.000000000000,
-834.000000000000,-100.000000000000,
998.000000000000,198.000000000000,
-168.000000000000,-377.000000000000,
-505.000000000000,336.000000000000,
-93.0000000000000,-612.000000000000,
-62.0000000000000,-745.000000000000,
-485.000000000000,260.000000000000,
-91.0000000000000,-359.000000000000,
871.000000000000,-139.000000000000,
-306.000000000000,1289.00000000000,
449.000000000000,409.000000000000,
224.000000000000,381.000000000000,
-45.0000000000000,-229.000000000000,
839.000000000000,-924.000000000000,
-141.000000000000,662.000000000000,
-101.000000000000,-534.000000000000,
196.000000000000,-8.00000000000000,
-130.000000000000,771.000000000000,
-935.000000000000,-179.000000000000,
13.0000000000000,690.000000000000,
-229.000000000000,171.000000000000,
-362.000000000000,285.000000000000,
1002.00000000000,-573.000000000000,
145.000000000000,-692.000000000000,
-142.000000000000,574.000000000000,
-506.000000000000,291.000000000000,
-296.000000000000,790.000000000000,
173.000000000000,389.000000000000,
340.000000000000,30.0000000000000,
451.000000000000,-443.000000000000,
501.000000000000,9.00000000000000,
431.000000000000,-467.000000000000,
-521.000000000000,-458.000000000000,
-106.000000000000,1086.00000000000,
-750.000000000000,-268.000000000000,
-1402.00000000000,-456.000000000000,
-73.0000000000000,-19.0000000000000,
209.000000000000,-281.000000000000,
-533.000000000000,-717.000000000000,
297.000000000000,65.0000000000000,
244.000000000000,791.000000000000,
-607.000000000000,-958.000000000000,
544.000000000000,-265.000000000000,
570.000000000000,780.000000000000,
473.000000000000,-41.0000000000000,
920.000000000000,-530.000000000000,
67.0000000000000,-550.000000000000,
1099.00000000000,-172.000000000000,
340.000000000000,544.000000000000,
41.0000000000000,1207.00000000000,
656.000000000000,-70.0000000000000,
-637.000000000000,-165.000000000000,
681.000000000000,-780.000000000000,
-67.0000000000000,-259.000000000000,
212.000000000000,-260.000000000000,
1382.00000000000,-811.000000000000,
268.000000000000,1529.00000000000,
-683.000000000000,-380.000000000000,
226.000000000000,-211.000000000000,
1403.00000000000,1417.00000000000,
132.000000000000,302.000000000000,
-156.000000000000,-102.000000000000,
854.000000000000,-313.000000000000,
409.000000000000,952.000000000000,
-696.000000000000,609.000000000000,
329.000000000000,751.000000000000,
-57.0000000000000,317.000000000000,
-1165.00000000000,-969.000000000000,
-164.000000000000,-421.000000000000,
-706.000000000000,-978.000000000000,
138.000000000000,-1094.00000000000,
81.0000000000000,111.000000000000,
-726.000000000000,-524.000000000000,
984.000000000000,-523.000000000000,
-527.000000000000,1033.00000000000,
-630.000000000000,337.000000000000,
-687.000000000000,212.000000000000,
-8.00000000000000,-301.000000000000,
799.000000000000,-199.000000000000,
-836.000000000000,368.000000000000,
774.000000000000,-1275.00000000000,
439.000000000000,115.000000000000,
-52.0000000000000,-12.0000000000000,
767.000000000000,-948.000000000000,
98.0000000000000,822.000000000000,
-551.000000000000,-537.000000000000,
-734.000000000000,-456.000000000000,
-320.000000000000,122.000000000000,
288.000000000000,467.000000000000,
-367.000000000000,939.000000000000,
0.00000000000000,-759.000000000000,
721.000000000000,292.000000000000,
-961.000000000000,-275.000000000000,
-641.000000000000,145.000000000000,
-547.000000000000,836.000000000000,
-119.000000000000,-170.000000000000,
534.000000000000,-512.000000000000,
-767.000000000000,45.0000000000000,
-356.000000000000,902.000000000000,
-207.000000000000,-491.000000000000,
395.000000000000,219.000000000000,
543.000000000000,-309.000000000000,
-310.000000000000,-1199.00000000000,
891.000000000000,-394.000000000000,
-512.000000000000,43.0000000000000,
-1025.00000000000,-290.000000000000,
131.000000000000,-894.000000000000,
87.0000000000000,-80.0000000000000,
471.000000000000,-780.000000000000,
553.000000000000,-253.000000000000,
994.000000000000,553.000000000000,
695.000000000000,619.000000000000,
728.000000000000,880.000000000000,
-965.000000000000,358.000000000000,
-683.000000000000,285.000000000000,
285.000000000000,-643.000000000000,
-1056.00000000000,559.000000000000,
627.000000000000,-501.000000000000,
-196.000000000000,-937.000000000000,
-73.0000000000000,803.000000000000,
23.0000000000000,-647.000000000000,
-360.000000000000,169.000000000000,
413.000000000000,-480.000000000000,
63.0000000000000,-756.000000000000,
1310.00000000000,159.000000000000,
30.0000000000000,273.000000000000,
-516.000000000000,-303.000000000000,
-93.0000000000000,-561.000000000000,
-497.000000000000,1082.00000000000,
-407.000000000000,-299.000000000000,
774.000000000000,587.000000000000,
823.000000000000,573.000000000000,
-1226.00000000000,-406.000000000000,
-512.000000000000,797.000000000000,
405.000000000000,-352.000000000000,
121.000000000000,-18.0000000000000,
-716.000000000000,226.000000000000,
269.000000000000,-644.000000000000,
1125.00000000000,-422.000000000000,
192.000000000000,575.000000000000,
515.000000000000,413.000000000000,
-356.000000000000,-63.0000000000000,
-206.000000000000,585.000000000000,
634.000000000000,432.000000000000,
-1054.00000000000,948.000000000000,
-956.000000000000,304.000000000000,
184.000000000000,582.000000000000,
-580.000000000000,891.000000000000,
-572.000000000000,-1341.00000000000,
547.000000000000,-1000.00000000000,
-328.000000000000,326.000000000000,
9.00000000000000,962.000000000000,
890.000000000000,578.000000000000,
483.000000000000,392.000000000000,
594.000000000000,272.000000000000,
-389.000000000000,-190.000000000000,
-843.000000000000,955.000000000000,
-586.000000000000,233.000000000000,
-320.000000000000,-948.000000000000,
149.000000000000,-249.000000000000,
-298.000000000000,5.00000000000000,
-438.000000000000,97.0000000000000,
-981.000000000000,514.000000000000,
-763.000000000000,-315.000000000000,
-51.0000000000000,306.000000000000,
130.000000000000,676.000000000000,
644.000000000000,202.000000000000,
197.000000000000,1046.00000000000,
-16.0000000000000,758.000000000000,
-980.000000000000,-345.000000000000,
-733.000000000000,-917.000000000000,
754.000000000000,-497.000000000000,
655.000000000000,345.000000000000,
25.0000000000000,47.0000000000000,
-997.000000000000,513.000000000000,
-697.000000000000,-705.000000000000,
-94.0000000000000,-1097.00000000000,
834.000000000000,591.000000000000,
-73.0000000000000,-463.000000000000,
-420.000000000000,-329.000000000000,
543.000000000000,-826.000000000000,
-180.000000000000,-640.000000000000,
-279.000000000000,-193.000000000000,
-412.000000000000,-1122.00000000000,
587.000000000000,471.000000000000,
-357.000000000000,958.000000000000,
-814.000000000000,-469.000000000000,
944.000000000000,-496.000000000000,
292.000000000000,940.000000000000,
170.000000000000,1118.00000000000,
-19.0000000000000,347.000000000000,
349.000000000000,177.000000000000,
-325.000000000000,572.000000000000,
-937.000000000000,-143.000000000000,
623.000000000000,-659.000000000000,
343.000000000000,474.000000000000,
218.000000000000,-512.000000000000,
27.0000000000000,-181.000000000000,
-272.000000000000,-4.00000000000000,
-1023.00000000000,-965.000000000000,
-325.000000000000,728.000000000000,
744.000000000000,-875.000000000000,
462.000000000000,-323.000000000000,
402.000000000000,728.000000000000,
397.000000000000,-456.000000000000,
-244.000000000000,959.000000000000,
-641.000000000000,-340.000000000000,
44.0000000000000,-484.000000000000,
-775.000000000000,474.000000000000,
-645.000000000000,511.000000000000,
-78.0000000000000,191.000000000000,
-445.000000000000,700.000000000000,
-550.000000000000,776.000000000000,
-13.0000000000000,-735.000000000000,
869.000000000000,738.000000000000,
217.000000000000,-40.0000000000000,
497.000000000000,-1075.00000000000,
452.000000000000,-189.000000000000,
-385.000000000000,621.000000000000,
-181.000000000000,-174.000000000000,
236.000000000000,-959.000000000000,
486.000000000000,1349.00000000000,
-689.000000000000,-164.000000000000,
-117.000000000000,288.000000000000,
508.000000000000,-151.000000000000,
-1117.00000000000,-365.000000000000,
-212.000000000000,505.000000000000,
134.000000000000,-1457.00000000000,
296.000000000000,863.000000000000,
266.000000000000,777.000000000000,
-45.0000000000000,220.000000000000,
-153.000000000000,541.000000000000,
-338.000000000000,474.000000000000,
233.000000000000,425.000000000000,
-941.000000000000,-253.000000000000,
-351.000000000000,184.000000000000,
-2.00000000000000,-768.000000000000,
13.0000000000000,230.000000000000,
464.000000000000,499.000000000000,
-1274.00000000000,67.0000000000000,
-370.000000000000,-494.000000000000,
-617.000000000000,-825.000000000000,
-529.000000000000,218.000000000000,
737.000000000000,-736.000000000000,
147.000000000000,-815.000000000000,
167.000000000000,204.000000000000,
-510.000000000000,-14.0000000000000,
-333.000000000000,-455.000000000000,
231.000000000000,116.000000000000,
-405.000000000000,-82.0000000000000,
-165.000000000000,-134.000000000000,
657.000000000000,159.000000000000,
-697.000000000000,-532.000000000000,
-1069.00000000000,-1009.00000000000,
655.000000000000,-829.000000000000,
64.0000000000000,-51.0000000000000,
-1046.00000000000,236.000000000000,
175.000000000000,415.000000000000,
353.000000000000,105.000000000000,
-37.0000000000000,-1284.00000000000,
773.000000000000,381.000000000000,
-332.000000000000,314.000000000000,
-650.000000000000,-1123.00000000000,
1656.00000000000,360.000000000000,
-216.000000000000,-280.000000000000,
-55.0000000000000,604.000000000000,
966.000000000000,-372.000000000000,
-916.000000000000,449.000000000000,
74.0000000000000,154.000000000000,
-902.000000000000,-821.000000000000,
-572.000000000000,1134.00000000000,
-628.000000000000,-660.000000000000,
-465.000000000000,372.000000000000,
152.000000000000,26.0000000000000,
-1134.00000000000,418.000000000000,
-164.000000000000,1143.00000000000,
79.0000000000000,250.000000000000,
853.000000000000,598.000000000000,
759.000000000000,-239.000000000000,
209.000000000000,661.000000000000,
-210.000000000000,530.000000000000,
-286.000000000000,89.0000000000000,
499.000000000000,110.000000000000,
104.000000000000,142.000000000000,
857.000000000000,309.000000000000,
243.000000000000,615.000000000000,
-190.000000000000,719.000000000000,
14.0000000000000,460.000000000000,
-638.000000000000,127.000000000000,
-123.000000000000,-1106.00000000000,
-772.000000000000,-978.000000000000,
-866.000000000000,-750.000000000000,
-426.000000000000,-141.000000000000,
-658.000000000000,1169.00000000000,
134.000000000000,465.000000000000,
-223.000000000000,279.000000000000,
-669.000000000000,-56.0000000000000,
650.000000000000,-1097.00000000000,
448.000000000000,204.000000000000,
-248.000000000000,742.000000000000,
-569.000000000000,-821.000000000000,
-332.000000000000,7.00000000000000,
688.000000000000,601.000000000000,
-273.000000000000,58.0000000000000,
-541.000000000000,171.000000000000,
-334.000000000000,-219.000000000000,
-542.000000000000,-27.0000000000000,
106.000000000000,730.000000000000,
-238.000000000000,420.000000000000,
-851.000000000000,-80.0000000000000,
-470.000000000000,-401.000000000000,
-515.000000000000,909.000000000000,
-827.000000000000,434.000000000000,
-933.000000000000,-1273.00000000000,
-64.0000000000000,783.000000000000,
182.000000000000,415.000000000000,
-487.000000000000,-345.000000000000,
-192.000000000000,41.0000000000000,
644.000000000000,-340.000000000000,
666.000000000000,-939.000000000000,
37.0000000000000,-497.000000000000,
962.000000000000,168.000000000000,
653.000000000000,-1084.00000000000,
56.0000000000000,710.000000000000,
-501.000000000000,160.000000000000,
-1049.00000000000,-432.000000000000,
-278.000000000000,486.000000000000,
-1366.00000000000,-1217.00000000000,
-197.000000000000,-572.000000000000,
530.000000000000,668.000000000000,
-287.000000000000,464.000000000000,
580.000000000000,131.000000000000,
-119.000000000000,104.000000000000,
-321.000000000000,-179.000000000000,
-383.000000000000,430.000000000000,
540.000000000000,-48.0000000000000,
908.000000000000,-719.000000000000,
694.000000000000,146.000000000000,
446.000000000000,-444.000000000000,
-1185.00000000000,-525.000000000000,
-432.000000000000,170.000000000000,
-1115.00000000000,482.000000000000,
-123.000000000000,393.000000000000,
1170.00000000000,601.000000000000,
316.000000000000,60.0000000000000,
502.000000000000,33.0000000000000,
275.000000000000,1201.00000000000,
928.000000000000,218.000000000000,
-678.000000000000,-470.000000000000,
-887.000000000000,-87.0000000000000,
614.000000000000,-449.000000000000,
80.0000000000000,-346.000000000000,
380.000000000000,615.000000000000,
798.000000000000,614.000000000000,
-89.0000000000000,-92.0000000000000,
-174.000000000000,597.000000000000,
-426.000000000000,-48.0000000000000,
-284.000000000000,-728.000000000000,
201.000000000000,229.000000000000,
-1114.00000000000,-928.000000000000,
-390.000000000000,147.000000000000,
857.000000000000,-39.0000000000000,
594.000000000000,-701.000000000000,
-114.000000000000,1322.00000000000,
-17.0000000000000,-196.000000000000,
308.000000000000,636.000000000000,
-803.000000000000,571.000000000000,
-821.000000000000,-604.000000000000,
-681.000000000000,-39.0000000000000,
66.0000000000000,-468.000000000000,
274.000000000000,160.000000000000,
26.0000000000000,231.000000000000,
1178.00000000000,-247.000000000000,
338.000000000000,-60.0000000000000,
-150.000000000000,157.000000000000,
722.000000000000,-267.000000000000,
-219.000000000000,85.0000000000000,
-494.000000000000,84.0000000000000,
-181.000000000000,-337.000000000000,
255.000000000000,-21.0000000000000,
888.000000000000,314.000000000000,
-324.000000000000,606.000000000000,
-571.000000000000,-503.000000000000,
735.000000000000,-478.000000000000,
646.000000000000,1085.00000000000,
-1058.00000000000,762.000000000000,
-246.000000000000,254.000000000000,
-528.000000000000,438.000000000000,
-1022.00000000000,-848.000000000000,
1131.00000000000,-117.000000000000,
-627.000000000000,397.000000000000,
-579.000000000000,-274.000000000000,
-357.000000000000,691.000000000000,
-457.000000000000,-117.000000000000,
-185.000000000000,530.000000000000,
-735.000000000000,-49.0000000000000,
937.000000000000,-673.000000000000,
-229.000000000000,1824.00000000000,
-39.0000000000000,-6.00000000000000,
576.000000000000,-859.000000000000,
275.000000000000,482.000000000000,
244.000000000000,-487.000000000000,
335.000000000000,737.000000000000,
353.000000000000,-209.000000000000,
-345.000000000000,-311.000000000000,
520.000000000000,941.000000000000,
-262.000000000000,401.000000000000,
128.000000000000,1114.00000000000,
208.000000000000,86.0000000000000,
-266.000000000000,927.000000000000,
143.000000000000,10.0000000000000,
128.000000000000,-852.000000000000,
1217.00000000000,-488.000000000000,
348.000000000000,-845.000000000000,
429.000000000000,-171.000000000000,
939.000000000000,-556.000000000000,
135.000000000000,1188.00000000000,
-564.000000000000,529.000000000000,
-276.000000000000,-660.000000000000,
243.000000000000,723.000000000000,
-1074.00000000000,452.000000000000,
33.0000000000000,-686.000000000000,
-435.000000000000,106.000000000000,
-617.000000000000,-89.0000000000000,
902.000000000000,-1501.00000000000,
-103.000000000000,-65.0000000000000,
-70.0000000000000,-594.000000000000,
-182.000000000000,-527.000000000000,
-640.000000000000,690.000000000000,
-770.000000000000,-1023.00000000000,
-472.000000000000,-193.000000000000,
838.000000000000,27.0000000000000,
690.000000000000,1107.00000000000,
-616.000000000000,95.0000000000000,
726.000000000000,-845.000000000000,
48.0000000000000,798.000000000000,
-561.000000000000,-1216.00000000000,
1120.00000000000,166.000000000000,
-761.000000000000,-584.000000000000,
-587.000000000000,-416.000000000000,
-2.00000000000000,-400.000000000000,
-210.000000000000,-893.000000000000,
621.000000000000,544.000000000000,
178.000000000000,-1196.00000000000,
263.000000000000,176.000000000000,
-393.000000000000,-350.000000000000,
170.000000000000,-659.000000000000,
607.000000000000,769.000000000000,
-710.000000000000,885.000000000000,
104.000000000000,886.000000000000,
-8.00000000000000,41.0000000000000,
27.0000000000000,-318.000000000000,
492.000000000000,-103.000000000000,
-95.0000000000000,-74.0000000000000,
267.000000000000,-1516.00000000000,
-157.000000000000,-339.000000000000,
-388.000000000000,243.000000000000,
-122.000000000000,-1075.00000000000,
-103.000000000000,-230.000000000000,
666.000000000000,-115.000000000000,
741.000000000000,561.000000000000,
-738.000000000000,345.000000000000,
-1110.00000000000,-904.000000000000,
110.000000000000,-463.000000000000,
137.000000000000,-180.000000000000,
925.000000000000,-6.00000000000000,
1004.00000000000,212.000000000000,
580.000000000000,93.0000000000000,
955.000000000000,386.000000000000,
-419.000000000000,757.000000000000,
-634.000000000000,-209.000000000000,
-278.000000000000,-767.000000000000,
907.000000000000,-347.000000000000,
126.000000000000,471.000000000000,
-783.000000000000,-159.000000000000,
1236.00000000000,-1446.00000000000,
642.000000000000,-155.000000000000,
662.000000000000,142.000000000000,
-142.000000000000,-656.000000000000,
-485.000000000000,-502.000000000000,
195.000000000000,578.000000000000,
263.000000000000,1219.00000000000,
643.000000000000,-162.000000000000,
-276.000000000000,159.000000000000,
650.000000000000,-194.000000000000,
390.000000000000,-333.000000000000,
-89.0000000000000,592.000000000000,
-983.000000000000,-818.000000000000,
-651.000000000000,203.000000000000,
339.000000000000,139.000000000000,
-390.000000000000,-1217.00000000000,
1056.00000000000,59.0000000000000,
31.0000000000000,371.000000000000,
136.000000000000,-666.000000000000,
-133.000000000000,-77.0000000000000,
-796.000000000000,-75.0000000000000,
236.000000000000,-554.000000000000,
-590.000000000000,1245.00000000000,
422.000000000000,498.000000000000,
565.000000000000,67.0000000000000,
1015.00000000000,474.000000000000,
496.000000000000,-14.0000000000000,
-658.000000000000,1076.00000000000,
-679.000000000000,-665.000000000000,
-1177.00000000000,-871.000000000000,
-497.000000000000,-892.000000000000,
566.000000000000,-594.000000000000,
996.000000000000,1053.00000000000,
127.000000000000,236.000000000000,
998.000000000000,1370.00000000000,
486.000000000000,-686.000000000000,
-334.000000000000,393.000000000000,
1108.00000000000,342.000000000000,
471.000000000000,-949.000000000000,
-82.0000000000000,621.000000000000,
-649.000000000000,-823.000000000000,
53.0000000000000,1029.00000000000,
107.000000000000,-424.000000000000,
-284.000000000000,-993.000000000000,
-248.000000000000,604.000000000000,
87.0000000000000,352.000000000000,
1492.00000000000,1148.00000000000,
-1105.00000000000,776.000000000000,
-317.000000000000,-292.000000000000,
738.000000000000,225.000000000000,
-1103.00000000000,793.000000000000,
1149.00000000000,-323.000000000000,
-69.0000000000000,357.000000000000,
-942.000000000000,-389.000000000000,
-529.000000000000,-977.000000000000,
-168.000000000000,-356.000000000000,
-32.0000000000000,-1312.00000000000,
-552.000000000000,-207.000000000000,
1309.00000000000,487.000000000000,
637.000000000000,226.000000000000,
162.000000000000,312.000000000000,
-163.000000000000,167.000000000000,
92.0000000000000,227.000000000000,
181.000000000000,362.000000000000,
427.000000000000,309.000000000000,
554.000000000000,-1153.00000000000,
-884.000000000000,197.000000000000,
931.000000000000,282.000000000000,
352.000000000000,-482.000000000000,
180.000000000000,844.000000000000,
-271.000000000000,-4.00000000000000,
-1299.00000000000,279.000000000000,
446.000000000000,58.0000000000000,
218.000000000000,-1163.00000000000,
1050.00000000000,-76.0000000000000,
-34.0000000000000,902.000000000000,
-983.000000000000,-417.000000000000,
-100.000000000000,-1123.00000000000,
-532.000000000000,-266.000000000000,
-524.000000000000,-83.0000000000000,
-746.000000000000,574.000000000000,
-650.000000000000,-706.000000000000,
-603.000000000000,-909.000000000000,
-267.000000000000,450.000000000000,
-528.000000000000,-665.000000000000,
-144.000000000000,407.000000000000,
696.000000000000,650.000000000000,
571.000000000000,58.0000000000000,
-4.00000000000000,377.000000000000,
-1266.00000000000,670.000000000000,
124.000000000000,619.000000000000,
-5.00000000000000,-840.000000000000,
152.000000000000,-237.000000000000,
288.000000000000,13.0000000000000,
-971.000000000000,-102.000000000000,
972.000000000000,-407.000000000000,
339.000000000000,271.000000000000,
-472.000000000000,948.000000000000,
507.000000000000,-507.000000000000,
481.000000000000,-256.000000000000,
261.000000000000,-616.000000000000,
-4.00000000000000,-667.000000000000,
636.000000000000,-718.000000000000,
309.000000000000,418.000000000000,
-768.000000000000,865.000000000000,
-240.000000000000,-897.000000000000,
413.000000000000,1030.00000000000,
-509.000000000000,-26.0000000000000,
24.0000000000000,-680.000000000000,
-147.000000000000,-314.000000000000,
-235.000000000000,-1341.00000000000,
1220.00000000000,216.000000000000,
724.000000000000,224.000000000000,
-236.000000000000,-276.000000000000,
-360.000000000000,-856.000000000000,
-28.0000000000000,708.000000000000,
-415.000000000000,764.000000000000,
-845.000000000000,502.000000000000,
0.00000000000000,620.000000000000,
-242.000000000000,-1002.00000000000,
761.000000000000,7.00000000000000,
535.000000000000,-177.000000000000,
-624.000000000000,214.000000000000,
-316.000000000000,-579.000000000000,
-1020.00000000000,-1133.00000000000,
-265.000000000000,-787.000000000000,
-264.000000000000,-706.000000000000,
331.000000000000,1165.00000000000,
514.000000000000,-814.000000000000,
-877.000000000000,23.0000000000000,
99.0000000000000,133.000000000000,
544.000000000000,-495.000000000000,
858.000000000000,1583.00000000000,
494.000000000000,598.000000000000,
374.000000000000,62.0000000000000,
555.000000000000,-221.000000000000,
643.000000000000,-544.000000000000,
-430.000000000000,231.000000000000,
-1424.00000000000,13.0000000000000,
1000.00000000000,-1078.00000000000,
-294.000000000000,354.000000000000,
-1028.00000000000,1019.00000000000,
-287.000000000000,-151.000000000000,
-376.000000000000,-655.000000000000,
1020.00000000000,-429.000000000000,
159.000000000000,896.000000000000,
474.000000000000,648.000000000000,
-743.000000000000,-26.0000000000000,
-562.000000000000,43.0000000000000,
1241.00000000000,428.000000000000,
137.000000000000,744.000000000000,
185.000000000000,753.000000000000,
395.000000000000,70.0000000000000,
944.000000000000,-532.000000000000,
-141.000000000000,1292.00000000000,
-151.000000000000,833.000000000000,
-205.000000000000,-1116.00000000000,
-972.000000000000,578.000000000000,
-577.000000000000,821.000000000000,
-1014.00000000000,-91.0000000000000,
159.000000000000,118.000000000000,
707.000000000000,102.000000000000,
-290.000000000000,-679.000000000000,
216.000000000000,-1194.00000000000,
1039.00000000000,514.000000000000,
-235.000000000000,2.00000000000000,
-512.000000000000,-703.000000000000,
-125.000000000000,524.000000000000,
-695.000000000000,447.000000000000,
330.000000000000,48.0000000000000,
-299.000000000000,345.000000000000,
-474.000000000000,180.000000000000,
579.000000000000,-884.000000000000,
-406.000000000000,341.000000000000,
-307.000000000000,-484.000000000000,
-164.000000000000,-1039.00000000000,
-83.0000000000000,872.000000000000,
34.0000000000000,77.0000000000000,
1090.00000000000,656.000000000000,
468.000000000000,-627.000000000000,
-722.000000000000,539.000000000000,
761.000000000000,463.000000000000,
4.00000000000000,47.0000000000000,
-529.000000000000,1231.00000000000,
-786.000000000000,-941.000000000000,
16.0000000000000,647.000000000000,
185.000000000000,-658.000000000000,
281.000000000000,224.000000000000,
842.000000000000,716.000000000000,
-1181.00000000000,-990.000000000000,
410.000000000000,-143.000000000000,
-326.000000000000,-1041.00000000000,
-469.000000000000,360.000000000000,
-34.0000000000000,496.000000000000,
-1336.00000000000,-271.000000000000,
1128.00000000000,-21.0000000000000,
-156.000000000000,51.0000000000000,
-40.0000000000000,-868.000000000000,
-43.0000000000000,-834.000000000000,
-37.0000000000000,55.0000000000000,
36.0000000000000,-258.000000000000,
-1107.00000000000,-591.000000000000,
1079.00000000000,-465.000000000000,
-542.000000000000,1091.00000000000,
-626.000000000000,765.000000000000,
692.000000000000,106.000000000000,
-567.000000000000,411.000000000000,
-325.000000000000,361.000000000000,
7.00000000000000,-690.000000000000,
-491.000000000000,-422.000000000000,
149.000000000000,1185.00000000000,
-258.000000000000,365.000000000000,
-989.000000000000,-838.000000000000,
-175.000000000000,-700.000000000000,
681.000000000000,-243.000000000000,
571.000000000000,438.000000000000,
-290.000000000000,-291.000000000000,
512.000000000000,-1257.00000000000,
798.000000000000,175.000000000000,
-353.000000000000,965.000000000000,
405.000000000000,125.000000000000,
-201.000000000000,-147.000000000000,
-690.000000000000,-425.000000000000,
-5.00000000000000,-623.000000000000,
-1032.00000000000,269.000000000000,
148.000000000000,-851.000000000000,
-328.000000000000,-526.000000000000,
-715.000000000000,1145.00000000000,
379.000000000000,-984.000000000000,
-288.000000000000,-475.000000000000,
-47.0000000000000,480.000000000000,
-350.000000000000,795.000000000000,
-1007.00000000000,422.000000000000,
237.000000000000,247.000000000000,
-341.000000000000,906.000000000000,
-787.000000000000,-1300.00000000000,
839.000000000000,427.000000000000,
-838.000000000000,720.000000000000,
-656.000000000000,-1091.00000000000,
1125.00000000000,-666.000000000000,
-545.000000000000,-86.0000000000000,
-300.000000000000,738.000000000000,
-427.000000000000,-747.000000000000,
-1073.00000000000,-604.000000000000,
19.0000000000000,-702.000000000000,
-262.000000000000,-766.000000000000,
-75.0000000000000,-891.000000000000,
463.000000000000,-294.000000000000,
1145.00000000000,877.000000000000,
-667.000000000000,656.000000000000,
-374.000000000000,951.000000000000,
594.000000000000,-1327.00000000000,
-912.000000000000,450.000000000000,
843.000000000000,-96.0000000000000,
628.000000000000,-746.000000000000,
1098.00000000000,1521.00000000000,
425.000000000000,-985.000000000000,
162.000000000000,-357.000000000000,
89.0000000000000,-475.000000000000,
-1027.00000000000,-348.000000000000,
461.000000000000,971.000000000000,
-1331.00000000000,207.000000000000,
-222.000000000000,-531.000000000000,
1308.00000000000,-992.000000000000,
-114.000000000000,-201.000000000000,
-157.000000000000,508.000000000000,
247.000000000000,564.000000000000,
399.000000000000,951.000000000000,
-1045.00000000000,474.000000000000,
143.000000000000,-673.000000000000,
-379.000000000000,663.000000000000,
-560.000000000000,65.0000000000000,
528.000000000000,101.000000000000,
147.000000000000,1194.00000000000,
615.000000000000,91.0000000000000,
-705.000000000000,627.000000000000,
-164.000000000000,799.000000000000,
-612.000000000000,-97.0000000000000,
-531.000000000000,-783.000000000000,
1414.00000000000,-71.0000000000000,
65.0000000000000,711.000000000000,
-646.000000000000,261.000000000000,
218.000000000000,-418.000000000000,
489.000000000000,131.000000000000,
-350.000000000000,594.000000000000,
-652.000000000000,-461.000000000000,
-472.000000000000,-724.000000000000,
-689.000000000000,-722.000000000000,
-556.000000000000,-824.000000000000,
-379.000000000000,-622.000000000000,
-13.0000000000000,-787.000000000000,
538.000000000000,483.000000000000,
99.0000000000000,948.000000000000,
-420.000000000000,-674.000000000000,
733.000000000000,245.000000000000,
605.000000000000,-23.0000000000000,
-134.000000000000,-1276.00000000000,
121.000000000000,-342.000000000000,
-440.000000000000,-549.000000000000,
817.000000000000,-742.000000000000,
236.000000000000,-482.000000000000,
-871.000000000000,-714.000000000000,
143.000000000000,-541.000000000000,
-677.000000000000,-83.0000000000000,
222.000000000000,527.000000000000,
-112.000000000000,421.000000000000,
-814.000000000000,-665.000000000000,
215.000000000000,168.000000000000,
8.00000000000000,446.000000000000,
448.000000000000,-1136.00000000000,
1054.00000000000,-526.000000000000,
984.000000000000,-795.000000000000,
-345.000000000000,-170.000000000000,
-488.000000000000,842.000000000000,
-277.000000000000,-1137.00000000000,
-243.000000000000,369.000000000000,
-166.000000000000,284.000000000000,
-832.000000000000,-87.0000000000000,
-627.000000000000,-310.000000000000,
316.000000000000,-1189.00000000000,
1200.00000000000,855.000000000000,
351.000000000000,418.000000000000,
873.000000000000,229.000000000000,
991.000000000000,-428.000000000000,
-84.0000000000000,0.00000000000000,
990.000000000000,421.000000000000,
754.000000000000,-808.000000000000,
605.000000000000,-157.000000000000,
698.000000000000,568.000000000000,
-598.000000000000,634.000000000000,
-554.000000000000,430.000000000000,
339.000000000000,1202.00000000000,
-596.000000000000,-267.000000000000,
-1496.00000000000,-688.000000000000,
591.000000000000,217.000000000000,
-555.000000000000,-953.000000000000,
-73.0000000000000,440.000000000000,
292.000000000000,643.000000000000,
-1302.00000000000,355.000000000000,
1103.00000000000,312.000000000000,
-750.000000000000,200.000000000000,
-637.000000000000,321.000000000000,
428.000000000000,-237.000000000000,
-301.000000000000,-632.000000000000,
450.000000000000,-1127.00000000000,
-305.000000000000,62.0000000000000,
-65.0000000000000,120.000000000000,
25.0000000000000,553.000000000000,
64.0000000000000,1212.00000000000,
-638.000000000000,435.000000000000,
-766.000000000000,542.000000000000,
-1074.00000000000,90.0000000000000,
-1035.00000000000,-441.000000000000,
394.000000000000,-1089.00000000000,
-65.0000000000000,589.000000000000,
-229.000000000000,523.000000000000,
-584.000000000000,-901.000000000000,
-292.000000000000,737.000000000000,
-595.000000000000,-784.000000000000,
-264.000000000000,-359.000000000000,
1050.00000000000,1151.00000000000,
-914.000000000000,-547.000000000000,
-947.000000000000,-385.000000000000,
344.000000000000,344.000000000000,
418.000000000000,-732.000000000000,
175.000000000000,-955.000000000000,
-209.000000000000,348.000000000000,
-358.000000000000,-214.000000000000,
-346.000000000000,109.000000000000,
-394.000000000000,-249.000000000000,
-1298.00000000000,-939.000000000000,
102.000000000000,507.000000000000,
440.000000000000,273.000000000000,
-883.000000000000,835.000000000000,
-729.000000000000,13.0000000000000,
-989.000000000000,-912.000000000000,
-623.000000000000,-806.000000000000,
182.000000000000,-1445.00000000000,
1204.00000000000,-508.000000000000,
-238.000000000000,717.000000000000,
-1019.00000000000,1231.00000000000,
-709.000000000000,116.000000000000,
-1059.00000000000,706.000000000000,
643.000000000000,-71.0000000000000,
18.0000000000000,-1215.00000000000,
383.000000000000,-2.00000000000000,
1048.00000000000,-691.000000000000,
-119.000000000000,841.000000000000,
124.000000000000,1023.00000000000,
-268.000000000000,-871.000000000000,
677.000000000000,93.0000000000000,
784.000000000000,695.000000000000,
-182.000000000000,-611.000000000000,
-1213.00000000000,-317.000000000000,
49.0000000000000,478.000000000000,
699.000000000000,115.000000000000,
-297.000000000000,-122.000000000000,
1024.00000000000,-455.000000000000,
-315.000000000000,484.000000000000,
-805.000000000000,449.000000000000,
-556.000000000000,-747.000000000000,
-872.000000000000,-646.000000000000,
425.000000000000,-106.000000000000,
-106.000000000000,345.000000000000,
-296.000000000000,-904.000000000000,
783.000000000000,-600.000000000000,
726.000000000000,500.000000000000,
276.000000000000,-641.000000000000,
627.000000000000,20.0000000000000,
290.000000000000,411.000000000000,
-524.000000000000,-103.000000000000,
-593.000000000000,-103.000000000000,
476.000000000000,-375.000000000000,
863.000000000000,11.0000000000000,
-952.000000000000,-195.000000000000,
-10.0000000000000,-635.000000000000,
1128.00000000000,-39.0000000000000,
-338.000000000000,730.000000000000,
-268.000000000000,-486.000000000000,
-48.0000000000000,-172.000000000000,
143.000000000000,531.000000000000,
-154.000000000000,-322.000000000000,
-148.000000000000,-5.00000000000000,
203.000000000000,-192.000000000000,
-586.000000000000,662.000000000000,
-796.000000000000,486.000000000000,
-657.000000000000,-1092.00000000000,
-4.00000000000000,-484.000000000000,
382.000000000000,671.000000000000,
380.000000000000,924.000000000000,
-267.000000000000,159.000000000000,
-530.000000000000,-121.000000000000,
278.000000000000,448.000000000000,
260.000000000000,-13.0000000000000,
-128.000000000000,-377.000000000000,
524.000000000000,132.000000000000,
514.000000000000,-614.000000000000,
-1113.00000000000,-698.000000000000,
-417.000000000000,-237.000000000000,
335.000000000000,-594.000000000000,
-974.000000000000,313.000000000000,
305.000000000000,855.000000000000,
-328.000000000000,371.000000000000,
-1428.00000000000,883.000000000000,
688.000000000000,483.000000000000,
-39.0000000000000,-321.000000000000,
-515.000000000000,-746.000000000000,
1163.00000000000,-345.000000000000,
514.000000000000,410.000000000000,
-27.0000000000000,518.000000000000,
381.000000000000,1220.00000000000,
-346.000000000000,784.000000000000,
435.000000000000,-296.000000000000,
700.000000000000,-244.000000000000,
-71.0000000000000,-505.000000000000,
734.000000000000,-455.000000000000,
-936.000000000000,1166.00000000000,
-379.000000000000,813.000000000000,
323.000000000000,-361.000000000000,
305.000000000000,-212.000000000000,
1115.00000000000,-879.000000000000,
-887.000000000000,-23.0000000000000,
733.000000000000,29.0000000000000,
1050.00000000000,-1039.00000000000,
8.00000000000000,-164.000000000000,
359.000000000000,647.000000000000,
743.000000000000,1332.00000000000,
494.000000000000,459.000000000000,
-477.000000000000,858.000000000000,
663.000000000000,635.000000000000,
-996.000000000000,-223.000000000000,
-352.000000000000,-633.000000000000,
1361.00000000000,-1238.00000000000,
-89.0000000000000,1097.00000000000,
-684.000000000000,-197.000000000000,
485.000000000000,-352.000000000000,
778.000000000000,917.000000000000,
-1349.00000000000,-354.000000000000,
279.000000000000,-322.000000000000,
1029.00000000000,-115.000000000000,
-81.0000000000000,799.000000000000,
211.000000000000,-685.000000000000,
45.0000000000000,-482.000000000000,
-322.000000000000,-103.000000000000,
-959.000000000000,-134.000000000000,
833.000000000000,-14.0000000000000,
-360.000000000000,-821.000000000000,
-389.000000000000,411.000000000000,
792.000000000000,-15.0000000000000,
-1231.00000000000,174.000000000000,
-331.000000000000,166.000000000000,
-583.000000000000,41.0000000000000,
-1136.00000000000,-37.0000000000000,
71.0000000000000,-1161.00000000000,
87.0000000000000,-262.000000000000,
-42.0000000000000,-1072.00000000000,
863.000000000000,-366.000000000000,
55.0000000000000,772.000000000000,
-1228.00000000000,-406.000000000000,
290.000000000000,-909.000000000000,
157.000000000000,189.000000000000,
-335.000000000000,787.000000000000,
92.0000000000000,-874.000000000000,
505.000000000000,483.000000000000,
323.000000000000,569.000000000000,
-903.000000000000,-366.000000000000,
450.000000000000,326.000000000000,
-640.000000000000,-205.000000000000,
-702.000000000000,141.000000000000,
726.000000000000,-245.000000000000,
552.000000000000,-553.000000000000,
480.000000000000,521.000000000000,
-1149.00000000000,282.000000000000,
426.000000000000,-1479.00000000000,
614.000000000000,-778.000000000000,
392.000000000000,763.000000000000,
387.000000000000,496.000000000000,
-647.000000000000,-500.000000000000,
716.000000000000,63.0000000000000,
457.000000000000,1139.00000000000,
812.000000000000,868.000000000000,
-503.000000000000,831.000000000000,
-540.000000000000,-317.000000000000,
554.000000000000,-1330.00000000000,
144.000000000000,-3.00000000000000,
356.000000000000,425.000000000000,
156.000000000000,1039.00000000000,
403.000000000000,1025.00000000000,
-1005.00000000000,575.000000000000,
-479.000000000000,582.000000000000,
621.000000000000,-682.000000000000,
339.000000000000,-28.0000000000000,
307.000000000000,76.0000000000000,
-410.000000000000,-622.000000000000,
576.000000000000,-125.000000000000,
146.000000000000,1083.00000000000,
-1133.00000000000,1021.00000000000,
-561.000000000000,-1209.00000000000,
782.000000000000,-458.000000000000,
410.000000000000,60.0000000000000,
-120.000000000000,-121.000000000000,
1119.00000000000,85.0000000000000,
439.000000000000,236.000000000000,
350.000000000000,1478.00000000000,
-221.000000000000,372.000000000000,
-376.000000000000,-675.000000000000,
389.000000000000,-64.0000000000000,
-1133.00000000000,48.0000000000000,
-270.000000000000,-1578.00000000000,
372.000000000000,-793.000000000000,
-244.000000000000,-294.000000000000,
-651.000000000000,-976.000000000000,
347.000000000000,942.000000000000,
877.000000000000,-695.000000000000,
744.000000000000,605.000000000000,
451.000000000000,1031.00000000000,
-1186.00000000000,-1130.00000000000,
856.000000000000,618.000000000000,
222.000000000000,282.000000000000,
-1153.00000000000,-228.000000000000,
-218.000000000000,-1115.00000000000,
-822.000000000000,238.000000000000,
-73.0000000000000,542.000000000000,
-908.000000000000,-1532.00000000000,
-280.000000000000,-431.000000000000,
182.000000000000,420.000000000000,
374.000000000000,-300.000000000000,
465.000000000000,-208.000000000000,
-560.000000000000,528.000000000000,
-260.000000000000,-473.000000000000,
-1060.00000000000,-442.000000000000,
526.000000000000,211.000000000000,
-133.000000000000,162.000000000000,
-1144.00000000000,-128.000000000000,
544.000000000000,-885.000000000000,
586.000000000000,-305.000000000000,
441.000000000000,690.000000000000,
-265.000000000000,680.000000000000,
-626.000000000000,706.000000000000,
-1047.00000000000,472.000000000000,
69.0000000000000,-916.000000000000,
796.000000000000,275.000000000000,
310.000000000000,1060.00000000000,
430.000000000000,54.0000000000000,
-415.000000000000,171.000000000000,
929.000000000000,-136.000000000000,
563.000000000000,43.0000000000000,
339.000000000000,6.00000000000000,
152.000000000000,-745.000000000000,
-304.000000000000,-201.000000000000,
1010.00000000000,-1055.00000000000,
-388.000000000000,132.000000000000,
-375.000000000000,898.000000000000,
-792.000000000000,-975.000000000000,
-753.000000000000,139.000000000000,
307.000000000000,248.000000000000,
-304.000000000000,669.000000000000,
268.000000000000,691.000000000000,
493.000000000000,963.000000000000,
655.000000000000,418.000000000000,
-84.0000000000000,-471.000000000000,
-605.000000000000,534.000000000000,
-463.000000000000,-744.000000000000,
248.000000000000,299.000000000000,
-288.000000000000,-97.0000000000000,
-125.000000000000,-949.000000000000,
1441.00000000000,-625.000000000000,
246.000000000000,-710.000000000000,
842.000000000000,-171.000000000000,
294.000000000000,-944.000000000000,
-538.000000000000,166.000000000000,
855.000000000000,-340.000000000000,
-313.000000000000,-287.000000000000,
-473.000000000000,891.000000000000,
-21.0000000000000,-276.000000000000,
79.0000000000000,-275.000000000000,
320.000000000000,579.000000000000,
-308.000000000000,831.000000000000,
-320.000000000000,203.000000000000,
24.0000000000000,18.0000000000000,
-374.000000000000,-338.000000000000,
-715.000000000000,-516.000000000000,
-325.000000000000,-868.000000000000,
222.000000000000,-1320.00000000000,
947.000000000000,223.000000000000,
107.000000000000,210.000000000000,
-337.000000000000,383.000000000000,
517.000000000000,1156.00000000000,
-200.000000000000,-149.000000000000,
952.000000000000,-123.000000000000,
9.00000000000000,889.000000000000,
-1299.00000000000,-216.000000000000,
-517.000000000000,-839.000000000000,
-629.000000000000,-659.000000000000,
1162.00000000000,-211.000000000000,
643.000000000000,939.000000000000,
270.000000000000,182.000000000000,
393.000000000000,714.000000000000,
645.000000000000,1406.00000000000,
-227.000000000000,-62.0000000000000,
-1270.00000000000,786.000000000000,
739.000000000000,-62.0000000000000,
-248.000000000000,-220.000000000000,
36.0000000000000,1045.00000000000,
590.000000000000,2.00000000000000,
119.000000000000,907.000000000000,
470.000000000000,-68.0000000000000,
-260.000000000000,-224.000000000000,
375.000000000000,-772.000000000000,
695.000000000000,-568.000000000000,
-562.000000000000,589.000000000000,
-343.000000000000,-1121.00000000000,
321.000000000000,51.0000000000000,
-384.000000000000,312.000000000000,
-974.000000000000,921.000000000000,
-730.000000000000,-517.000000000000,
907.000000000000,-932.000000000000,
423.000000000000,659.000000000000,
499.000000000000,-1139.00000000000,
552.000000000000,-507.000000000000,
-663.000000000000,-164.000000000000,
708.000000000000,-586.000000000000,
767.000000000000,112.000000000000,
384.000000000000,688.000000000000,
-63.0000000000000,-577.000000000000,
-1057.00000000000,-707.000000000000,
438.000000000000,907.000000000000,
135.000000000000,-35.0000000000000,
-685.000000000000,164.000000000000,
776.000000000000,143.000000000000,
128.000000000000,-88.0000000000000,
410.000000000000,1058.00000000000,
225.000000000000,75.0000000000000,
654.000000000000,-290.000000000000,
-98.0000000000000,605.000000000000,
-681.000000000000,-423.000000000000,
895.000000000000,-586.000000000000,
-334.000000000000,-171.000000000000,
1057.00000000000,282.000000000000,
-426.000000000000,804.000000000000,
-576.000000000000,-520.000000000000,
640.000000000000,-251.000000000000,
-467.000000000000,-226.000000000000,
610.000000000000,-1246.00000000000,
-62.0000000000000,283.000000000000,
30.0000000000000,-333.000000000000,
-628.000000000000,-460.000000000000,
-137.000000000000,1119.00000000000,
470.000000000000,35.0000000000000,
-344.000000000000,722.000000000000,
-668.000000000000,41.0000000000000,
-751.000000000000,-401.000000000000,
-67.0000000000000,-891.000000000000,
-575.000000000000,-953.000000000000,
-294.000000000000,94.0000000000000,
314.000000000000,-1217.00000000000,
750.000000000000,680.000000000000,
243.000000000000,-649.000000000000,
-995.000000000000,260.000000000000,
-324.000000000000,233.000000000000,
-91.0000000000000,-1345.00000000000,
-55.0000000000000,1277.00000000000,
109.000000000000,-1343.00000000000,
1240.00000000000,-521.000000000000,
646.000000000000,1157.00000000000,
-807.000000000000,696.000000000000,
230.000000000000,388.000000000000,
-176.000000000000,241.000000000000,
592.000000000000,681.000000000000,
-550.000000000000,-104.000000000000,
-293.000000000000,226.000000000000,
341.000000000000,165.000000000000,
-1368.00000000000,582.000000000000,
456.000000000000,-217.000000000000,
289.000000000000,-298.000000000000,
-201.000000000000,700.000000000000,
-713.000000000000,453.000000000000,
-530.000000000000,-415.000000000000,
1192.00000000000,-1147.00000000000,
224.000000000000,294.000000000000,
-102.000000000000,-613.000000000000,
552.000000000000,-341.000000000000,
208.000000000000,1314.00000000000,
297.000000000000,-566.000000000000,
-476.000000000000,-392.000000000000,
-91.0000000000000,107.000000000000,
692.000000000000,-72.0000000000000,
-732.000000000000,-339.000000000000,
759.000000000000,-497.000000000000,
121.000000000000,-724.000000000000,
-876.000000000000,-626.000000000000,
310.000000000000,423.000000000000,
-564.000000000000,-602.000000000000,
72.0000000000000,228.000000000000,
340.000000000000,1269.00000000000,
-835.000000000000,167.000000000000,
-63.0000000000000,-111.000000000000,
605.000000000000,129.000000000000,
-199.000000000000,293.000000000000,
284.000000000000,293.000000000000,
640.000000000000,136.000000000000,
-443.000000000000,136.000000000000,
-637.000000000000,675.000000000000,
110.000000000000,-138.000000000000,
-545.000000000000,-1168.00000000000,
-2.00000000000000,-552.000000000000,
89.0000000000000,-123.000000000000,
-1051.00000000000,740.000000000000,
-35.0000000000000,729.000000000000,
156.000000000000,340.000000000000,
-146.000000000000,22.0000000000000,
-675.000000000000,-91.0000000000000,
202.000000000000,89.0000000000000,
-21.0000000000000,-642.000000000000,
-185.000000000000,-115.000000000000,
794.000000000000,-1066.00000000000,
-717.000000000000,-266.000000000000,
-391.000000000000,866.000000000000,
-257.000000000000,-1001.00000000000,
-68.0000000000000,-268.000000000000,
421.000000000000,365.000000000000,
485.000000000000,-630.000000000000,
1244.00000000000,57.0000000000000,
637.000000000000,168.000000000000,
-590.000000000000,180.000000000000,
-835.000000000000,223.000000000000,
-171.000000000000,-418.000000000000,
100.000000000000,607.000000000000,
-1.00000000000000,-388.000000000000,
-288.000000000000,-524.000000000000,
-611.000000000000,1117.00000000000,
168.000000000000,37.0000000000000,
673.000000000000,2.00000000000000,
142.000000000000,903.000000000000,
128.000000000000,236.000000000000,
315.000000000000,589.000000000000,
-599.000000000000,-656.000000000000,
-939.000000000000,-399.000000000000,
-582.000000000000,32.0000000000000,
-1314.00000000000,-498.000000000000,
624.000000000000,243.000000000000,
998.000000000000,-544.000000000000,
892.000000000000,295.000000000000,
883.000000000000,-415.000000000000,
-503.000000000000,-560.000000000000,
484.000000000000,-643.000000000000,
-901.000000000000,-1168.00000000000,
528.000000000000,-138.000000000000,
1289.00000000000,-504.000000000000,
224.000000000000,197.000000000000,
423.000000000000,-241.000000000000,
137.000000000000,-327.000000000000,
1367.00000000000,-118.000000000000,
-37.0000000000000,210.000000000000,
220.000000000000,424.000000000000,
876.000000000000,-191.000000000000,
77.0000000000000,403.000000000000,
-310.000000000000,-358.000000000000,
-677.000000000000,-716.000000000000,
-288.000000000000,-658.000000000000,
-948.000000000000,3.00000000000000,
2.00000000000000,384.000000000000,
314.000000000000,-945.000000000000,
862.000000000000,-294.000000000000,
61.0000000000000,518.000000000000,
-672.000000000000,208.000000000000,
1116.00000000000,-131.000000000000,
-517.000000000000,1096.00000000000,
-1170.00000000000,461.000000000000,
112.000000000000,-860.000000000000,
956.000000000000,459.000000000000,
-278.000000000000,72.0000000000000,
-942.000000000000,470.000000000000,
89.0000000000000,35.0000000000000,
-1218.00000000000,-409.000000000000,
-245.000000000000,-359.000000000000,
-514.000000000000,-1114.00000000000,
263.000000000000,-154.000000000000,
99.0000000000000,-349.000000000000,
-692.000000000000,-68.0000000000000,
579.000000000000,-912.000000000000,
-657.000000000000,-589.000000000000,
926.000000000000,-454.000000000000,
-291.000000000000,-440.000000000000,
158.000000000000,1253.00000000000,
426.000000000000,-383.000000000000,
-857.000000000000,184.000000000000,
1500.00000000000,-92.0000000000000,
-428.000000000000,-61.0000000000000,
-673.000000000000,219.000000000000,
-327.000000000000,-266.000000000000,
-286.000000000000,1110.00000000000,
-196.000000000000,-828.000000000000,
-197.000000000000,-935.000000000000,
590.000000000000,550.000000000000,
30.0000000000000,-260.000000000000,
-190.000000000000,-479.000000000000,
-383.000000000000,513.000000000000,
-297.000000000000,-20.0000000000000,
-788.000000000000,-1089.00000000000,
-145.000000000000,-798.000000000000,
58.0000000000000,-221.000000000000,
-945.000000000000,240.000000000000,
-159.000000000000,-260.000000000000,
3.00000000000000,-863.000000000000,
-197.000000000000,-425.000000000000,
-45.0000000000000,380.000000000000,
13.0000000000000,-524.000000000000,
-636.000000000000,-668.000000000000,
-6.00000000000000,-484.000000000000,
1001.00000000000,-140.000000000000,
-711.000000000000,-150.000000000000,
728.000000000000,-728.000000000000,
1063.00000000000,-24.0000000000000,
-44.0000000000000,-101.000000000000,
314.000000000000,325.000000000000,
-1335.00000000000,972.000000000000,
-195.000000000000,-648.000000000000,
664.000000000000,-623.000000000000,
118.000000000000,-402.000000000000,
-102.000000000000,-1009.00000000000,
-468.000000000000,752.000000000000,
67.0000000000000,724.000000000000,
375.000000000000,-288.000000000000,
496.000000000000,618.000000000000,
560.000000000000,746.000000000000,
-232.000000000000,964.000000000000,
-385.000000000000,353.000000000000,
1336.00000000000,-676.000000000000,
526.000000000000,330.000000000000,
-41.0000000000000,55.0000000000000,
107.000000000000,-196.000000000000,
-1523.00000000000,844.000000000000,
571.000000000000,-329.000000000000,
107.000000000000,-800.000000000000,
-308.000000000000,-370.000000000000,
863.000000000000,198.000000000000,
-1730.00000000000,1188.00000000000,
-869.000000000000,-697.000000000000,
16.0000000000000,-382.000000000000,
-325.000000000000,718.000000000000,
-884.000000000000,-646.000000000000,
-336.000000000000,554.000000000000,
1016.00000000000,-646.000000000000,
649.000000000000,-52.0000000000000,
187.000000000000,588.000000000000,
-21.0000000000000,-677.000000000000,
641.000000000000,-307.000000000000,
-1145.00000000000,-629.000000000000,
441.000000000000,-75.0000000000000,
356.000000000000,-52.0000000000000,
-992.000000000000,498.000000000000,
1316.00000000000,-544.000000000000,
-380.000000000000,-796.000000000000,
1097.00000000000,-325.000000000000,
363.000000000000,117.000000000000,
-199.000000000000,1255.00000000000,
679.000000000000,-301.000000000000,
186.000000000000,485.000000000000,
583.000000000000,1182.00000000000,
-1288.00000000000,476.000000000000,
435.000000000000,492.000000000000,
286.000000000000,271.000000000000,
550.000000000000,396.000000000000,
16.0000000000000,446.000000000000,
-673.000000000000,643.000000000000,
499.000000000000,612.000000000000,
-1109.00000000000,-197.000000000000,
937.000000000000,102.000000000000,
-449.000000000000,557.000000000000,
-758.000000000000,-1016.00000000000,
-291.000000000000,-532.000000000000,
-1008.00000000000,620.000000000000,
737.000000000000,-412.000000000000,
599.000000000000,485.000000000000,
1191.00000000000,278.000000000000,
367.000000000000,-794.000000000000,
708.000000000000,166.000000000000,
762.000000000000,-9.00000000000000,
51.0000000000000,270.000000000000,
742.000000000000,764.000000000000,
73.0000000000000,149.000000000000,
-207.000000000000,-556.000000000000,
-465.000000000000,470.000000000000,
-600.000000000000,577.000000000000,
-117.000000000000,-202.000000000000,
92.0000000000000,1043.00000000000,
66.0000000000000,585.000000000000,
-224.000000000000,-60.0000000000000,
-850.000000000000,384.000000000000,
49.0000000000000,-298.000000000000,
-123.000000000000,-255.000000000000,
-420.000000000000,270.000000000000,
73.0000000000000,543.000000000000,
-842.000000000000,478.000000000000,
-451.000000000000,50.0000000000000,
-130.000000000000,-872.000000000000,
-543.000000000000,-655.000000000000,
368.000000000000,-84.0000000000000,
357.000000000000,-186.000000000000,
-385.000000000000,385.000000000000,
-3.00000000000000,624.000000000000,
-179.000000000000,657.000000000000,
-489.000000000000,-1035.00000000000,
-263.000000000000,-350.000000000000,
167.000000000000,740.000000000000,
-276.000000000000,-1158.00000000000,
-41.0000000000000,-260.000000000000,
-524.000000000000,-467.000000000000,
-931.000000000000,-502.000000000000,
25.0000000000000,-270.000000000000,
-516.000000000000,-856.000000000000,
388.000000000000,-37.0000000000000,
-511.000000000000,-2.00000000000000,
-537.000000000000,-95.0000000000000,
974.000000000000,-824.000000000000,
-10.0000000000000,157.000000000000,
571.000000000000,93.0000000000000,
-491.000000000000,-1036.00000000000,
-586.000000000000,-474.000000000000,
452.000000000000,264.000000000000,
177.000000000000,-295.000000000000,
7.00000000000000,-1325.00000000000,
27.0000000000000,948.000000000000,
-249.000000000000,-186.000000000000,
263.000000000000,-185.000000000000,
856.000000000000,255.000000000000,
-602.000000000000,-796.000000000000,
-931.000000000000,980.000000000000,
-518.000000000000,-977.000000000000,
161.000000000000,423.000000000000,
392.000000000000,949.000000000000,
-894.000000000000,-412.000000000000,
587.000000000000,371.000000000000,
1175.00000000000,-508.000000000000,
158.000000000000,171.000000000000,
192.000000000000,-37.0000000000000,
-389.000000000000,-315.000000000000,
-516.000000000000,-35.0000000000000,
109.000000000000,-48.0000000000000,
-449.000000000000,-686.000000000000,
-596.000000000000,-1017.00000000000,
643.000000000000,-627.000000000000,
-98.0000000000000,-361.000000000000,
-351.000000000000,104.000000000000,
1138.00000000000,685.000000000000,
170.000000000000,686.000000000000,
-797.000000000000,-680.000000000000,
546.000000000000,-335.000000000000,
-427.000000000000,17.0000000000000,
-127.000000000000,-622.000000000000,
851.000000000000,616.000000000000,
-1086.00000000000,847.000000000000,
-417.000000000000,165.000000000000,
675.000000000000,-17.0000000000000,
776.000000000000,-731.000000000000,
872.000000000000,-77.0000000000000,
573.000000000000,904.000000000000,
375.000000000000,407.000000000000,
-549.000000000000,122.000000000000,
-779.000000000000,509.000000000000,
-257.000000000000,23.0000000000000,
-454.000000000000,373.000000000000,
274.000000000000,600.000000000000,
1179.00000000000,-326.000000000000,
-269.000000000000,644.000000000000,
-729.000000000000,634.000000000000,
628.000000000000,-368.000000000000,
878.000000000000,354.000000000000,
553.000000000000,901.000000000000,
-149.000000000000,735.000000000000,
-1003.00000000000,703.000000000000,
56.0000000000000,337.000000000000,
-37.0000000000000,-110.000000000000,
-568.000000000000,-1100.00000000000,
713.000000000000,-92.0000000000000,
751.000000000000,25.0000000000000,
989.000000000000,-49.0000000000000,
-217.000000000000,1025.00000000000,
-932.000000000000,-613.000000000000,
716.000000000000,379.000000000000,
480.000000000000,25.0000000000000,
84.0000000000000,-430.000000000000,
-361.000000000000,580.000000000000,
97.0000000000000,-116.000000000000,
-480.000000000000,415.000000000000,
747.000000000000,68.0000000000000,
374.000000000000,-134.000000000000,
-862.000000000000,-571.000000000000,
1474.00000000000,-206.000000000000,
-276.000000000000,583.000000000000,
13.0000000000000,614.000000000000,
574.000000000000,829.000000000000,
-488.000000000000,407.000000000000,
-744.000000000000,-516.000000000000,
-473.000000000000,-1432.00000000000,
630.000000000000,-137.000000000000,
-857.000000000000,478.000000000000,
-727.000000000000,-359.000000000000,
-993.000000000000,-106.000000000000,
-316.000000000000,-326.000000000000,
701.000000000000,-863.000000000000,
-829.000000000000,-397.000000000000,
395.000000000000,-936.000000000000,
812.000000000000,-249.000000000000,
-526.000000000000,347.000000000000,
128.000000000000,-788.000000000000,
1374.00000000000,348.000000000000,
347.000000000000,290.000000000000,
-626.000000000000,-741.000000000000,
531.000000000000,103.000000000000,
659.000000000000,535.000000000000,
-856.000000000000,235.000000000000,
-861.000000000000,612.000000000000,
-884.000000000000,233.000000000000,
-266.000000000000,-959.000000000000,
1211.00000000000,-633.000000000000,
-443.000000000000,-427.000000000000,
-632.000000000000,-865.000000000000,
747.000000000000,-645.000000000000,
-639.000000000000,-4.00000000000000,
250.000000000000,-297.000000000000,
1296.00000000000,-949.000000000000,
-414.000000000000,-198.000000000000,
42.0000000000000,214.000000000000,
-208.000000000000,918.000000000000,
-1023.00000000000,221.000000000000,
367.000000000000,-684.000000000000,
880.000000000000,924.000000000000,
-120.000000000000,677.000000000000,
387.000000000000,126.000000000000,
306.000000000000,-70.0000000000000,
-780.000000000000,-632.000000000000,
-137.000000000000,133.000000000000,
-62.0000000000000,-409.000000000000,
656.000000000000,-577.000000000000,
131.000000000000,771.000000000000,
151.000000000000,-116.000000000000,
444.000000000000,-212.000000000000,
-855.000000000000,391.000000000000,
-309.000000000000,-442.000000000000,
-907.000000000000,775.000000000000,
382.000000000000,606.000000000000,
697.000000000000,-844.000000000000,
73.0000000000000,860.000000000000,
220.000000000000,680.000000000000,
-1482.00000000000,747.000000000000,
209.000000000000,-333.000000000000,
-441.000000000000,-587.000000000000,
-1174.00000000000,91.0000000000000,
335.000000000000,-1326.00000000000,
920.000000000000,1373.00000000000,
-38.0000000000000,-163.000000000000,
-1062.00000000000,-75.0000000000000,
727.000000000000,-1.00000000000000,
643.000000000000,-240.000000000000,
421.000000000000,1583.00000000000,
29.0000000000000,-552.000000000000,
-331.000000000000,50.0000000000000,
-427.000000000000,-491.000000000000,
-389.000000000000,385.000000000000,
-289.000000000000,-233.000000000000,
-801.000000000000,-1553.00000000000,
1169.00000000000,305.000000000000,
-202.000000000000,-247.000000000000,
-963.000000000000,-743.000000000000,
193.000000000000,-938.000000000000,
-1034.00000000000,-610.000000000000,
-313.000000000000,-286.000000000000,
78.0000000000000,329.000000000000,
63.0000000000000,741.000000000000,
632.000000000000,252.000000000000,
322.000000000000,-296.000000000000,
-487.000000000000,-167.000000000000,
-323.000000000000,831.000000000000,
-370.000000000000,-362.000000000000,
-1178.00000000000,-351.000000000000,
-850.000000000000,210.000000000000,
-1082.00000000000,-102.000000000000,
-992.000000000000,440.000000000000,
124.000000000000,-1091.00000000000,
902.000000000000,-355.000000000000,
637.000000000000,647.000000000000,
220.000000000000,-181.000000000000,
615.000000000000,-913.000000000000,
-236.000000000000,-490.000000000000,
-136.000000000000,-17.0000000000000,
233.000000000000,-1228.00000000000,
389.000000000000,825.000000000000,
860.000000000000,548.000000000000,
-112.000000000000,297.000000000000,
661.000000000000,72.0000000000000,
190.000000000000,-436.000000000000,
-1130.00000000000,465.000000000000,
341.000000000000,-1427.00000000000,
504.000000000000,450.000000000000,
-164.000000000000,-437.000000000000,
76.0000000000000,-154.000000000000,
-125.000000000000,1405.00000000000,
-93.0000000000000,52.0000000000000,
637.000000000000,808.000000000000,
284.000000000000,-800.000000000000,
25.0000000000000,50.0000000000000,
-711.000000000000,585.000000000000,
-1396.00000000000,29.0000000000000,
-630.000000000000,407.000000000000,
-656.000000000000,237.000000000000,
742.000000000000,541.000000000000,
-36.0000000000000,-229.000000000000,
156.000000000000,-743.000000000000,
1066.00000000000,183.000000000000,
-631.000000000000,456.000000000000,
1029.00000000000,-616.000000000000,
-480.000000000000,617.000000000000,
-1526.00000000000,534.000000000000,
-372.000000000000,-1243.00000000000,
-372.000000000000,699.000000000000,
406.000000000000,634.000000000000,
-572.000000000000,815.000000000000,
-588.000000000000,-761.000000000000,
65.0000000000000,-811.000000000000,
1120.00000000000,934.000000000000,
-604.000000000000,-1156.00000000000,
-176.000000000000,533.000000000000,
978.000000000000,-321.000000000000,
-205.000000000000,84.0000000000000,
1094.00000000000,463.000000000000,
285.000000000000,36.0000000000000,
383.000000000000,1019.00000000000,
376.000000000000,-1019.00000000000,
369.000000000000,481.000000000000,
15.0000000000000,753.000000000000,
-1545.00000000000,597.000000000000,
10.0000000000000,-563.000000000000,
-175.000000000000,-965.000000000000,
-191.000000000000,260.000000000000,
663.000000000000,-545.000000000000,
930.000000000000,-1.00000000000000,
797.000000000000,212.000000000000,
-52.0000000000000,255.000000000000,
-143.000000000000,-798.000000000000,
95.0000000000000,-101.000000000000,
-302.000000000000,-241.000000000000,
-668.000000000000,-1257.00000000000,
-252.000000000000,734.000000000000,
-92.0000000000000,-87.0000000000000,
28.0000000000000,-195.000000000000,
-94.0000000000000,-136.000000000000,
-479.000000000000,125.000000000000,
-414.000000000000,493.000000000000,
426.000000000000,-786.000000000000,
865.000000000000,-439.000000000000,
457.000000000000,368.000000000000,
235.000000000000,841.000000000000,
431.000000000000,107.000000000000,
411.000000000000,136.000000000000,
-541.000000000000,335.000000000000,
262.000000000000,-150.000000000000,
83.0000000000000,373.000000000000,
-1162.00000000000,-15.0000000000000,
339.000000000000,127.000000000000,
279.000000000000,238.000000000000,
-672.000000000000,94.0000000000000,
400.000000000000,471.000000000000,
-1116.00000000000,437.000000000000,
-229.000000000000,34.0000000000000,
1245.00000000000,-400.000000000000,
-204.000000000000,78.0000000000000,
-42.0000000000000,147.000000000000,
-467.000000000000,-709.000000000000,
227.000000000000,-722.000000000000,
696.000000000000,358.000000000000,
-177.000000000000,335.000000000000,
-474.000000000000,-368.000000000000,
732.000000000000,550.000000000000,
477.000000000000,1224.00000000000,
-433.000000000000,27.0000000000000,
1210.00000000000,-548.000000000000,
319.000000000000,-389.000000000000,
664.000000000000,-458.000000000000,
-79.0000000000000,92.0000000000000,
-450.000000000000,914.000000000000,
713.000000000000,748.000000000000,
-636.000000000000,-632.000000000000,
905.000000000000,123.000000000000,
-227.000000000000,369.000000000000,
144.000000000000,-123.000000000000,
218.000000000000,713.000000000000,
-651.000000000000,-650.000000000000,
74.0000000000000,-947.000000000000,
-218.000000000000,-541.000000000000,
1226.00000000000,-478.000000000000,
444.000000000000,866.000000000000,
848.000000000000,927.000000000000,
220.000000000000,309.000000000000,
-72.0000000000000,193.000000000000,
743.000000000000,-121.000000000000,
-312.000000000000,-915.000000000000,
278.000000000000,77.0000000000000,
-863.000000000000,610.000000000000,
25.0000000000000,-565.000000000000,
-247.000000000000,-780.000000000000,
-430.000000000000,-508.000000000000,
1421.00000000000,-891.000000000000,
570.000000000000,202.000000000000,
-233.000000000000,585.000000000000,
-879.000000000000,-814.000000000000,
714.000000000000,-485.000000000000,
1205.00000000000,701.000000000000,
-57.0000000000000,464.000000000000,
64.0000000000000,-828.000000000000,
-3.00000000000000,126.000000000000,
-384.000000000000,129.000000000000,
-757.000000000000,-192.000000000000,
-416.000000000000,-54.0000000000000,
-708.000000000000,-488.000000000000,
-492.000000000000,701.000000000000,
-1296.00000000000,338.000000000000,
-858.000000000000,388.000000000000,
1032.00000000000,-22.0000000000000,
-153.000000000000,-271.000000000000,
-173.000000000000,-633.000000000000,
-96.0000000000000,-1487.00000000000,
-335.000000000000,640.000000000000,
-296.000000000000,264.000000000000,
-713.000000000000,-506.000000000000,
478.000000000000,490.000000000000,
465.000000000000,35.0000000000000,
188.000000000000,-133.000000000000,
-145.000000000000,309.000000000000,
-262.000000000000,-668.000000000000,
-267.000000000000,-955.000000000000,
-483.000000000000,833.000000000000,
-15.0000000000000,-298.000000000000,
731.000000000000,-883.000000000000,
950.000000000000,321.000000000000,
-757.000000000000,327.000000000000,
-70.0000000000000,58.0000000000000,
195.000000000000,-519.000000000000,
304.000000000000,-146.000000000000,
1049.00000000000,-333.000000000000,
-386.000000000000,-614.000000000000,
775.000000000000,1.00000000000000,
76.0000000000000,221.000000000000,
363.000000000000,944.000000000000,
384.000000000000,683.000000000000,
-559.000000000000,-528.000000000000,
848.000000000000,-729.000000000000,
159.000000000000,224.000000000000,
579.000000000000,670.000000000000,
-551.000000000000,508.000000000000,
2.00000000000000,356.000000000000,
1062.00000000000,763.000000000000,
-1062.00000000000,1115.00000000000,
-293.000000000000,-438.000000000000,
570.000000000000,515.000000000000,
-955.000000000000,983.000000000000,
-996.000000000000,-368.000000000000,
-322.000000000000,-1145.00000000000,
-335.000000000000,-1485.00000000000,
448.000000000000,467.000000000000,
68.0000000000000,-190.000000000000,
-100.000000000000,-90.0000000000000,
750.000000000000,1196.00000000000,
252.000000000000,273.000000000000,
-136.000000000000,-609.000000000000,
-589.000000000000,-1420.00000000000,
185.000000000000,-847.000000000000,
1089.00000000000,-820.000000000000,
-441.000000000000,718.000000000000,
-382.000000000000,-350.000000000000,
-170.000000000000,-811.000000000000,
-776.000000000000,541.000000000000,
88.0000000000000,-1145.00000000000,
-231.000000000000,405.000000000000,
-500.000000000000,-80.0000000000000,
-47.0000000000000,-1094.00000000000,
-679.000000000000,174.000000000000,
141.000000000000,342.000000000000,
1205.00000000000,445.000000000000,
-178.000000000000,1025.00000000000,
-460.000000000000,985.000000000000,
232.000000000000,-993.000000000000,
814.000000000000,356.000000000000,
820.000000000000,536.000000000000,
-846.000000000000,281.000000000000,
-688.000000000000,553.000000000000,
-840.000000000000,-1402.00000000000,
-326.000000000000,67.0000000000000,
1302.00000000000,417.000000000000,
258.000000000000,-284.000000000000,
-282.000000000000,183.000000000000,
-664.000000000000,320.000000000000,
389.000000000000,-415.000000000000,
255.000000000000,-1101.00000000000,
673.000000000000,-374.000000000000,
1502.00000000000,-831.000000000000,
702.000000000000,817.000000000000,
179.000000000000,-497.000000000000,
-971.000000000000,-366.000000000000,
422.000000000000,13.0000000000000,
184.000000000000,-1028.00000000000,
-1183.00000000000,798.000000000000,
271.000000000000,-1036.00000000000,
92.0000000000000,629.000000000000,
-278.000000000000,397.000000000000,
898.000000000000,-912.000000000000,
1105.00000000000,861.000000000000,
843.000000000000,431.000000000000,
-410.000000000000,1477.00000000000,
-536.000000000000,804.000000000000,
161.000000000000,-556.000000000000,
-48.0000000000000,-895.000000000000,
714.000000000000,-607.000000000000,
212.000000000000,-205.000000000000,
-178.000000000000,324.000000000000,
396.000000000000,204.000000000000,
-526.000000000000,-722.000000000000,
333.000000000000,-20.0000000000000,
1089.00000000000,-104.000000000000,
-582.000000000000,1120.00000000000,
-286.000000000000,390.000000000000,
-641.000000000000,-707.000000000000,
535.000000000000,317.000000000000,
911.000000000000,-826.000000000000,
-96.0000000000000,971.000000000000,
-105.000000000000,442.000000000000,
-726.000000000000,-65.0000000000000,
757.000000000000,1500.00000000000,
-1003.00000000000,100.000000000000,
-520.000000000000,-791.000000000000,
-14.0000000000000,-1424.00000000000,
-390.000000000000,-255.000000000000,
1312.00000000000,576.000000000000,
438.000000000000,-227.000000000000,
750.000000000000,146.000000000000,
-486.000000000000,915.000000000000,
-50.0000000000000,671.000000000000,
844.000000000000,-104.000000000000,
437.000000000000,88.0000000000000,
-15.0000000000000,744.000000000000,
-963.000000000000,152.000000000000,
59.0000000000000,-835.000000000000,
-219.000000000000,-176.000000000000,
295.000000000000,-200.000000000000,
675.000000000000,-261.000000000000,
-419.000000000000,55.0000000000000,
-131.000000000000,-756.000000000000,
78.0000000000000,969.000000000000,
-516.000000000000,-47.0000000000000,
686.000000000000,-930.000000000000,
1027.00000000000,618.000000000000,
-408.000000000000,-261.000000000000,
0.00000000000000,594.000000000000,
410.000000000000,863.000000000000,
-1036.00000000000,949.000000000000,
-948.000000000000,15.0000000000000,
209.000000000000,-1181.00000000000,
-168.000000000000,453.000000000000,
-590.000000000000,165.000000000000,
642.000000000000,-210.000000000000,
524.000000000000,852.000000000000,
-721.000000000000,238.000000000000,
-33.0000000000000,-1047.00000000000,
-2.00000000000000,-78.0000000000000,
276.000000000000,258.000000000000,
-38.0000000000000,301.000000000000,
-706.000000000000,655.000000000000,
-489.000000000000,-630.000000000000,
377.000000000000,485.000000000000,
190.000000000000,609.000000000000,
-1119.00000000000,-736.000000000000,
738.000000000000,-416.000000000000,
-114.000000000000,449.000000000000,
-612.000000000000,1054.00000000000,
290.000000000000,-410.000000000000,
-440.000000000000,289.000000000000,
-240.000000000000,300.000000000000,
-1042.00000000000,-55.0000000000000,
107.000000000000,498.000000000000,
-454.000000000000,-389.000000000000,
167.000000000000,669.000000000000,
-403.000000000000,461.000000000000,
-1366.00000000000,511.000000000000,
949.000000000000,23.0000000000000,
-229.000000000000,545.000000000000,
979.000000000000,61.0000000000000,
281.000000000000,-841.000000000000,
631.000000000000,881.000000000000,
663.000000000000,-661.000000000000,
-645.000000000000,249.000000000000,
696.000000000000,-422.000000000000,
-1084.00000000000,-744.000000000000,
-565.000000000000,1193.00000000000,
-1233.00000000000,-383.000000000000,
-679.000000000000,-710.000000000000,
137.000000000000,-790.000000000000,
-844.000000000000,-646.000000000000,
-67.0000000000000,-86.0000000000000,
483.000000000000,-12.0000000000000,
1335.00000000000,-124.000000000000,
610.000000000000,941.000000000000,
145.000000000000,681.000000000000,
-1000.00000000000,-723.000000000000,
-482.000000000000,101.000000000000,
517.000000000000,73.0000000000000,
-201.000000000000,-481.000000000000,
649.000000000000,-629.000000000000,
-129.000000000000,-345.000000000000,
327.000000000000,178.000000000000,
1216.00000000000,-95.0000000000000,
44.0000000000000,701.000000000000,
-488.000000000000,725.000000000000,
-755.000000000000,549.000000000000,
-609.000000000000,-480.000000000000,
-177.000000000000,-1390.00000000000,
867.000000000000,-479.000000000000,
-293.000000000000,-394.000000000000,
-545.000000000000,288.000000000000,
520.000000000000,22.0000000000000,
-162.000000000000,-321.000000000000,
147.000000000000,-810.000000000000,
295.000000000000,-344.000000000000,
170.000000000000,60.0000000000000,
-157.000000000000,-123.000000000000,
197.000000000000,903.000000000000,
756.000000000000,-701.000000000000,
416.000000000000,717.000000000000,
679.000000000000,1020.00000000000,
-437.000000000000,-718.000000000000,
-503.000000000000,-450.000000000000,
115.000000000000,-1292.00000000000,
-191.000000000000,674.000000000000,
-363.000000000000,316.000000000000,
-740.000000000000,-911.000000000000,
-237.000000000000,209.000000000000,
184.000000000000,916.000000000000,
-394.000000000000,254.000000000000,
-922.000000000000,-851.000000000000,
832.000000000000,-523.000000000000,
1186.00000000000,-606.000000000000,
14.0000000000000,360.000000000000,
1093.00000000000,-75.0000000000000,
462.000000000000,796.000000000000,
-209.000000000000,1207.00000000000,
144.000000000000,-788.000000000000,
-638.000000000000,-812.000000000000,
522.000000000000,-908.000000000000,
463.000000000000,945.000000000000,
-1071.00000000000,-357.000000000000,
-1.00000000000000,-382.000000000000,
425.000000000000,905.000000000000,
-657.000000000000,-495.000000000000,
-323.000000000000,518.000000000000,
411.000000000000,-879.000000000000,
803.000000000000,176.000000000000,
32.0000000000000,658.000000000000,
-975.000000000000,-443.000000000000,
720.000000000000,351.000000000000,
46.0000000000000,-196.000000000000,
-91.0000000000000,-66.0000000000000,
-104.000000000000,44.0000000000000,
-1099.00000000000,658.000000000000,
-61.0000000000000,-435.000000000000,
-799.000000000000,-865.000000000000,
76.0000000000000,-1272.00000000000,
295.000000000000,-1115.00000000000,
1190.00000000000,190.000000000000,
484.000000000000,-836.000000000000,
-509.000000000000,207.000000000000,
445.000000000000,-976.000000000000,
-862.000000000000,-196.000000000000,
279.000000000000,786.000000000000,
-869.000000000000,-198.000000000000,
-736.000000000000,1021.00000000000,
796.000000000000,-12.0000000000000,
-327.000000000000,990.000000000000,
-659.000000000000,122.000000000000,
-327.000000000000,-1232.00000000000,
1049.00000000000,1006.00000000000,
482.000000000000,440.000000000000,
360.000000000000,-11.0000000000000,
-245.000000000000,646.000000000000,
347.000000000000,49.0000000000000,
474.000000000000,289.000000000000,
-1141.00000000000,149.000000000000,
69.0000000000000,-1668.00000000000,
-766.000000000000,-461.000000000000,
120.000000000000,290.000000000000,
1121.00000000000,-739.000000000000,
465.000000000000,271.000000000000,
355.000000000000,849.000000000000,
-611.000000000000,1316.00000000000,
-748.000000000000,63.0000000000000,
-1076.00000000000,-679.000000000000,
203.000000000000,214.000000000000,
276.000000000000,-650.000000000000,
-327.000000000000,481.000000000000,
29.0000000000000,553.000000000000,
-514.000000000000,-368.000000000000,
122.000000000000,189.000000000000,
293.000000000000,1067.00000000000,
-641.000000000000,471.000000000000,
-986.000000000000,-1624.00000000000,
578.000000000000,-894.000000000000,
356.000000000000,39.0000000000000,
-1401.00000000000,153.000000000000,
-200.000000000000,-1005.00000000000,
693.000000000000,-940.000000000000,
1628.00000000000,-28.0000000000000,
-136.000000000000,-273.000000000000,
-788.000000000000,958.000000000000,
-62.0000000000000,654.000000000000,
67.0000000000000,581.000000000000,
825.000000000000,112.000000000000,
-732.000000000000,-697.000000000000,
468.000000000000,-595.000000000000,
-284.000000000000,-940.000000000000,
-152.000000000000,-467.000000000000,
544.000000000000,-942.000000000000,
-896.000000000000,-275.000000000000,
689.000000000000,982.000000000000,
-549.000000000000,5.00000000000000,
-635.000000000000,-1146.00000000000,
651.000000000000,-1123.00000000000,
-145.000000000000,-436.000000000000,
526.000000000000,-2.00000000000000,
635.000000000000,-423.000000000000,
-122.000000000000,-519.000000000000,
700.000000000000,1000.00000000000,
81.0000000000000,546.000000000000,
-127.000000000000,-420.000000000000,
55.0000000000000,566.000000000000,
-592.000000000000,340.000000000000,
-134.000000000000,214.000000000000,
-75.0000000000000,-300.000000000000,
513.000000000000,-847.000000000000,
1202.00000000000,21.0000000000000,
741.000000000000,695.000000000000,
-171.000000000000,92.0000000000000,
-718.000000000000,-740.000000000000,
221.000000000000,-880.000000000000,
303.000000000000,-429.000000000000,
-687.000000000000,524.000000000000,
358.000000000000,77.0000000000000,
-655.000000000000,-235.000000000000,
-827.000000000000,29.0000000000000,
-478.000000000000,-1582.00000000000,
-37.0000000000000,-596.000000000000,
1690.00000000000,-223.000000000000,
-94.0000000000000,-392.000000000000,
-341.000000000000,312.000000000000,
46.0000000000000,372.000000000000,
246.000000000000,141.000000000000,
136.000000000000,-907.000000000000,
-725.000000000000,262.000000000000,
144.000000000000,-920.000000000000,
218.000000000000,-142.000000000000,
703.000000000000,776.000000000000,
466.000000000000,692.000000000000,
-943.000000000000,1008.00000000000,
-200.000000000000,-617.000000000000,
1034.00000000000,1126.00000000000,
640.000000000000,-336.000000000000,
-206.000000000000,-56.0000000000000,
-921.000000000000,713.000000000000,
-344.000000000000,-358.000000000000,
203.000000000000,1056.00000000000,
-859.000000000000,-294.000000000000,
-75.0000000000000,-802.000000000000,
1418.00000000000,-314.000000000000,
81.0000000000000,576.000000000000,
-40.0000000000000,662.000000000000,
54.0000000000000,569.000000000000,
-530.000000000000,737.000000000000,
-257.000000000000,-256.000000000000,
-199.000000000000,-415.000000000000,
-444.000000000000,-944.000000000000,
-346.000000000000,-323.000000000000,
-189.000000000000,328.000000000000,
74.0000000000000,-189.000000000000,
501.000000000000,-334.000000000000,
-775.000000000000,349.000000000000,
-125.000000000000,1192.00000000000,
-16.0000000000000,15.0000000000000,
-1243.00000000000,450.000000000000,
349.000000000000,688.000000000000,
50.0000000000000,750.000000000000,
518.000000000000,793.000000000000,
482.000000000000,-548.000000000000,
-36.0000000000000,-398.000000000000,
443.000000000000,-879.000000000000,
-763.000000000000,427.000000000000,
-466.000000000000,440.000000000000,
194.000000000000,46.0000000000000,
268.000000000000,578.000000000000,
-943.000000000000,-160.000000000000,
-567.000000000000,878.000000000000,
0.00000000000000,-505.000000000000,
175.000000000000,-305.000000000000,
1007.00000000000,15.0000000000000,
-321.000000000000,-442.000000000000,
1101.00000000000,239.000000000000,
-162.000000000000,-78.0000000000000,
-1006.00000000000,842.000000000000,
578.000000000000,714.000000000000,
-5.00000000000000,107.000000000000,
-361.000000000000,-478.000000000000,
-619.000000000000,-587.000000000000,
305.000000000000,-820.000000000000,
-199.000000000000,239.000000000000,
633.000000000000,1023.00000000000,
641.000000000000,-655.000000000000,
-146.000000000000,802.000000000000,
863.000000000000,-319.000000000000,
-572.000000000000,-342.000000000000,
399.000000000000,1239.00000000000,
729.000000000000,-541.000000000000,
-402.000000000000,-189.000000000000,
-483.000000000000,217.000000000000,
-956.000000000000,518.000000000000,
-84.0000000000000,-692.000000000000,
1028.00000000000,-491.000000000000,
1023.00000000000,823.000000000000,
-142.000000000000,337.000000000000,
-171.000000000000,-209.000000000000,
-322.000000000000,-1050.00000000000,
522.000000000000,304.000000000000,
749.000000000000,640.000000000000,
273.000000000000,205.000000000000,
1426.00000000000,-177.000000000000,
-517.000000000000,-229.000000000000,
54.0000000000000,391.000000000000,
-73.0000000000000,-459.000000000000,
-404.000000000000,-332.000000000000,
1604.00000000000,209.000000000000,
-93.0000000000000,-117.000000000000,
-88.0000000000000,-671.000000000000,
-138.000000000000,-998.000000000000,
449.000000000000,-654.000000000000,
1201.00000000000,134.000000000000,
-190.000000000000,1357.00000000000,
-479.000000000000,842.000000000000,
417.000000000000,639.000000000000,
739.000000000000,543.000000000000,
-161.000000000000,980.000000000000,
740.000000000000,675.000000000000,
428.000000000000,-709.000000000000,
-682.000000000000,535.000000000000,
-926.000000000000,-642.000000000000,
-732.000000000000,-735.000000000000,
807.000000000000,402.000000000000,
-152.000000000000,1029.00000000000,
-106.000000000000,824.000000000000,
-115.000000000000,-1146.00000000000,
95.0000000000000,620.000000000000,
-218.000000000000,231.000000000000,
-1190.00000000000,-633.000000000000,
722.000000000000,-439.000000000000,
186.000000000000,463.000000000000,
314.000000000000,779.000000000000,
29.0000000000000,-414.000000000000,
-314.000000000000,1123.00000000000,
924.000000000000,410.000000000000,
-112.000000000000,169.000000000000,
30.0000000000000,829.000000000000,
-407.000000000000,224.000000000000,
-1025.00000000000,-427.000000000000,
460.000000000000,-601.000000000000,
201.000000000000,449.000000000000,
-512.000000000000,-598.000000000000,
633.000000000000,-772.000000000000,
-460.000000000000,-399.000000000000,
-945.000000000000,-526.000000000000,
340.000000000000,-392.000000000000,
-905.000000000000,362.000000000000,
-224.000000000000,900.000000000000,
346.000000000000,15.0000000000000,
-1087.00000000000,-201.000000000000,
121.000000000000,-1393.00000000000,
174.000000000000,-326.000000000000,
-606.000000000000,511.000000000000,
-228.000000000000,174.000000000000,
-742.000000000000,817.000000000000,
185.000000000000,-799.000000000000,
196.000000000000,-541.000000000000,
-275.000000000000,-693.000000000000,
696.000000000000,174.000000000000,
-317.000000000000,174.000000000000,
-186.000000000000,-763.000000000000,
-318.000000000000,879.000000000000,
-1147.00000000000,-857.000000000000,
-529.000000000000,-840.000000000000,
-251.000000000000,-623.000000000000,
-145.000000000000,-1097.00000000000,
572.000000000000,-626.000000000000,
1112.00000000000,-233.000000000000,
702.000000000000,-311.000000000000,
646.000000000000,-442.000000000000,
445.000000000000,1289.00000000000,
161.000000000000,-143.000000000000,
-249.000000000000,-55.0000000000000,
-653.000000000000,275.000000000000,
-502.000000000000,-579.000000000000,
779.000000000000,544.000000000000,
691.000000000000,252.000000000000,
235.000000000000,1417.00000000000,
155.000000000000,583.000000000000,
-611.000000000000,263.000000000000,
917.000000000000,-198.000000000000,
249.000000000000,-400.000000000000,
-928.000000000000,689.000000000000,
-7.00000000000000,-1008.00000000000,
-112.000000000000,422.000000000000,
670.000000000000,482.000000000000,
506.000000000000,-145.000000000000,
-119.000000000000,-590.000000000000,
-155.000000000000,-800.000000000000,
-335.000000000000,-765.000000000000,
1041.00000000000,-917.000000000000,
-207.000000000000,1310.00000000000,
-600.000000000000,-312.000000000000,
950.000000000000,-164.000000000000,
-214.000000000000,-82.0000000000000,
653.000000000000,-140.000000000000,
1010.00000000000,1597.00000000000,
-68.0000000000000,957.000000000000,
189.000000000000,745.000000000000,
48.0000000000000,-557.000000000000,
-616.000000000000,464.000000000000,
-650.000000000000,-164.000000000000,
-400.000000000000,-282.000000000000,
-488.000000000000,423.000000000000,
-968.000000000000,-1216.00000000000,
24.0000000000000,881.000000000000,
6.00000000000000,479.000000000000,
-1262.00000000000,608.000000000000,
1177.00000000000,-31.0000000000000,
1066.00000000000,-547.000000000000,
-325.000000000000,592.000000000000,
-154.000000000000,-162.000000000000,
102.000000000000,681.000000000000,
-212.000000000000,-699.000000000000,
-1090.00000000000,69.0000000000000,
-368.000000000000,-640.000000000000,
-497.000000000000,-292.000000000000,
189.000000000000,1230.00000000000,
-875.000000000000,-222.000000000000,
-179.000000000000,1158.00000000000,
-46.0000000000000,254.000000000000,
-1649.00000000000,532.000000000000,
76.0000000000000,-244.000000000000,
-532.000000000000,-1335.00000000000,
510.000000000000,-881.000000000000,
1229.00000000000,-689.000000000000,
-366.000000000000,424.000000000000,
191.000000000000,-748.000000000000,
759.000000000000,600.000000000000,
973.000000000000,409.000000000000,
337.000000000000,306.000000000000,
-362.000000000000,910.000000000000,
216.000000000000,405.000000000000,
-454.000000000000,291.000000000000,
-562.000000000000,-978.000000000000,
209.000000000000,823.000000000000,
613.000000000000,266.000000000000,
730.000000000000,-267.000000000000,
-514.000000000000,137.000000000000,
108.000000000000,-913.000000000000,
377.000000000000,-337.000000000000,
-842.000000000000,-373.000000000000,
-270.000000000000,-58.0000000000000,
-734.000000000000,382.000000000000,
-915.000000000000,-841.000000000000,
466.000000000000,-595.000000000000,
692.000000000000,149.000000000000,
513.000000000000,-285.000000000000,
-457.000000000000,146.000000000000,
86.0000000000000,-408.000000000000,
133.000000000000,-482.000000000000,
-670.000000000000,405.000000000000,
1017.00000000000,-96.0000000000000,
-152.000000000000,452.000000000000,
252.000000000000,640.000000000000,
452.000000000000,-798.000000000000,
-1380.00000000000,-375.000000000000,
314.000000000000,-505.000000000000,
-119.000000000000,-298.000000000000,
-869.000000000000,250.000000000000,
52.0000000000000,539.000000000000,
413.000000000000,1309.00000000000,
592.000000000000,307.000000000000,
160.000000000000,118.000000000000,
-308.000000000000,-389.000000000000,
365.000000000000,149.000000000000,
508.000000000000,216.000000000000,
16.0000000000000,-71.0000000000000,
-20.0000000000000,563.000000000000,
-844.000000000000,194.000000000000,
-374.000000000000,673.000000000000,
976.000000000000,408.000000000000,
233.000000000000,197.000000000000,
-457.000000000000,-673.000000000000,
-622.000000000000,-451.000000000000,
-810.000000000000,651.000000000000,
123.000000000000,149.000000000000,
128.000000000000,238.000000000000,
-310.000000000000,-285.000000000000,
39.0000000000000,-118.000000000000,
-365.000000000000,-8.00000000000000,
-597.000000000000,-205.000000000000,
234.000000000000,-254.000000000000,
-153.000000000000,2.00000000000000,
-960.000000000000,784.000000000000,
354.000000000000,-1023.00000000000,
357.000000000000,-744.000000000000,
-226.000000000000,-163.000000000000,
1169.00000000000,-924.000000000000,
1266.00000000000,256.000000000000,
532.000000000000,603.000000000000,
573.000000000000,243.000000000000,
-250.000000000000,328.000000000000,
-571.000000000000,-415.000000000000,
-72.0000000000000,-768.000000000000,
-76.0000000000000,-916.000000000000,
-356.000000000000,-280.000000000000,
-195.000000000000,724.000000000000,
-521.000000000000,144.000000000000,
-178.000000000000,699.000000000000,
288.000000000000,720.000000000000,
-166.000000000000,725.000000000000,
505.000000000000,738.000000000000,
42.0000000000000,-629.000000000000,
-102.000000000000,-981.000000000000,
-229.000000000000,-1023.00000000000,
-401.000000000000,-84.0000000000000,
-48.0000000000000,301.000000000000,
-137.000000000000,-1181.00000000000,
362.000000000000,-38.0000000000000,
540.000000000000,129.000000000000,
46.0000000000000,-713.000000000000,
580.000000000000,1236.00000000000,
27.0000000000000,-141.000000000000,
-298.000000000000,-509.000000000000,
847.000000000000,957.000000000000,
292.000000000000,14.0000000000000,
184.000000000000,-486.000000000000,
-441.000000000000,324.000000000000,
381.000000000000,1048.00000000000,
452.000000000000,-231.000000000000,
140.000000000000,-596.000000000000,
698.000000000000,-704.000000000000,
-180.000000000000,-1175.00000000000,
806.000000000000,403.000000000000,
-472.000000000000,737.000000000000,
-957.000000000000,-471.000000000000,
31.0000000000000,112.000000000000,
44.0000000000000,557.000000000000,
369.000000000000,-623.000000000000,
-238.000000000000,-210.000000000000,
-413.000000000000,-22.0000000000000,
-470.000000000000,-585.000000000000,
979.000000000000,-3.00000000000000,
756.000000000000,-592.000000000000,
-265.000000000000,-103.000000000000,
785.000000000000,140.000000000000,
529.000000000000,36.0000000000000,
551.000000000000,-848.000000000000,
-125.000000000000,-481.000000000000,
-423.000000000000,507.000000000000,
466.000000000000,-1155.00000000000,
1256.00000000000,89.0000000000000,
-49.0000000000000,331.000000000000,
-653.000000000000,-603.000000000000,
757.000000000000,565.000000000000,
-632.000000000000,-333.000000000000,
99.0000000000000,-373.000000000000,
330.000000000000,548.000000000000,
416.000000000000,-323.000000000000,
1152.00000000000,-287.000000000000,
414.000000000000,-29.0000000000000,
851.000000000000,-371.000000000000,
-338.000000000000,-859.000000000000,
-293.000000000000,-823.000000000000,
-28.0000000000000,-164.000000000000,
428.000000000000,-214.000000000000,
627.000000000000,-344.000000000000,
-254.000000000000,688.000000000000,
328.000000000000,-510.000000000000,
-513.000000000000,-1033.00000000000,
-330.000000000000,-222.000000000000,
-397.000000000000,-871.000000000000,
346.000000000000,5.00000000000000,
1073.00000000000,123.000000000000,
-259.000000000000,1129.00000000000,
122.000000000000,711.000000000000,
186.000000000000,223.000000000000,
-185.000000000000,1419.00000000000,
-527.000000000000,-249.000000000000,
-587.000000000000,-1084.00000000000,
-301.000000000000,-33.0000000000000,
-426.000000000000,957.000000000000,
-386.000000000000,418.000000000000,
-208.000000000000,-193.000000000000,
-43.0000000000000,-647.000000000000,
-782.000000000000,-1382.00000000000,
719.000000000000,-755.000000000000,
-263.000000000000,293.000000000000,
-1179.00000000000,728.000000000000,
672.000000000000,-650.000000000000,
-739.000000000000,-113.000000000000,
482.000000000000,545.000000000000,
1325.00000000000,-655.000000000000,
636.000000000000,651.000000000000,
1010.00000000000,597.000000000000,
330.000000000000,193.000000000000,
-121.000000000000,-163.000000000000,
-169.000000000000,-807.000000000000,
984.000000000000,371.000000000000,
-215.000000000000,801.000000000000,
-525.000000000000,662.000000000000,
-203.000000000000,291.000000000000,
-308.000000000000,-386.000000000000,
-337.000000000000,-73.0000000000000,
-1241.00000000000,529.000000000000,
-440.000000000000,-507.000000000000,
-406.000000000000,-384.000000000000,
-499.000000000000,463.000000000000,
-790.000000000000,-995.000000000000,
-304.000000000000,-789.000000000000,
271.000000000000,-312.000000000000,
-575.000000000000,-886.000000000000,
640.000000000000,-970.000000000000,
711.000000000000,213.000000000000,
749.000000000000,1170.00000000000,
230.000000000000,-699.000000000000,
-740.000000000000,-517.000000000000,
88.0000000000000,246.000000000000,
-121.000000000000,-228.000000000000,
293.000000000000,-865.000000000000,
-159.000000000000,377.000000000000,
361.000000000000,926.000000000000,
150.000000000000,-611.000000000000,
-610.000000000000,605.000000000000,
-430.000000000000,-1322.00000000000,
-243.000000000000,-913.000000000000,
881.000000000000,839.000000000000,
-627.000000000000,-805.000000000000,
582.000000000000,-17.0000000000000,
533.000000000000,579.000000000000,
-180.000000000000,1084.00000000000,
29.0000000000000,287.000000000000,
-983.000000000000,135.000000000000,
471.000000000000,764.000000000000,
-1057.00000000000,-193.000000000000,
-743.000000000000,-220.000000000000,
-763.000000000000,-306.000000000000,
-368.000000000000,-1087.00000000000,
1403.00000000000,-923.000000000000,
127.000000000000,1243.00000000000,
270.000000000000,145.000000000000,
-503.000000000000,-386.000000000000,
-992.000000000000,529.000000000000,
-53.0000000000000,-1606.00000000000,
1075.00000000000,-426.000000000000,
1203.00000000000,986.000000000000,
139.000000000000,951.000000000000,
-412.000000000000,803.000000000000,
-1015.00000000000,-290.000000000000,
-198.000000000000,-1009.00000000000,
148.000000000000,-928.000000000000,
182.000000000000,-349.000000000000,
-726.000000000000,222.000000000000,
-668.000000000000,921.000000000000,
681.000000000000,566.000000000000,
185.000000000000,327.000000000000,
149.000000000000,445.000000000000,
-986.000000000000,-347.000000000000,
49.0000000000000,312.000000000000,
674.000000000000,761.000000000000,
-316.000000000000,68.0000000000000,
26.0000000000000,234.000000000000,
-1001.00000000000,447.000000000000,
485.000000000000,-377.000000000000,
277.000000000000,-933.000000000000,
-55.0000000000000,-128.000000000000,
988.000000000000,-15.0000000000000,
334.000000000000,135.000000000000,
-199.000000000000,356.000000000000,
-328.000000000000,539.000000000000,
942.000000000000,277.000000000000,
380.000000000000,-737.000000000000,
1005.00000000000,-45.0000000000000,
-125.000000000000,455.000000000000,
-876.000000000000,-86.0000000000000,
779.000000000000,-292.000000000000,
-163.000000000000,-662.000000000000,
-191.000000000000,235.000000000000,
704.000000000000,-14.0000000000000,
915.000000000000,-17.0000000000000,
371.000000000000,1477.00000000000,
45.0000000000000,-138.000000000000,
-264.000000000000,48.0000000000000,
-754.000000000000,687.000000000000,
-398.000000000000,-1390.00000000000,
-371.000000000000,-503.000000000000,
-2.00000000000000,745.000000000000,
188.000000000000,-6.00000000000000,
-232.000000000000,688.000000000000,
-475.000000000000,59.0000000000000,
-453.000000000000,-24.0000000000000,
524.000000000000,-584.000000000000,
221.000000000000,-513.000000000000,
-500.000000000000,962.000000000000,
-536.000000000000,-498.000000000000,
57.0000000000000,139.000000000000,
1227.00000000000,-351.000000000000,
977.000000000000,-253.000000000000,
444.000000000000,617.000000000000,
-441.000000000000,-195.000000000000,
-42.0000000000000,782.000000000000,
208.000000000000,294.000000000000,
-281.000000000000,-682.000000000000,
-268.000000000000,-383.000000000000,
-35.0000000000000,-183.000000000000,
1037.00000000000,115.000000000000,
765.000000000000,385.000000000000,
251.000000000000,-190.000000000000,
-372.000000000000,-948.000000000000,
-653.000000000000,-965.000000000000,
-379.000000000000,-32.0000000000000,
-236.000000000000,1259.00000000000,
-258.000000000000,48.0000000000000,
-856.000000000000,-601.000000000000,
-260.000000000000,323.000000000000,
-483.000000000000,-769.000000000000,
481.000000000000,-292.000000000000,
103.000000000000,574.000000000000,
-823.000000000000,-548.000000000000,
996.000000000000,-361.000000000000,
46.0000000000000,-102.000000000000,
605.000000000000,515.000000000000,
607.000000000000,970.000000000000,
-297.000000000000,-191.000000000000,
-633.000000000000,-376.000000000000,
-526.000000000000,493.000000000000,
545.000000000000,688.000000000000,
85.0000000000000,-375.000000000000,
726.000000000000,56.0000000000000,
18.0000000000000,685.000000000000,
382.000000000000,-241.000000000000,
1248.00000000000,-339.000000000000,
115.000000000000,721.000000000000,
59.0000000000000,439.000000000000,
-526.000000000000,969.000000000000,
544.000000000000,763.000000000000,
62.0000000000000,-1073.00000000000,
293.000000000000,-417.000000000000,
265.000000000000,-685.000000000000,
-396.000000000000,700.000000000000,
812.000000000000,881.000000000000,
61.0000000000000,-81.0000000000000,
789.000000000000,190.000000000000,
328.000000000000,-486.000000000000,
644.000000000000,-49.0000000000000,
-216.000000000000,-489.000000000000,
-1052.00000000000,666.000000000000,
925.000000000000,690.000000000000,
-663.000000000000,752.000000000000,
-1017.00000000000,430.000000000000,
-761.000000000000,-1216.00000000000,
8.00000000000000,-270.000000000000,
1651.00000000000,-579.000000000000,
-18.0000000000000,-745.000000000000,
-18.0000000000000,-32.0000000000000,
553.000000000000,142.000000000000,
-773.000000000000,-377.000000000000,
523.000000000000,92.0000000000000,
289.000000000000,630.000000000000,
-541.000000000000,297.000000000000,
-1.00000000000000,619.000000000000,
-832.000000000000,-249.000000000000,
333.000000000000,-216.000000000000,
796.000000000000,274.000000000000,
-256.000000000000,535.000000000000,
-227.000000000000,187.000000000000,
-572.000000000000,-308.000000000000,
-330.000000000000,227.000000000000,
371.000000000000,-884.000000000000,
-277.000000000000,-623.000000000000,
366.000000000000,-326.000000000000,
1129.00000000000,-923.000000000000,
602.000000000000,50.0000000000000,
-283.000000000000,-254.000000000000,
-179.000000000000,-576.000000000000,
1118.00000000000,15.0000000000000,
553.000000000000,486.000000000000,
322.000000000000,-450.000000000000,
432.000000000000,538.000000000000,
-50.0000000000000,220.000000000000,
-590.000000000000,-1355.00000000000,
-136.000000000000,728.000000000000,
346.000000000000,-992.000000000000,
-1163.00000000000,66.0000000000000,
-599.000000000000,168.000000000000,
-297.000000000000,-1024.00000000000,
-429.000000000000,840.000000000000,
831.000000000000,-849.000000000000,
917.000000000000,-235.000000000000,
798.000000000000,320.000000000000,
73.0000000000000,-425.000000000000,
284.000000000000,-1087.00000000000,
803.000000000000,-236.000000000000,
-185.000000000000,144.000000000000,
-696.000000000000,-366.000000000000,
-159.000000000000,782.000000000000,
-448.000000000000,-375.000000000000,
-109.000000000000,193.000000000000,
282.000000000000,1219.00000000000,
-777.000000000000,-170.000000000000,
292.000000000000,-744.000000000000,
-54.0000000000000,-400.000000000000,
69.0000000000000,-499.000000000000,
787.000000000000,-1003.00000000000,
-249.000000000000,-352.000000000000,
-141.000000000000,-963.000000000000,
-885.000000000000,-156.000000000000,
663.000000000000,818.000000000000,
513.000000000000,-502.000000000000,
-490.000000000000,-100.000000000000,
731.000000000000,-507.000000000000,
34.0000000000000,329.000000000000,
-37.0000000000000,-241.000000000000,
694.000000000000,-768.000000000000,
867.000000000000,88.0000000000000,
-914.000000000000,-386.000000000000,
-12.0000000000000,888.000000000000,
810.000000000000,228.000000000000,
-247.000000000000,92.0000000000000,
723.000000000000,481.000000000000,
209.000000000000,568.000000000000,
173.000000000000,-390.000000000000,
581.000000000000,-717.000000000000,
854.000000000000,753.000000000000,
199.000000000000,617.000000000000,
-809.000000000000,1066.00000000000,
-428.000000000000,-88.0000000000000,
-78.0000000000000,169.000000000000,
753.000000000000,934.000000000000,
-631.000000000000,-464.000000000000,
-690.000000000000,-1011.00000000000,
635.000000000000,-1160.00000000000,
-324.000000000000,391.000000000000,
-896.000000000000,-383.000000000000,
-565.000000000000,149.000000000000,
-4.00000000000000,1035.00000000000,
-1186.00000000000,229.000000000000,
-799.000000000000,-33.0000000000000,
-280.000000000000,-763.000000000000,
-791.000000000000,673.000000000000,
76.0000000000000,-1121.00000000000,
-771.000000000000,-357.000000000000,
249.000000000000,-18.0000000000000,
581.000000000000,-762.000000000000,
-198.000000000000,1814.00000000000,
-244.000000000000,213.000000000000,
140.000000000000,406.000000000000,
206.000000000000,346.000000000000,
-749.000000000000,176.000000000000,
-388.000000000000,-509.000000000000,
-1195.00000000000,-457.000000000000,
458.000000000000,510.000000000000,
860.000000000000,-792.000000000000,
-553.000000000000,777.000000000000,
273.000000000000,-774.000000000000,
153.000000000000,-1085.00000000000,
147.000000000000,777.000000000000,
-494.000000000000,-761.000000000000,
287.000000000000,-510.000000000000,
-586.000000000000,611.000000000000,
-470.000000000000,680.000000000000,
709.000000000000,219.000000000000,
422.000000000000,500.000000000000,
437.000000000000,268.000000000000,
-877.000000000000,-996.000000000000,
311.000000000000,-923.000000000000,
37.0000000000000,-1447.00000000000,
-74.0000000000000,-1016.00000000000,
122.000000000000,754.000000000000,
-366.000000000000,-294.000000000000,
1201.00000000000,453.000000000000,
714.000000000000,690.000000000000,
-401.000000000000,-622.000000000000,
28.0000000000000,625.000000000000,
1031.00000000000,175.000000000000,
-454.000000000000,347.000000000000,
-1097.00000000000,571.000000000000,
559.000000000000,-407.000000000000,
342.000000000000,584.000000000000,
-90.0000000000000,977.000000000000,
428.000000000000,-62.0000000000000,
21.0000000000000,194.000000000000,
-121.000000000000,252.000000000000,
-381.000000000000,118.000000000000,
-1111.00000000000,192.000000000000,
-547.000000000000,-115.000000000000,
274.000000000000,-223.000000000000,
693.000000000000,234.000000000000,
640.000000000000,426.000000000000,
325.000000000000,-617.000000000000,
553.000000000000,-354.000000000000,
625.000000000000,305.000000000000,
-172.000000000000,-75.0000000000000,
-776.000000000000,-112.000000000000,
-752.000000000000,109.000000000000,
-745.000000000000,-38.0000000000000,
-539.000000000000,70.0000000000000,
-506.000000000000,399.000000000000,
-217.000000000000,-781.000000000000,
-193.000000000000,-339.000000000000,
-73.0000000000000,-140.000000000000,
217.000000000000,-1107.00000000000,
-438.000000000000,14.0000000000000,
-641.000000000000,294.000000000000,
281.000000000000,-419.000000000000,
385.000000000000,-963.000000000000,
763.000000000000,-413.000000000000,
1515.00000000000,32.0000000000000,
17.0000000000000,-496.000000000000,
22.0000000000000,-458.000000000000,
-185.000000000000,-1287.00000000000,
-536.000000000000,150.000000000000,
587.000000000000,1230.00000000000,
-34.0000000000000,760.000000000000,
1178.00000000000,-35.0000000000000,
288.000000000000,-58.0000000000000,
-583.000000000000,409.000000000000,
119.000000000000,-381.000000000000,
-320.000000000000,985.000000000000,
251.000000000000,-249.000000000000,
399.000000000000,-49.0000000000000,
950.000000000000,225.000000000000,
-757.000000000000,-315.000000000000,
-841.000000000000,583.000000000000,
369.000000000000,-1302.00000000000,
-395.000000000000,51.0000000000000,
71.0000000000000,197.000000000000,
-89.0000000000000,-47.0000000000000,
-555.000000000000,-506.000000000000,
93.0000000000000,-1422.00000000000,
1420.00000000000,196.000000000000,
678.000000000000,748.000000000000,
-175.000000000000,258.000000000000,
538.000000000000,-479.000000000000,
838.000000000000,-19.0000000000000,
93.0000000000000,686.000000000000,
-1412.00000000000,384.000000000000,
-458.000000000000,-271.000000000000,
713.000000000000,-445.000000000000,
566.000000000000,33.0000000000000,
638.000000000000,296.000000000000,
477.000000000000,720.000000000000,
711.000000000000,145.000000000000,
-145.000000000000,-84.0000000000000,
-613.000000000000,-646.000000000000,
360.000000000000,-311.000000000000,
561.000000000000,1552.00000000000,
433.000000000000,215.000000000000,
710.000000000000,-151.000000000000,
296.000000000000,-77.0000000000000,
-715.000000000000,-565.000000000000,
187.000000000000,-496.000000000000,
-53.0000000000000,47.0000000000000,
-385.000000000000,802.000000000000,
605.000000000000,-518.000000000000,
513.000000000000,747.000000000000,
-336.000000000000,659.000000000000,
-109.000000000000,-668.000000000000,
1087.00000000000,953.000000000000,
-578.000000000000,-517.000000000000,
412.000000000000,-649.000000000000,
510.000000000000,1003.00000000000,
-703.000000000000,-340.000000000000,
1219.00000000000,-67.0000000000000,
-686.000000000000,870.000000000000,
-947.000000000000,550.000000000000,
342.000000000000,541.000000000000,
-77.0000000000000,-279.000000000000,
662.000000000000,-213.000000000000,
-144.000000000000,1023.00000000000,
-1338.00000000000,488.000000000000,
-107.000000000000,-350.000000000000,
648.000000000000,-806.000000000000,
590.000000000000,189.000000000000,
-30.0000000000000,806.000000000000,
-354.000000000000,-1079.00000000000,
-5.00000000000000,-767.000000000000,
56.0000000000000,8.00000000000000,
452.000000000000,-2.00000000000000,
196.000000000000,548.000000000000,
-153.000000000000,-59.0000000000000,
-156.000000000000,-894.000000000000,
-717.000000000000,41.0000000000000,
-426.000000000000,725.000000000000,
556.000000000000,-149.000000000000,
177.000000000000,-582.000000000000,
-327.000000000000,-525.000000000000,
-244.000000000000,-624.000000000000,
-198.000000000000,-86.0000000000000,
-127.000000000000,383.000000000000,
-179.000000000000,758.000000000000,
27.0000000000000,-283.000000000000,
-21.0000000000000,-471.000000000000,
635.000000000000,859.000000000000,
224.000000000000,968.000000000000,
-640.000000000000,522.000000000000,
-1072.00000000000,53.0000000000000,
375.000000000000,254.000000000000,
508.000000000000,-236.000000000000,
-1074.00000000000,-555.000000000000,
-452.000000000000,163.000000000000,
-756.000000000000,-15.0000000000000,
369.000000000000,-122.000000000000,
-179.000000000000,-870.000000000000,
-8.00000000000000,-992.000000000000,
650.000000000000,-898.000000000000,
-248.000000000000,-1012.00000000000,
1100.00000000000,710.000000000000,
-187.000000000000,878.000000000000,
-67.0000000000000,418.000000000000,
248.000000000000,388.000000000000,
-372.000000000000,-834.000000000000,
472.000000000000,-1119.00000000000,
561.000000000000,410.000000000000,
787.000000000000,290.000000000000,
807.000000000000,-126.000000000000,
923.000000000000,443.000000000000,
-132.000000000000,-192.000000000000,
-590.000000000000,-258.000000000000,
340.000000000000,266.000000000000,
-468.000000000000,718.000000000000,
-382.000000000000,-723.000000000000,
711.000000000000,-824.000000000000,
39.0000000000000,-36.0000000000000,
628.000000000000,-680.000000000000,
665.000000000000,7.00000000000000,
-789.000000000000,223.000000000000,
-522.000000000000,410.000000000000,
-750.000000000000,384.000000000000,
-1024.00000000000,-752.000000000000,
656.000000000000,-1051.00000000000,
104.000000000000,-516.000000000000,
660.000000000000,6.00000000000000,
1645.00000000000,-133.000000000000,
-396.000000000000,634.000000000000,
-1072.00000000000,493.000000000000,
-702.000000000000,-638.000000000000,
363.000000000000,-21.0000000000000,
585.000000000000,589.000000000000,
-52.0000000000000,-116.000000000000,
197.000000000000,-905.000000000000,
-440.000000000000,-713.000000000000,
347.000000000000,-1342.00000000000,
915.000000000000,-191.000000000000,
-273.000000000000,-15.0000000000000,
696.000000000000,-555.000000000000,
797.000000000000,490.000000000000,
154.000000000000,428.000000000000,
-101.000000000000,1082.00000000000,
-489.000000000000,-263.000000000000,
85.0000000000000,30.0000000000000,
-45.0000000000000,470.000000000000,
-879.000000000000,-693.000000000000,
27.0000000000000,-456.000000000000,
1276.00000000000,-639.000000000000,
264.000000000000,1232.00000000000,
489.000000000000,336.000000000000,
814.000000000000,-362.000000000000,
608.000000000000,-9.00000000000000,
-214.000000000000,-1103.00000000000,
-15.0000000000000,-79.0000000000000,
240.000000000000,666.000000000000,
-149.000000000000,966.000000000000,
490.000000000000,603.000000000000,
-473.000000000000,1202.00000000000,
-973.000000000000,315.000000000000,
-521.000000000000,28.0000000000000,
-335.000000000000,818.000000000000,
367.000000000000,-676.000000000000,
326.000000000000,-17.0000000000000,
837.000000000000,647.000000000000,
-74.0000000000000,702.000000000000,
-719.000000000000,-609.000000000000,
775.000000000000,-403.000000000000,
661.000000000000,1281.00000000000,
-35.0000000000000,303.000000000000,
-422.000000000000,302.000000000000,
-876.000000000000,-43.0000000000000,
-538.000000000000,789.000000000000,
-303.000000000000,198.000000000000,
-144.000000000000,-1084.00000000000,
1342.00000000000,259.000000000000,
5.00000000000000,675.000000000000,
-382.000000000000,1028.00000000000,
363.000000000000,-481.000000000000,
-757.000000000000,-1003.00000000000,
1025.00000000000,-78.0000000000000,
636.000000000000,267.000000000000,
400.000000000000,406.000000000000,
274.000000000000,-282.000000000000,
-989.000000000000,-191.000000000000,
-201.000000000000,-522.000000000000,
296.000000000000,-35.0000000000000,
139.000000000000,-127.000000000000,
109.000000000000,-735.000000000000,
848.000000000000,78.0000000000000,
-282.000000000000,-182.000000000000,
-1140.00000000000,40.0000000000000,
5.00000000000000,520.000000000000,
-298.000000000000,-344.000000000000,
-622.000000000000,49.0000000000000,
423.000000000000,759.000000000000,
649.000000000000,242.000000000000,
105.000000000000,480.000000000000,
1003.00000000000,639.000000000000,
188.000000000000,304.000000000000,
-597.000000000000,990.000000000000,
-42.0000000000000,-737.000000000000,
-1119.00000000000,-96.0000000000000,
457.000000000000,868.000000000000,
-222.000000000000,-741.000000000000,
-1362.00000000000,282.000000000000,
-76.0000000000000,-83.0000000000000,
-833.000000000000,638.000000000000,
36.0000000000000,-347.000000000000,
84.0000000000000,-278.000000000000,
-267.000000000000,695.000000000000,
-185.000000000000,-1278.00000000000,
423.000000000000,165.000000000000,
1407.00000000000,350.000000000000,
256.000000000000,-220.000000000000,
-445.000000000000,-214.000000000000,
-217.000000000000,322.000000000000,
-180.000000000000,829.000000000000,
-812.000000000000,-60.0000000000000,
-82.0000000000000,-769.000000000000,
629.000000000000,-1077.00000000000,
562.000000000000,-142.000000000000,
1189.00000000000,-434.000000000000,
363.000000000000,-295.000000000000,
-309.000000000000,-201.000000000000,
-549.000000000000,-445.000000000000,
-136.000000000000,-994.000000000000,
135.000000000000,-1045.00000000000,
-482.000000000000,978.000000000000,
525.000000000000,-150.000000000000,
335.000000000000,860.000000000000,
-579.000000000000,4.00000000000000,
-668.000000000000,-1469.00000000000,
-323.000000000000,625.000000000000,
-331.000000000000,-1197.00000000000,
-141.000000000000,-510.000000000000,
1117.00000000000,252.000000000000,
43.0000000000000,1027.00000000000,
-20.0000000000000,387.000000000000,
570.000000000000,-663.000000000000,
33.0000000000000,537.000000000000,
165.000000000000,-269.000000000000,
-65.0000000000000,859.000000000000,
451.000000000000,531.000000000000,
11.0000000000000,-641.000000000000,
-661.000000000000,9.00000000000000,
24.0000000000000,171.000000000000,
-576.000000000000,113.000000000000,
-290.000000000000,449.000000000000,
197.000000000000,-343.000000000000,
-213.000000000000,-353.000000000000,
-248.000000000000,422.000000000000,
-695.000000000000,-476.000000000000,
172.000000000000,409.000000000000,
-40.0000000000000,-169.000000000000,
187.000000000000,-1127.00000000000,
952.000000000000,108.000000000000,
554.000000000000,16.0000000000000,
257.000000000000,-537.000000000000,
-610.000000000000,-70.0000000000000,
-92.0000000000000,-149.000000000000,
924.000000000000,37.0000000000000,
960.000000000000,128.000000000000,
83.0000000000000,-451.000000000000,
-764.000000000000,160.000000000000,
-93.0000000000000,70.0000000000000,
-38.0000000000000,-695.000000000000,
-1267.00000000000,203.000000000000,
316.000000000000,315.000000000000,
362.000000000000,-378.000000000000,
-420.000000000000,464.000000000000,
-165.000000000000,-857.000000000000,
-18.0000000000000,-200.000000000000,
729.000000000000,827.000000000000,
-1294.00000000000,-67.0000000000000,
-524.000000000000,-238.000000000000,
502.000000000000,55.0000000000000,
85.0000000000000,1267.00000000000,
-150.000000000000,-856.000000000000,
213.000000000000,-1124.00000000000,
1115.00000000000,153.000000000000,
-407.000000000000,-118.000000000000,
326.000000000000,376.000000000000,
110.000000000000,587.000000000000,
-590.000000000000,1267.00000000000,
-1120.00000000000,334.000000000000,
-902.000000000000,183.000000000000,
750.000000000000,740.000000000000,
-634.000000000000,-616.000000000000,
-691.000000000000,-269.000000000000,
275.000000000000,472.000000000000,
229.000000000000,104.000000000000,
-800.000000000000,202.000000000000,
-1165.00000000000,-2.00000000000000,
817.000000000000,-512.000000000000,
1092.00000000000,-363.000000000000,
15.0000000000000,-252.000000000000,
278.000000000000,374.000000000000,
172.000000000000,-300.000000000000,
177.000000000000,-709.000000000000,
-239.000000000000,672.000000000000,
-567.000000000000,-372.000000000000,
1031.00000000000,-548.000000000000,
947.000000000000,598.000000000000,
26.0000000000000,560.000000000000,
-341.000000000000,321.000000000000,
-613.000000000000,-782.000000000000,
157.000000000000,-951.000000000000,
853.000000000000,-383.000000000000,
678.000000000000,-461.000000000000,
686.000000000000,-122.000000000000,
574.000000000000,30.0000000000000,
423.000000000000,-215.000000000000,
-106.000000000000,350.000000000000,
-6.00000000000000,1065.00000000000,
387.000000000000,-502.000000000000,
-703.000000000000,-199.000000000000,
-98.0000000000000,-119.000000000000,
-553.000000000000,-175.000000000000,
-405.000000000000,-301.000000000000,
507.000000000000,-1210.00000000000,
-82.0000000000000,1247.00000000000,
216.000000000000,-799.000000000000,
-836.000000000000,-291.000000000000,
142.000000000000,473.000000000000,
580.000000000000,-163.000000000000,
-204.000000000000,428.000000000000,
-44.0000000000000,-1735.00000000000,
1003.00000000000,-70.0000000000000,
1340.00000000000,-468.000000000000,
-856.000000000000,548.000000000000,
23.0000000000000,461.000000000000,
214.000000000000,-666.000000000000,
-795.000000000000,1391.00000000000,
-50.0000000000000,311.000000000000,
8.00000000000000,-322.000000000000,
648.000000000000,-14.0000000000000,
478.000000000000,6.00000000000000,
-268.000000000000,-962.000000000000,
736.000000000000,-448.000000000000,
1422.00000000000,312.000000000000,
-997.000000000000,83.0000000000000,
-562.000000000000,539.000000000000,
494.000000000000,-643.000000000000,
-176.000000000000,828.000000000000,
223.000000000000,1491.00000000000,
-1492.00000000000,-212.000000000000,
-242.000000000000,-687.000000000000,
914.000000000000,-954.000000000000,
319.000000000000,1113.00000000000,
149.000000000000,1205.00000000000,
-220.000000000000,-184.000000000000,
-486.000000000000,-29.0000000000000,
-1358.00000000000,418.000000000000,
-186.000000000000,361.000000000000,
-871.000000000000,162.000000000000,
-1343.00000000000,213.000000000000,
204.000000000000,-429.000000000000,
51.0000000000000,-246.000000000000,
574.000000000000,-432.000000000000,
394.000000000000,826.000000000000,
-578.000000000000,672.000000000000,
-1044.00000000000,-816.000000000000,
-463.000000000000,-301.000000000000,
-186.000000000000,-1113.00000000000,
-1223.00000000000,9.00000000000000,
-742.000000000000,161.000000000000,
593.000000000000,-946.000000000000,
307.000000000000,157.000000000000,
-526.000000000000,99.0000000000000,
1163.00000000000,36.0000000000000,
-138.000000000000,127.000000000000,
-716.000000000000,-109.000000000000,
1099.00000000000,-476.000000000000,
-495.000000000000,366.000000000000,
71.0000000000000,117.000000000000,
-396.000000000000,-965.000000000000,
-482.000000000000,-35.0000000000000,
80.0000000000000,-618.000000000000,
-508.000000000000,-674.000000000000,
314.000000000000,-153.000000000000,
318.000000000000,-709.000000000000,
230.000000000000,-10.0000000000000,
271.000000000000,911.000000000000,
652.000000000000,515.000000000000,
-116.000000000000,741.000000000000,
-228.000000000000,1167.00000000000,
894.000000000000,-572.000000000000,
178.000000000000,176.000000000000,
68.0000000000000,638.000000000000,
346.000000000000,245.000000000000,
-765.000000000000,1357.00000000000,
-893.000000000000,125.000000000000,
-550.000000000000,-1025.00000000000,
188.000000000000,-758.000000000000,
463.000000000000,-153.000000000000,
-132.000000000000,-531.000000000000,
-23.0000000000000,-1369.00000000000,
76.0000000000000,-625.000000000000,
-321.000000000000,297.000000000000,
-893.000000000000,219.000000000000,
-682.000000000000,168.000000000000,
698.000000000000,118.000000000000,
-262.000000000000,287.000000000000,
-1305.00000000000,119.000000000000,
-21.0000000000000,-116.000000000000,
-848.000000000000,-407.000000000000,
-34.0000000000000,-539.000000000000,
576.000000000000,471.000000000000,
-310.000000000000,739.000000000000,
16.0000000000000,323.000000000000,
-1139.00000000000,-363.000000000000,
721.000000000000,-641.000000000000,
589.000000000000,-446.000000000000,
-1041.00000000000,444.000000000000,
-200.000000000000,244.000000000000,
-537.000000000000,-379.000000000000,
699.000000000000,-328.000000000000,
609.000000000000,616.000000000000,
-210.000000000000,1090.00000000000,
-78.0000000000000,430.000000000000,
-337.000000000000,1269.00000000000,
-850.000000000000,95.0000000000000,
-1302.00000000000,15.0000000000000,
-106.000000000000,-345.000000000000,
643.000000000000,-567.000000000000,
985.000000000000,282.000000000000,
302.000000000000,149.000000000000,
-870.000000000000,543.000000000000,
-885.000000000000,-805.000000000000,
-470.000000000000,-961.000000000000,
1416.00000000000,-697.000000000000,
1026.00000000000,170.000000000000,
13.0000000000000,-259.000000000000,
1003.00000000000,-421.000000000000,
132.000000000000,808.000000000000,
-200.000000000000,-876.000000000000,
737.000000000000,-155.000000000000,
540.000000000000,1115.00000000000,
117.000000000000,541.000000000000,
-319.000000000000,-127.000000000000,
411.000000000000,-337.000000000000,
1216.00000000000,172.000000000000,
730.000000000000,397.000000000000,
-101.000000000000,-60.0000000000000,
-568.000000000000,-568.000000000000,
-659.000000000000,-317.000000000000,
-526.000000000000,-578.000000000000,
-316.000000000000,-1072.00000000000,
538.000000000000,-1045.00000000000,
1026.00000000000,-446.000000000000,
-507.000000000000,200.000000000000,
-606.000000000000,605.000000000000,
640.000000000000,92.0000000000000,
-48.0000000000000,-230.000000000000,
146.000000000000,130.000000000000,
740.000000000000,40.0000000000000,
302.000000000000,-251.000000000000,
964.000000000000,-117.000000000000,
-235.000000000000,361.000000000000,
-970.000000000000,-91.0000000000000,
281.000000000000,-594.000000000000,
-788.000000000000,-583.000000000000,
43.0000000000000,-153.000000000000,
-57.0000000000000,-969.000000000000,
136.000000000000,-697.000000000000,
824.000000000000,1160.00000000000,
-536.000000000000,48.0000000000000,
-67.0000000000000,-658.000000000000,
-1040.00000000000,-183.000000000000,
670.000000000000,465.000000000000,
582.000000000000,-555.000000000000,
241.000000000000,-483.000000000000,
1060.00000000000,-300.000000000000,
-909.000000000000,-504.000000000000,
591.000000000000,-319.000000000000,
-843.000000000000,126.000000000000,
-835.000000000000,150.000000000000,
731.000000000000,-962.000000000000,
-353.000000000000,737.000000000000,
-202.000000000000,90.0000000000000,
-635.000000000000,224.000000000000,
-262.000000000000,988.000000000000,
229.000000000000,357.000000000000,
569.000000000000,-164.000000000000,
788.000000000000,-836.000000000000,
546.000000000000,223.000000000000,
643.000000000000,-585.000000000000,
286.000000000000,916.000000000000,
978.000000000000,-6.00000000000000,
133.000000000000,5.00000000000000,
-507.000000000000,751.000000000000,
-262.000000000000,-1311.00000000000,
-341.000000000000,-303.000000000000,
1065.00000000000,-833.000000000000,
299.000000000000,1402.00000000000,
-204.000000000000,-125.000000000000,
-316.000000000000,-824.000000000000,
710.000000000000,1259.00000000000,
-267.000000000000,-358.000000000000,
-632.000000000000,1211.00000000000,
551.000000000000,-553.000000000000,
-512.000000000000,-628.000000000000,
531.000000000000,-503.000000000000,
328.000000000000,-361.000000000000,
954.000000000000,981.000000000000,
-341.000000000000,-232.000000000000,
-877.000000000000,1101.00000000000,
-77.0000000000000,265.000000000000,
-1072.00000000000,-111.000000000000,
-450.000000000000,-347.000000000000,
-523.000000000000,-91.0000000000000,
488.000000000000,736.000000000000,
-723.000000000000,583.000000000000,
-305.000000000000,627.000000000000,
363.000000000000,-652.000000000000,
-1020.00000000000,261.000000000000,
166.000000000000,-461.000000000000,
-10.0000000000000,-872.000000000000,
474.000000000000,187.000000000000,
812.000000000000,35.0000000000000,
561.000000000000,-140.000000000000,
712.000000000000,-719.000000000000,
-477.000000000000,357.000000000000,
-65.0000000000000,-530.000000000000,
526.000000000000,-382.000000000000,
213.000000000000,681.000000000000,
345.000000000000,605.000000000000,
-926.000000000000,1016.00000000000,
-912.000000000000,247.000000000000,
165.000000000000,-899.000000000000,
-542.000000000000,-491.000000000000,
359.000000000000,-108.000000000000,
516.000000000000,-308.000000000000,
-823.000000000000,843.000000000000,
345.000000000000,377.000000000000,
134.000000000000,-353.000000000000,
-1028.00000000000,624.000000000000,
756.000000000000,-633.000000000000,
1109.00000000000,-837.000000000000,
-5.00000000000000,283.000000000000,
-682.000000000000,592.000000000000,
-580.000000000000,-601.000000000000,
-371.000000000000,-1236.00000000000,
145.000000000000,1088.00000000000,
886.000000000000,-525.000000000000,
-568.000000000000,58.0000000000000,
-6.00000000000000,-127.000000000000,
-219.000000000000,-1632.00000000000,
16.0000000000000,405.000000000000,
1060.00000000000,-812.000000000000,
958.000000000000,-80.0000000000000,
163.000000000000,64.0000000000000,
-741.000000000000,-534.000000000000,
882.000000000000,-423.000000000000,
821.000000000000,-256.000000000000,
328.000000000000,925.000000000000,
-737.000000000000,-71.0000000000000,
-1151.00000000000,-41.0000000000000,
327.000000000000,558.000000000000,
-486.000000000000,22.0000000000000,
13.0000000000000,-669.000000000000,
646.000000000000,740.000000000000,
-373.000000000000,532.000000000000,
-176.000000000000,243.000000000000,
483.000000000000,1331.00000000000,
379.000000000000,-402.000000000000,
-310.000000000000,-187.000000000000,
-178.000000000000,-799.000000000000,
-309.000000000000,-690.000000000000,
-294.000000000000,783.000000000000,
-569.000000000000,-366.000000000000,
-543.000000000000,595.000000000000,
176.000000000000,-211.000000000000,
262.000000000000,-672.000000000000,
764.000000000000,703.000000000000,
589.000000000000,364.000000000000,
605.000000000000,234.000000000000,
-284.000000000000,750.000000000000,
249.000000000000,164.000000000000,
741.000000000000,83.0000000000000,
-994.000000000000,1164.00000000000,
-470.000000000000,-990.000000000000,
-741.000000000000,-714.000000000000,
-629.000000000000,-20.0000000000000,
487.000000000000,-332.000000000000,
-396.000000000000,1367.00000000000,
-599.000000000000,-19.0000000000000,
297.000000000000,-56.0000000000000,
41.0000000000000,-452.000000000000,
-740.000000000000,-412.000000000000,
-114.000000000000,424.000000000000,
-522.000000000000,-1163.00000000000,
629.000000000000,-537.000000000000,
302.000000000000,-625.000000000000,
-781.000000000000,-359.000000000000,
133.000000000000,822.000000000000,
-168.000000000000,218.000000000000,
180.000000000000,260.000000000000,
-534.000000000000,272.000000000000,
493.000000000000,361.000000000000,
-224.000000000000,817.000000000000,
-1608.00000000000,-305.000000000000,
-103.000000000000,-586.000000000000,
-477.000000000000,942.000000000000,
-39.0000000000000,-232.000000000000,
497.000000000000,-959.000000000000,
158.000000000000,434.000000000000,
699.000000000000,463.000000000000,
-389.000000000000,869.000000000000,
-1143.00000000000,256.000000000000,
-142.000000000000,-280.000000000000,
649.000000000000,-500.000000000000,
473.000000000000,31.0000000000000,
-118.000000000000,422.000000000000,
791.000000000000,-240.000000000000,
-74.0000000000000,822.000000000000,
-1242.00000000000,185.000000000000,
101.000000000000,-499.000000000000,
162.000000000000,-206.000000000000,
297.000000000000,-187.000000000000,
1033.00000000000,259.000000000000,
251.000000000000,-153.000000000000,
398.000000000000,-477.000000000000,
540.000000000000,687.000000000000,
-1055.00000000000,1118.00000000000,
-981.000000000000,-535.000000000000,
-811.000000000000,102.000000000000,
-680.000000000000,-223.000000000000,
-79.0000000000000,-1455.00000000000,
-482.000000000000,32.0000000000000,
398.000000000000,-270.000000000000,
372.000000000000,945.000000000000,
498.000000000000,66.0000000000000,
474.000000000000,-254.000000000000,
-1028.00000000000,851.000000000000,
-1042.00000000000,-1009.00000000000,
-264.000000000000,-17.0000000000000,
1011.00000000000,296.000000000000,
214.000000000000,8.00000000000000,
110.000000000000,-1093.00000000000,
445.000000000000,14.0000000000000,
-502.000000000000,831.000000000000,
459.000000000000,-970.000000000000,
679.000000000000,830.000000000000,
-367.000000000000,1049.00000000000,
662.000000000000,207.000000000000,
354.000000000000,877.000000000000,
-1318.00000000000,674.000000000000,
-577.000000000000,433.000000000000,
-634.000000000000,-272.000000000000,
108.000000000000,-191.000000000000,
432.000000000000,729.000000000000,
-135.000000000000,-308.000000000000,
126.000000000000,99.0000000000000,
-458.000000000000,1010.00000000000,
99.0000000000000,315.000000000000,
-721.000000000000,-25.0000000000000,
-568.000000000000,277.000000000000,
277.000000000000,-356.000000000000,
-713.000000000000,-443.000000000000,
-394.000000000000,-379.000000000000,
-222.000000000000,-426.000000000000,
94.0000000000000,-603.000000000000,
-194.000000000000,-1229.00000000000,
742.000000000000,-783.000000000000,
1015.00000000000,-666.000000000000,
-413.000000000000,403.000000000000,
103.000000000000,-694.000000000000,
-248.000000000000,-41.0000000000000,
-441.000000000000,1085.00000000000,
-825.000000000000,-562.000000000000,
-36.0000000000000,-514.000000000000,
487.000000000000,-1104.00000000000,
179.000000000000,120.000000000000,
763.000000000000,-553.000000000000,
-292.000000000000,-737.000000000000,
876.000000000000,597.000000000000,
672.000000000000,290.000000000000,
-36.0000000000000,509.000000000000,
142.000000000000,-967.000000000000,
-660.000000000000,-30.0000000000000,
-480.000000000000,-246.000000000000,
-514.000000000000,-1349.00000000000,
1142.00000000000,-630.000000000000,
584.000000000000,196.000000000000,
-390.000000000000,842.000000000000,
352.000000000000,-183.000000000000,
337.000000000000,-117.000000000000,
-38.0000000000000,-72.0000000000000,
-83.0000000000000,1035.00000000000,
367.000000000000,581.000000000000,
-413.000000000000,-1498.00000000000,
-121.000000000000,-371.000000000000,
-1111.00000000000,-153.000000000000,
-855.000000000000,316.000000000000,
19.0000000000000,168.000000000000,
-141.000000000000,-809.000000000000,
195.000000000000,272.000000000000,
-1137.00000000000,366.000000000000,
630.000000000000,636.000000000000,
-756.000000000000,448.000000000000,
-1190.00000000000,-79.0000000000000,
222.000000000000,115.000000000000,
-1283.00000000000,240.000000000000,
-197.000000000000,434.000000000000,
-969.000000000000,49.0000000000000,
-691.000000000000,-459.000000000000,
513.000000000000,-1196.00000000000,
-202.000000000000,-949.000000000000,
955.000000000000,-809.000000000000,
473.000000000000,-92.0000000000000,
-447.000000000000,-349.000000000000,
675.000000000000,-38.0000000000000,
601.000000000000,-10.0000000000000,
-532.000000000000,-63.0000000000000,
-175.000000000000,796.000000000000,
470.000000000000,-765.000000000000,
607.000000000000,802.000000000000,
336.000000000000,216.000000000000,
-1374.00000000000,-239.000000000000,
-199.000000000000,377.000000000000,
682.000000000000,-1047.00000000000,
-504.000000000000,715.000000000000,
-506.000000000000,-176.000000000000,
-856.000000000000,-1134.00000000000,
-104.000000000000,-701.000000000000,
-20.0000000000000,-490.000000000000,
229.000000000000,-781.000000000000,
277.000000000000,-1006.00000000000,
-129.000000000000,180.000000000000,
223.000000000000,-1300.00000000000,
124.000000000000,-821.000000000000,
465.000000000000,288.000000000000,
22.0000000000000,15.0000000000000,
473.000000000000,231.000000000000,
-195.000000000000,598.000000000000,
-856.000000000000,666.000000000000,
-402.000000000000,-400.000000000000,
-286.000000000000,166.000000000000,
432.000000000000,-536.000000000000,
295.000000000000,482.000000000000,
193.000000000000,1634.00000000000,
-882.000000000000,-142.000000000000,
-753.000000000000,-570.000000000000,
378.000000000000,-29.0000000000000,
-889.000000000000,610.000000000000,
-245.000000000000,-1120.00000000000,
669.000000000000,264.000000000000,
-308.000000000000,1638.00000000000,
-828.000000000000,-189.000000000000,
-61.0000000000000,-493.000000000000,
50.0000000000000,-1299.00000000000,
769.000000000000,-252.000000000000,
772.000000000000,763.000000000000,
-1033.00000000000,281.000000000000,
-127.000000000000,951.000000000000,
-64.0000000000000,287.000000000000,
-528.000000000000,-257.000000000000,
31.0000000000000,272.000000000000,
424.000000000000,-367.000000000000,
666.000000000000,-453.000000000000,
27.0000000000000,986.000000000000,
-356.000000000000,265.000000000000,
-698.000000000000,-1113.00000000000,
-748.000000000000,-430.000000000000,
-604.000000000000,-103.000000000000,
-495.000000000000,-1021.00000000000,
287.000000000000,-867.000000000000,
-454.000000000000,129.000000000000,
-391.000000000000,-793.000000000000,
1250.00000000000,-773.000000000000,
49.0000000000000,-397.000000000000,
333.000000000000,79.0000000000000,
330.000000000000,413.000000000000,
-257.000000000000,-684.000000000000,
208.000000000000,115.000000000000,
-609.000000000000,-34.0000000000000,
-210.000000000000,677.000000000000,
-49.0000000000000,902.000000000000,
-556.000000000000,-472.000000000000,
347.000000000000,634.000000000000,
578.000000000000,-620.000000000000,
-1062.00000000000,196.000000000000,
183.000000000000,289.000000000000,
240.000000000000,-768.000000000000,
-765.000000000000,476.000000000000,
112.000000000000,625.000000000000,
-747.000000000000,193.000000000000,
-340.000000000000,-760.000000000000,
249.000000000000,-638.000000000000,
530.000000000000,-1120.00000000000,
1124.00000000000,172.000000000000,
571.000000000000,1453.00000000000,
172.000000000000,219.000000000000,
-411.000000000000,27.0000000000000,
-325.000000000000,-694.000000000000,
-25.0000000000000,226.000000000000,
389.000000000000,877.000000000000,
92.0000000000000,284.000000000000,
-421.000000000000,478.000000000000,
-162.000000000000,513.000000000000,
-581.000000000000,-39.0000000000000,
-669.000000000000,-478.000000000000,
614.000000000000,264.000000000000,
423.000000000000,303.000000000000,
-1310.00000000000,419.000000000000,
-433.000000000000,-130.000000000000,
-133.000000000000,-1895.00000000000,
428.000000000000,-574.000000000000,
787.000000000000,136.000000000000,
265.000000000000,-446.000000000000,
1042.00000000000,-519.000000000000,
639.000000000000,-61.0000000000000,
778.000000000000,376.000000000000,
121.000000000000,-521.000000000000,
390.000000000000,-441.000000000000,
940.000000000000,529.000000000000,
-537.000000000000,862.000000000000,
-627.000000000000,-196.000000000000,
-137.000000000000,22.0000000000000,
698.000000000000,49.0000000000000,
-350.000000000000,-795.000000000000,
-627.000000000000,-270.000000000000,
-244.000000000000,-1023.00000000000,
-865.000000000000,45.0000000000000,
134.000000000000,250.000000000000,
788.000000000000,-981.000000000000,
-321.000000000000,13.0000000000000,
-615.000000000000,-612.000000000000,
1298.00000000000,-259.000000000000,
-453.000000000000,441.000000000000,
-345.000000000000,113.000000000000,
637.000000000000,109.000000000000,
-1043.00000000000,-547.000000000000,
1534.00000000000,14.0000000000000,
556.000000000000,1128.00000000000,
-985.000000000000,481.000000000000,
226.000000000000,-355.000000000000,
-371.000000000000,683.000000000000,
13.0000000000000,123.000000000000,
-212.000000000000,54.0000000000000,
-635.000000000000,-83.0000000000000,
-552.000000000000,278.000000000000,
-534.000000000000,-414.000000000000,
78.0000000000000,-1569.00000000000,
-738.000000000000,509.000000000000,
-257.000000000000,-1074.00000000000,
565.000000000000,-569.000000000000,
60.0000000000000,493.000000000000,
218.000000000000,-916.000000000000,
1228.00000000000,208.000000000000,
1109.00000000000,543.000000000000,
-126.000000000000,983.000000000000,
-47.0000000000000,449.000000000000,
41.0000000000000,112.000000000000,
270.000000000000,904.000000000000,
-11.0000000000000,806.000000000000,
-143.000000000000,80.0000000000000,
-333.000000000000,479.000000000000,
443.000000000000,462.000000000000,
756.000000000000,-710.000000000000,
-484.000000000000,826.000000000000,
338.000000000000,-470.000000000000,
-847.000000000000,-517.000000000000,
-954.000000000000,210.000000000000,
285.000000000000,-1795.00000000000,
160.000000000000,1228.00000000000,
130.000000000000,1021.00000000000,
-27.0000000000000,-371.000000000000,
95.0000000000000,636.000000000000,
-553.000000000000,-1021.00000000000,
-59.0000000000000,-677.000000000000,
-474.000000000000,424.000000000000,
583.000000000000,-40.0000000000000,
1237.00000000000,259.000000000000,
-436.000000000000,1645.00000000000,
209.000000000000,-76.0000000000000,
325.000000000000,-932.000000000000,
602.000000000000,338.000000000000,
-728.000000000000,141.000000000000,
-729.000000000000,-84.0000000000000,
351.000000000000,-1215.00000000000,
159.000000000000,-423.000000000000,
596.000000000000,-244.000000000000,
-481.000000000000,-359.000000000000,
1003.00000000000,619.000000000000,
1312.00000000000,31.0000000000000,
-666.000000000000,137.000000000000,
-608.000000000000,315.000000000000,
-788.000000000000,667.000000000000,
-860.000000000000,-832.000000000000,
434.000000000000,-702.000000000000,
1300.00000000000,419.000000000000,
-363.000000000000,-421.000000000000,
-303.000000000000,-473.000000000000,
928.000000000000,-439.000000000000,
47.0000000000000,-592.000000000000,
123.000000000000,-776.000000000000,
488.000000000000,223.000000000000,
248.000000000000,462.000000000000,
-42.0000000000000,-990.000000000000,
-138.000000000000,-514.000000000000,
-241.000000000000,578.000000000000,
-24.0000000000000,1232.00000000000,
-108.000000000000,948.000000000000,
87.0000000000000,385.000000000000,
431.000000000000,1037.00000000000,
-730.000000000000,43.0000000000000,
-233.000000000000,-1474.00000000000,
633.000000000000,-697.000000000000,
346.000000000000,89.0000000000000,
-112.000000000000,-62.0000000000000,
-423.000000000000,177.000000000000,
-6.00000000000000,871.000000000000,
-244.000000000000,709.000000000000,
-77.0000000000000,-68.0000000000000,
39.0000000000000,267.000000000000,
-288.000000000000,676.000000000000,
-587.000000000000,-1082.00000000000,
-802.000000000000,-366.000000000000,
772.000000000000,557.000000000000,
373.000000000000,920.000000000000,
-1088.00000000000,833.000000000000,
-172.000000000000,-218.000000000000,
406.000000000000,688.000000000000,
785.000000000000,101.000000000000,
-709.000000000000,9.00000000000000,
-712.000000000000,-558.000000000000,
256.000000000000,127.000000000000,
-422.000000000000,577.000000000000,
564.000000000000,-984.000000000000,
402.000000000000,184.000000000000,
233.000000000000,-584.000000000000,
486.000000000000,-830.000000000000,
-602.000000000000,435.000000000000,
-288.000000000000,-392.000000000000,
-87.0000000000000,-837.000000000000,
-1249.00000000000,-112.000000000000,
-40.0000000000000,219.000000000000,
-53.0000000000000,-469.000000000000,
-242.000000000000,-718.000000000000,
664.000000000000,317.000000000000,
-824.000000000000,172.000000000000,
268.000000000000,-92.0000000000000,
583.000000000000,562.000000000000,
-342.000000000000,362.000000000000,
117.000000000000,-747.000000000000,
875.000000000000,-410.000000000000,
649.000000000000,1104.00000000000,
-320.000000000000,505.000000000000,
481.000000000000,106.000000000000,
206.000000000000,882.000000000000,
37.0000000000000,1050.00000000000,
45.0000000000000,774.000000000000,
-862.000000000000,382.000000000000,
145.000000000000,-341.000000000000,
-11.0000000000000,207.000000000000,
-1058.00000000000,737.000000000000,
194.000000000000,-352.000000000000,
-89.0000000000000,-100.000000000000,
-898.000000000000,307.000000000000,
60.0000000000000,-479.000000000000,
472.000000000000,-936.000000000000,
547.000000000000,-295.000000000000,
527.000000000000,-191.000000000000,
-610.000000000000,126.000000000000,
99.0000000000000,875.000000000000,
-231.000000000000,-204.000000000000,
-1184.00000000000,512.000000000000,
543.000000000000,-126.000000000000,
269.000000000000,-627.000000000000,
-354.000000000000,369.000000000000,
-1102.00000000000,-494.000000000000,
-104.000000000000,-472.000000000000,
28.0000000000000,-908.000000000000,
-338.000000000000,-464.000000000000,
1218.00000000000,-742.000000000000,
-518.000000000000,-442.000000000000,
362.000000000000,39.0000000000000,
1186.00000000000,-427.000000000000,
-1006.00000000000,665.000000000000,
-167.000000000000,-171.000000000000,
857.000000000000,-340.000000000000,
-368.000000000000,-170.000000000000,
-263.000000000000,-258.000000000000,
590.000000000000,663.000000000000,
-1097.00000000000,566.000000000000,
-1161.00000000000,308.000000000000,
-479.000000000000,-412.000000000000,
267.000000000000,-152.000000000000,
145.000000000000,731.000000000000,
-622.000000000000,366.000000000000,
-420.000000000000,-56.0000000000000,
-1249.00000000000,-516.000000000000,
182.000000000000,-460.000000000000,
269.000000000000,8.00000000000000,
-132.000000000000,583.000000000000,
364.000000000000,-385.000000000000,
-96.0000000000000,-299.000000000000,
610.000000000000,1135.00000000000,
-626.000000000000,847.000000000000,
-877.000000000000,584.000000000000,
-437.000000000000,-508.000000000000,
-213.000000000000,-1212.00000000000,
847.000000000000,-755.000000000000,
740.000000000000,413.000000000000,
1301.00000000000,224.000000000000,
621.000000000000,-122.000000000000,
190.000000000000,-350.000000000000,
-199.000000000000,-1014.00000000000,
-1268.00000000000,275.000000000000,
-529.000000000000,-378.000000000000,
-38.0000000000000,-158.000000000000,
41.0000000000000,-1139.00000000000,
-350.000000000000,-783.000000000000,
377.000000000000,1450.00000000000,
-467.000000000000,200.000000000000,
-1001.00000000000,729.000000000000,
900.000000000000,369.000000000000,
170.000000000000,145.000000000000,
-411.000000000000,746.000000000000,
-346.000000000000,-256.000000000000,
472.000000000000,-1275.00000000000,
724.000000000000,-87.0000000000000,
-200.000000000000,747.000000000000,
-950.000000000000,-1612.00000000000,
-51.0000000000000,-373.000000000000,
835.000000000000,677.000000000000,
-388.000000000000,528.000000000000,
168.000000000000,1234.00000000000,
-1131.00000000000,50.0000000000000,
-1026.00000000000,-39.0000000000000,
653.000000000000,-1115.00000000000,
264.000000000000,-876.000000000000,
1466.00000000000,-424.000000000000,
464.000000000000,-574.000000000000,
370.000000000000,-501.000000000000,
268.000000000000,-178.000000000000,
-18.0000000000000,1396.00000000000,
-25.0000000000000,-881.000000000000,
-745.000000000000,-147.000000000000,
262.000000000000,1128.00000000000,
-411.000000000000,109.000000000000,
-587.000000000000,-249.000000000000,
-435.000000000000,-850.000000000000,
363.000000000000,-916.000000000000,
278.000000000000,-1169.00000000000,
-446.000000000000,512.000000000000,
791.000000000000,-272.000000000000,
407.000000000000,-654.000000000000,
-112.000000000000,141.000000000000,
-1129.00000000000,-476.000000000000,
-83.0000000000000,-69.0000000000000,
1188.00000000000,-16.0000000000000,
227.000000000000,937.000000000000,
489.000000000000,90.0000000000000,
327.000000000000,-293.000000000000,
495.000000000000,-409.000000000000,
176.000000000000,-1085.00000000000,
971.000000000000,370.000000000000,
802.000000000000,416.000000000000,
-513.000000000000,528.000000000000,
-194.000000000000,-463.000000000000,
-651.000000000000,-687.000000000000,
-171.000000000000,1.00000000000000,
-298.000000000000,-399.000000000000,
196.000000000000,-22.0000000000000,
592.000000000000,288.000000000000,
14.0000000000000,298.000000000000,
413.000000000000,-1083.00000000000,
-617.000000000000,172.000000000000,
398.000000000000,-259.000000000000,
671.000000000000,-18.0000000000000,
-93.0000000000000,1352.00000000000,
890.000000000000,-147.000000000000,
-40.0000000000000,494.000000000000,
-528.000000000000,-606.000000000000,
-125.000000000000,-318.000000000000,
-2.00000000000000,49.0000000000000,
-563.000000000000,-814.000000000000,
-287.000000000000,-747.000000000000,
143.000000000000,-57.0000000000000,
-592.000000000000,985.000000000000,
-1088.00000000000,-956.000000000000,
-304.000000000000,250.000000000000,
824.000000000000,258.000000000000,
-681.000000000000,-715.000000000000,
128.000000000000,1514.00000000000,
-447.000000000000,130.000000000000,
0.00000000000000,-34.0000000000000,
1515.00000000000,-98.0000000000000,
-369.000000000000,-497.000000000000,
-219.000000000000,431.000000000000,
152.000000000000,-250.000000000000,
818.000000000000,646.000000000000,
-807.000000000000,419.000000000000,
-34.0000000000000,-300.000000000000,
1341.00000000000,610.000000000000,
-129.000000000000,479.000000000000,
42.0000000000000,184.000000000000,
32.0000000000000,-240.000000000000,
-394.000000000000,-676.000000000000,
-177.000000000000,110.000000000000,
270.000000000000,252.000000000000,
-615.000000000000,91.0000000000000,
-956.000000000000,-76.0000000000000,
521.000000000000,-911.000000000000,
267.000000000000,599.000000000000,
-802.000000000000,377.000000000000,
-304.000000000000,-1370.00000000000,
-192.000000000000,-93.0000000000000,
-810.000000000000,101.000000000000,
-539.000000000000,-28.0000000000000,
282.000000000000,-472.000000000000,
758.000000000000,-534.000000000000,
617.000000000000,1069.00000000000,
-703.000000000000,274.000000000000,
-858.000000000000,-590.000000000000,
-579.000000000000,-305.000000000000,
-415.000000000000,-84.0000000000000,
-130.000000000000,532.000000000000,
194.000000000000,-244.000000000000,
536.000000000000,-649.000000000000,
-470.000000000000,-241.000000000000,
-365.000000000000,-529.000000000000,
-355.000000000000,-362.000000000000,
-369.000000000000,78.0000000000000,
421.000000000000,691.000000000000,
249.000000000000,467.000000000000,
-30.0000000000000,48.0000000000000,
229.000000000000,-452.000000000000,
295.000000000000,-522.000000000000,
171.000000000000,-418.000000000000,
319.000000000000,-965.000000000000,
-653.000000000000,-179.000000000000,
-784.000000000000,804.000000000000,
103.000000000000,998.000000000000,
308.000000000000,627.000000000000,
-130.000000000000,280.000000000000,
-430.000000000000,-312.000000000000,
381.000000000000,-756.000000000000,
301.000000000000,747.000000000000,
-904.000000000000,685.000000000000,
-859.000000000000,270.000000000000,
179.000000000000,417.000000000000,
-221.000000000000,483.000000000000,
-335.000000000000,65.0000000000000,
834.000000000000,-576.000000000000,
-841.000000000000,28.0000000000000,
-508.000000000000,-704.000000000000,
559.000000000000,267.000000000000,
-615.000000000000,709.000000000000,
313.000000000000,34.0000000000000,
271.000000000000,204.000000000000,
829.000000000000,262.000000000000,
379.000000000000,42.0000000000000,
-268.000000000000,-407.000000000000,
827.000000000000,766.000000000000,
-528.000000000000,975.000000000000,
305.000000000000,663.000000000000,
-105.000000000000,-462.000000000000,
-805.000000000000,-846.000000000000,
-62.0000000000000,263.000000000000,
-1075.00000000000,648.000000000000,
-399.000000000000,-719.000000000000,
-188.000000000000,-1112.00000000000,
-172.000000000000,806.000000000000,
-336.000000000000,-364.000000000000,
-337.000000000000,75.0000000000000,
14.0000000000000,720.000000000000,
-430.000000000000,-782.000000000000,
174.000000000000,-424.000000000000,
994.000000000000,-133.000000000000,
86.0000000000000,17.0000000000000,
-1413.00000000000,-363.000000000000,
660.000000000000,-153.000000000000,
549.000000000000,165.000000000000,
-1070.00000000000,-788.000000000000,
-104.000000000000,152.000000000000,
1.00000000000000,567.000000000000,
-650.000000000000,-279.000000000000,
-948.000000000000,376.000000000000,
160.000000000000,110.000000000000,
368.000000000000,-891.000000000000,
32.0000000000000,-146.000000000000,
1369.00000000000,-234.000000000000,
362.000000000000,840.000000000000,
-370.000000000000,644.000000000000,
-310.000000000000,-670.000000000000,
-941.000000000000,257.000000000000,
-114.000000000000,-1290.00000000000,
161.000000000000,-840.000000000000,
332.000000000000,-770.000000000000,
-220.000000000000,-495.000000000000,
-193.000000000000,1331.00000000000,
-892.000000000000,-218.000000000000,
-869.000000000000,-371.000000000000,
241.000000000000,-13.0000000000000,
413.000000000000,139.000000000000,
-35.0000000000000,-122.000000000000,
-458.000000000000,-859.000000000000,
690.000000000000,-1201.00000000000,
80.0000000000000,-631.000000000000,
618.000000000000,712.000000000000,
836.000000000000,364.000000000000,
99.0000000000000,595.000000000000,
-173.000000000000,686.000000000000,
-966.000000000000,8.00000000000000,
505.000000000000,13.0000000000000,
721.000000000000,-80.0000000000000,
287.000000000000,1097.00000000000,
-438.000000000000,88.0000000000000,
23.0000000000000,-532.000000000000,
30.0000000000000,-165.000000000000,
-748.000000000000,-740.000000000000,
572.000000000000,937.000000000000,
204.000000000000,756.000000000000,
621.000000000000,-289.000000000000,
-154.000000000000,215.000000000000,
-580.000000000000,-159.000000000000,
1373.00000000000,-284.000000000000,
-121.000000000000,1140.00000000000,
-340.000000000000,128.000000000000,
798.000000000000,-158.000000000000,
89.0000000000000,392.000000000000,
-757.000000000000,-532.000000000000,
-1032.00000000000,-115.000000000000,
329.000000000000,-978.000000000000,
723.000000000000,-416.000000000000,
-203.000000000000,285.000000000000,
-78.0000000000000,194.000000000000,
-352.000000000000,692.000000000000,
-628.000000000000,-394.000000000000,
707.000000000000,264.000000000000,
206.000000000000,712.000000000000,
-736.000000000000,-445.000000000000,
464.000000000000,-958.000000000000,
40.0000000000000,-817.000000000000,
903.000000000000,-719.000000000000,
173.000000000000,-537.000000000000,
-9.00000000000000,763.000000000000,
805.000000000000,-244.000000000000,
-1134.00000000000,-817.000000000000,
142.000000000000,-527.000000000000,
812.000000000000,143.000000000000,
411.000000000000,603.000000000000,
-282.000000000000,-789.000000000000,
-242.000000000000,231.000000000000,
743.000000000000,-471.000000000000,
247.000000000000,-552.000000000000,
-253.000000000000,-75.0000000000000,
-497.000000000000,-313.000000000000,
-65.0000000000000,1031.00000000000,
-508.000000000000,225.000000000000,
108.000000000000,-522.000000000000,
788.000000000000,-213.000000000000,
-201.000000000000,-954.000000000000,
-93.0000000000000,-82.0000000000000,
-157.000000000000,558.000000000000,
107.000000000000,-704.000000000000,
593.000000000000,411.000000000000,
-423.000000000000,172.000000000000,
306.000000000000,-936.000000000000,
624.000000000000,174.000000000000,
-559.000000000000,-215.000000000000,
-287.000000000000,-97.0000000000000,
-448.000000000000,-623.000000000000,
169.000000000000,-1596.00000000000,
336.000000000000,-223.000000000000,
-631.000000000000,393.000000000000,
36.0000000000000,412.000000000000,
490.000000000000,579.000000000000,
-96.0000000000000,-336.000000000000,
269.000000000000,-620.000000000000,
79.0000000000000,-162.000000000000,
329.000000000000,673.000000000000,
397.000000000000,1585.00000000000,
-1259.00000000000,704.000000000000,
-836.000000000000,-464.000000000000,
458.000000000000,-392.000000000000,
-474.000000000000,-134.000000000000,
-798.000000000000,-96.0000000000000,
113.000000000000,-504.000000000000,
203.000000000000,416.000000000000,
-308.000000000000,1444.00000000000,
-521.000000000000,-466.000000000000,
-549.000000000000,-1141.00000000000,
152.000000000000,-855.000000000000,
-548.000000000000,-752.000000000000,
-341.000000000000,880.000000000000,
471.000000000000,728.000000000000,
-392.000000000000,432.000000000000,
-326.000000000000,-242.000000000000,
-132.000000000000,248.000000000000,
239.000000000000,564.000000000000,
-206.000000000000,-231.000000000000,
709.000000000000,-620.000000000000,
642.000000000000,-162.000000000000,
-717.000000000000,1077.00000000000,
884.000000000000,-451.000000000000,
-105.000000000000,60.0000000000000,
-465.000000000000,-345.000000000000,
-111.000000000000,-699.000000000000,
-366.000000000000,97.0000000000000,
762.000000000000,-728.000000000000,
-612.000000000000,1151.00000000000,
-1439.00000000000,156.000000000000,
-141.000000000000,-986.000000000000,
426.000000000000,11.0000000000000,
51.0000000000000,253.000000000000,
457.000000000000,1021.00000000000,
-392.000000000000,567.000000000000,
-618.000000000000,-147.000000000000,
135.000000000000,-228.000000000000,
-137.000000000000,668.000000000000,
-4.00000000000000,1260.00000000000,
-46.0000000000000,659.000000000000,
371.000000000000,422.000000000000,
9.00000000000000,-218.000000000000,
495.000000000000,-128.000000000000,
409.000000000000,943.000000000000,
-1019.00000000000,376.000000000000,
-1174.00000000000,-128.000000000000,
-231.000000000000,-5.00000000000000,
162.000000000000,475.000000000000,
-873.000000000000,60.0000000000000,
451.000000000000,-187.000000000000,
522.000000000000,1038.00000000000,
-884.000000000000,408.000000000000,
-254.000000000000,-669.000000000000,
-249.000000000000,-30.0000000000000,
-713.000000000000,589.000000000000,
-375.000000000000,409.000000000000,
19.0000000000000,1141.00000000000,
-671.000000000000,269.000000000000,
-439.000000000000,-1492.00000000000,
-171.000000000000,-500.000000000000,
-577.000000000000,355.000000000000,
566.000000000000,-416.000000000000,
-464.000000000000,-279.000000000000,
-265.000000000000,1084.00000000000,
303.000000000000,-327.000000000000,
-286.000000000000,537.000000000000,
566.000000000000,983.000000000000,
-143.000000000000,-20.0000000000000,
968.000000000000,569.000000000000,
-294.000000000000,-125.000000000000,
-295.000000000000,-347.000000000000,
959.000000000000,-755.000000000000,
-398.000000000000,1025.00000000000,
417.000000000000,64.0000000000000,
-571.000000000000,-69.0000000000000,
-1142.00000000000,685.000000000000,
-996.000000000000,-1251.00000000000,
34.0000000000000,-563.000000000000,
909.000000000000,-731.000000000000,
174.000000000000,-332.000000000000,
856.000000000000,-291.000000000000,
634.000000000000,-93.0000000000000,
790.000000000000,349.000000000000,
931.000000000000,59.0000000000000,
307.000000000000,863.000000000000,
-794.000000000000,400.000000000000,
-345.000000000000,-71.0000000000000,
-63.0000000000000,-843.000000000000,
-1136.00000000000,-153.000000000000,
830.000000000000,-150.000000000000,
448.000000000000,305.000000000000,
-297.000000000000,1758.00000000000,
-377.000000000000,685.000000000000,
-1874.00000000000,149.000000000000,
25.0000000000000,-745.000000000000,
130.000000000000,272.000000000000,
158.000000000000,-305.000000000000,
1025.00000000000,-627.000000000000,
218.000000000000,910.000000000000,
492.000000000000,641.000000000000,
-307.000000000000,-28.0000000000000,
-19.0000000000000,-664.000000000000,
292.000000000000,617.000000000000,
-1104.00000000000,-80.0000000000000,
-810.000000000000,10.0000000000000,
202.000000000000,877.000000000000,
858.000000000000,83.0000000000000,
8.00000000000000,132.000000000000,
-1160.00000000000,-279.000000000000,
-734.000000000000,-430.000000000000,
157.000000000000,592.000000000000,
-156.000000000000,290.000000000000,
-638.000000000000,-905.000000000000,
254.000000000000,455.000000000000,
-80.0000000000000,431.000000000000,
215.000000000000,-743.000000000000,
737.000000000000,-230.000000000000,
-307.000000000000,-611.000000000000,
248.000000000000,-123.000000000000,
1275.00000000000,393.000000000000,
-143.000000000000,476.000000000000,
-340.000000000000,1178.00000000000,
122.000000000000,-303.000000000000,
109.000000000000,17.0000000000000,
803.000000000000,812.000000000000,
603.000000000000,-213.000000000000,
919.000000000000,701.000000000000,
94.0000000000000,336.000000000000,
133.000000000000,176.000000000000,
243.000000000000,729.000000000000,
-305.000000000000,-27.0000000000000,
1088.00000000000,-43.0000000000000,
646.000000000000,64.0000000000000,
-803.000000000000,233.000000000000,
-1255.00000000000,-853.000000000000,
-205.000000000000,-452.000000000000,
-871.000000000000,-108.000000000000,
-312.000000000000,-720.000000000000,
991.000000000000,227.000000000000,
-220.000000000000,335.000000000000,
537.000000000000,338.000000000000,
691.000000000000,584.000000000000,
438.000000000000,-160.000000000000,
667.000000000000,-410.000000000000,
364.000000000000,1100.00000000000,
-216.000000000000,994.000000000000,
-1904.00000000000,262.000000000000,
-399.000000000000,-996.000000000000,
251.000000000000,-439.000000000000,
-809.000000000000,511.000000000000,
407.000000000000,-1644.00000000000,
454.000000000000,-181.000000000000,
842.000000000000,109.000000000000,
911.000000000000,-488.000000000000,
297.000000000000,174.000000000000,
-26.0000000000000,-1229.00000000000,
-377.000000000000,-333.000000000000,
96.0000000000000,476.000000000000,
550.000000000000,-333.000000000000,
-55.0000000000000,-608.000000000000,
253.000000000000,-1205.00000000000,
-56.0000000000000,-69.0000000000000,
-590.000000000000,-277.000000000000,
178.000000000000,-1067.00000000000,
98.0000000000000,867.000000000000,
458.000000000000,-269.000000000000,
270.000000000000,-548.000000000000,
16.0000000000000,-360.000000000000,
-18.0000000000000,-459.000000000000,
-192.000000000000,799.000000000000,
-800.000000000000,-181.000000000000,
291.000000000000,-304.000000000000,
695.000000000000,-430.000000000000,
-499.000000000000,-578.000000000000,
398.000000000000,421.000000000000,
354.000000000000,179.000000000000,
-836.000000000000,365.000000000000,
-917.000000000000,-62.0000000000000,
10.0000000000000,-821.000000000000,
40.0000000000000,419.000000000000,
-273.000000000000,893.000000000000,
300.000000000000,695.000000000000,
648.000000000000,-37.0000000000000,
79.0000000000000,-476.000000000000,
970.000000000000,676.000000000000,
-50.0000000000000,-683.000000000000,
-82.0000000000000,-302.000000000000,
398.000000000000,98.0000000000000,
-806.000000000000,-115.000000000000,
105.000000000000,56.0000000000000,
-736.000000000000,-996.000000000000,
802.000000000000,28.0000000000000,
576.000000000000,551.000000000000,
-618.000000000000,492.000000000000,
-181.000000000000,-413.000000000000,
-1191.00000000000,64.0000000000000,
-485.000000000000,-63.0000000000000,
-633.000000000000,-1303.00000000000,
-347.000000000000,118.000000000000,
266.000000000000,-156.000000000000,
501.000000000000,-409.000000000000,
76.0000000000000,280.000000000000,
221.000000000000,367.000000000000,
562.000000000000,398.000000000000,
-609.000000000000,724.000000000000,
204.000000000000,841.000000000000,
505.000000000000,220.000000000000,
-144.000000000000,-384.000000000000,
505.000000000000,-749.000000000000,
454.000000000000,-398.000000000000,
996.000000000000,-536.000000000000,
246.000000000000,1127.00000000000,
35.0000000000000,1245.00000000000,
148.000000000000,136.000000000000,
-789.000000000000,1173.00000000000,
-881.000000000000,-171.000000000000,
-132.000000000000,493.000000000000,
-241.000000000000,340.000000000000,
-1223.00000000000,-247.000000000000,
157.000000000000,798.000000000000,
-54.0000000000000,-834.000000000000,
95.0000000000000,51.0000000000000,
-402.000000000000,383.000000000000,
-1310.00000000000,-145.000000000000,
416.000000000000,-165.000000000000,
236.000000000000,-688.000000000000,
651.000000000000,-702.000000000000,
102.000000000000,-55.0000000000000,
157.000000000000,703.000000000000,
584.000000000000,-147.000000000000,
334.000000000000,476.000000000000,
412.000000000000,-344.000000000000,
-832.000000000000,206.000000000000,
275.000000000000,1283.00000000000,
44.0000000000000,-757.000000000000,
-127.000000000000,-413.000000000000,
-1026.00000000000,-763.000000000000,
-479.000000000000,642.000000000000,
507.000000000000,159.000000000000,
-307.000000000000,-635.000000000000,
1629.00000000000,397.000000000000,
-45.0000000000000,-518.000000000000,
-249.000000000000,1080.00000000000,
-356.000000000000,219.000000000000,
338.000000000000,-85.0000000000000,
1252.00000000000,-153.000000000000,
-334.000000000000,-1093.00000000000,
702.000000000000,483.000000000000,
-454.000000000000,523.000000000000,
222.000000000000,683.000000000000,
-179.000000000000,-273.000000000000,
-481.000000000000,-303.000000000000,
409.000000000000,714.000000000000,
259.000000000000,214.000000000000,
699.000000000000,49.0000000000000,
778.000000000000,-242.000000000000,
749.000000000000,965.000000000000,
-974.000000000000,151.000000000000,
-116.000000000000,-577.000000000000,
130.000000000000,479.000000000000,
-1037.00000000000,-163.000000000000,
590.000000000000,-408.000000000000,
40.0000000000000,600.000000000000,
-428.000000000000,436.000000000000,
-673.000000000000,-171.000000000000,
-1014.00000000000,-86.0000000000000,
-176.000000000000,-786.000000000000,
-205.000000000000,-22.0000000000000,
350.000000000000,-834.000000000000,
-58.0000000000000,-806.000000000000,
169.000000000000,191.000000000000,
1573.00000000000,-439.000000000000,
528.000000000000,528.000000000000,
-323.000000000000,68.0000000000000,
459.000000000000,-121.000000000000,
211.000000000000,596.000000000000,
-1238.00000000000,11.0000000000000,
-248.000000000000,-1209.00000000000,
977.000000000000,-346.000000000000,
-705.000000000000,890.000000000000,
-691.000000000000,63.0000000000000,
159.000000000000,-537.000000000000,
555.000000000000,-1486.00000000000,
209.000000000000,443.000000000000,
366.000000000000,1056.00000000000,
-48.0000000000000,-290.000000000000,
-318.000000000000,62.0000000000000,
912.000000000000,-351.000000000000,
-169.000000000000,1449.00000000000,
-238.000000000000,1254.00000000000,
-1.00000000000000,59.0000000000000,
330.000000000000,-883.000000000000,
210.000000000000,-436.000000000000,
141.000000000000,1099.00000000000,
252.000000000000,-578.000000000000,
-841.000000000000,168.000000000000,
725.000000000000,-485.000000000000,
204.000000000000,353.000000000000,
-177.000000000000,1221.00000000000,
294.000000000000,-1204.00000000000,
-291.000000000000,-383.000000000000,
-943.000000000000,-270.000000000000,
-172.000000000000,-353.000000000000,
1033.00000000000,-658.000000000000,
-121.000000000000,-337.000000000000,
233.000000000000,926.000000000000,
265.000000000000,-230.000000000000,
526.000000000000,20.0000000000000,
274.000000000000,854.000000000000,
-727.000000000000,98.0000000000000,
573.000000000000,-428.000000000000,
603.000000000000,207.000000000000,
209.000000000000,139.000000000000,
-247.000000000000,1016.00000000000,
-419.000000000000,1262.00000000000,
-817.000000000000,408.000000000000,
-950.000000000000,865.000000000000,
884.000000000000,-603.000000000000,
-823.000000000000,254.000000000000,
-522.000000000000,-599.000000000000,
688.000000000000,-335.000000000000,
-245.000000000000,1785.00000000000,
-257.000000000000,400.000000000000,
-427.000000000000,662.000000000000,
309.000000000000,-1164.00000000000,
-617.000000000000,66.0000000000000,
254.000000000000,443.000000000000,
849.000000000000,-1466.00000000000,
-134.000000000000,-98.0000000000000,
-247.000000000000,547.000000000000,
-226.000000000000,832.000000000000,
965.000000000000,-245.000000000000,
-312.000000000000,608.000000000000,
-888.000000000000,-57.0000000000000,
-169.000000000000,-1060.00000000000,
937.000000000000,222.000000000000,
-274.000000000000,-136.000000000000,
-758.000000000000,62.0000000000000,
376.000000000000,-1133.00000000000,
-886.000000000000,-241.000000000000,
80.0000000000000,-373.000000000000,
744.000000000000,-1128.00000000000,
801.000000000000,485.000000000000,
-50.0000000000000,-32.0000000000000,
-123.000000000000,-55.0000000000000,
933.000000000000,293.000000000000,
-641.000000000000,509.000000000000,
144.000000000000,-207.000000000000,
1108.00000000000,-244.000000000000,
202.000000000000,341.000000000000,
-457.000000000000,-127.000000000000,
-951.000000000000,-443.000000000000,
-523.000000000000,114.000000000000,
-400.000000000000,714.000000000000,
-45.0000000000000,104.000000000000,
416.000000000000,460.000000000000,
-52.0000000000000,-634.000000000000,
-598.000000000000,-583.000000000000,
-345.000000000000,650.000000000000,
-98.0000000000000,-968.000000000000,
71.0000000000000,727.000000000000,
-318.000000000000,723.000000000000,
-1280.00000000000,-406.000000000000,
227.000000000000,1252.00000000000,
-632.000000000000,407.000000000000,
-588.000000000000,982.000000000000,
-97.0000000000000,774.000000000000,
-617.000000000000,191.000000000000,
117.000000000000,270.000000000000,
-394.000000000000,-925.000000000000,
600.000000000000,-391.000000000000,
424.000000000000,-1118.00000000000,
57.0000000000000,-1022.00000000000,
-373.000000000000,206.000000000000,
-476.000000000000,-616.000000000000,
202.000000000000,-1191.00000000000,
59.0000000000000,-129.000000000000,
542.000000000000,902.000000000000,
638.000000000000,418.000000000000,
371.000000000000,424.000000000000,
-954.000000000000,255.000000000000,
-1132.00000000000,-146.000000000000,
-465.000000000000,-679.000000000000,
-1193.00000000000,-410.000000000000,
-645.000000000000,-439.000000000000,
-71.0000000000000,-718.000000000000,
524.000000000000,1040.00000000000,
-616.000000000000,354.000000000000,
-318.000000000000,-331.000000000000,
1476.00000000000,-239.000000000000,
-66.0000000000000,232.000000000000,
-51.0000000000000,602.000000000000,
313.000000000000,-844.000000000000,
-545.000000000000,-605.000000000000,
-442.000000000000,356.000000000000,
-391.000000000000,289.000000000000,
-652.000000000000,-214.000000000000,
-320.000000000000,-730.000000000000,
773.000000000000,-971.000000000000,
596.000000000000,653.000000000000,
184.000000000000,1581.00000000000,
36.0000000000000,-402.000000000000,
-12.0000000000000,-304.000000000000,
-352.000000000000,-618.000000000000,
-73.0000000000000,-510.000000000000,
588.000000000000,655.000000000000,
-1133.00000000000,47.0000000000000,
-632.000000000000,-287.000000000000,
-100.000000000000,-837.000000000000,
61.0000000000000,594.000000000000,
107.000000000000,291.000000000000,
-990.000000000000,-120.000000000000,
-527.000000000000,577.000000000000,
-773.000000000000,-517.000000000000,
831.000000000000,493.000000000000,
-64.0000000000000,-433.000000000000,
-387.000000000000,-438.000000000000,
734.000000000000,644.000000000000,
219.000000000000,315.000000000000,
170.000000000000,-65.0000000000000,
-603.000000000000,-168.000000000000,
166.000000000000,791.000000000000,
-91.0000000000000,-628.000000000000,
196.000000000000,66.0000000000000,
397.000000000000,1148.00000000000,
-15.0000000000000,-232.000000000000,
-481.000000000000,326.000000000000,
148.000000000000,-207.000000000000,
585.000000000000,363.000000000000,
-455.000000000000,832.000000000000,
852.000000000000,-118.000000000000,
689.000000000000,804.000000000000,
-336.000000000000,-186.000000000000,
-154.000000000000,-735.000000000000,
-140.000000000000,-56.0000000000000,
259.000000000000,265.000000000000,
-339.000000000000,1427.00000000000,
-907.000000000000,32.0000000000000,
622.000000000000,-846.000000000000,
367.000000000000,1488.00000000000,
-306.000000000000,742.000000000000,
-36.0000000000000,12.0000000000000,
70.0000000000000,-911.000000000000,
-216.000000000000,-1106.00000000000,
299.000000000000,900.000000000000,
729.000000000000,-644.000000000000,
-189.000000000000,-61.0000000000000,
159.000000000000,-565.000000000000,
213.000000000000,-993.000000000000,
791.000000000000,1063.00000000000,
295.000000000000,401.000000000000,
-136.000000000000,1042.00000000000,
-766.000000000000,619.000000000000,
-754.000000000000,-999.000000000000,
1470.00000000000,-708.000000000000,
112.000000000000,771.000000000000,
68.0000000000000,84.0000000000000,
460.000000000000,331.000000000000,
147.000000000000,1263.00000000000,
334.000000000000,-181.000000000000,
-877.000000000000,368.000000000000,
450.000000000000,-1051.00000000000,
-88.0000000000000,-188.000000000000,
-653.000000000000,572.000000000000,
-385.000000000000,-232.000000000000,
-763.000000000000,562.000000000000,
12.0000000000000,-829.000000000000,
348.000000000000,-340.000000000000,
643.000000000000,-301.000000000000,
-459.000000000000,-93.0000000000000,
682.000000000000,-481.000000000000,
476.000000000000,202.000000000000,
-801.000000000000,516.000000000000,
-377.000000000000,-1661.00000000000,
-241.000000000000,296.000000000000,
371.000000000000,407.000000000000,
99.0000000000000,-565.000000000000,
1074.00000000000,-320.000000000000,
442.000000000000,415.000000000000,
-363.000000000000,1838.00000000000,
-990.000000000000,54.0000000000000,
4.00000000000000,285.000000000000,
1205.00000000000,-87.0000000000000,
-110.000000000000,-726.000000000000,
-63.0000000000000,562.000000000000,
-524.000000000000,-82.0000000000000,
1.00000000000000,-305.000000000000,
-113.000000000000,-1056.00000000000,
332.000000000000,-979.000000000000,
531.000000000000,-507.000000000000,
-391.000000000000,-338.000000000000,
448.000000000000,-152.000000000000,
-86.0000000000000,-349.000000000000,
-175.000000000000,-381.000000000000,
-405.000000000000,-516.000000000000,
165.000000000000,-232.000000000000,
-135.000000000000,-507.000000000000,
-863.000000000000,548.000000000000,
514.000000000000,-78.0000000000000,
-435.000000000000,-1039.00000000000,
-1090.00000000000,135.000000000000,
-8.00000000000000,-396.000000000000,
1067.00000000000,657.000000000000,
-351.000000000000,595.000000000000,
-1170.00000000000,-321.000000000000,
-26.0000000000000,380.000000000000,
-603.000000000000,-154.000000000000,
-552.000000000000,38.0000000000000,
-401.000000000000,-36.0000000000000,
-52.0000000000000,-121.000000000000,
-496.000000000000,-61.0000000000000,
-756.000000000000,-1182.00000000000,
866.000000000000,-1051.00000000000,
901.000000000000,427.000000000000,
480.000000000000,-81.0000000000000,
622.000000000000,-196.000000000000,
542.000000000000,773.000000000000,
177.000000000000,351.000000000000,
-832.000000000000,-212.000000000000,
246.000000000000,-750.000000000000,
53.0000000000000,710.000000000000,
-251.000000000000,23.0000000000000,
553.000000000000,392.000000000000,
-407.000000000000,172.000000000000,
273.000000000000,-1079.00000000000,
-564.000000000000,729.000000000000,
-348.000000000000,-1273.00000000000,
213.000000000000,-183.000000000000,
-146.000000000000,1307.00000000000,
310.000000000000,-950.000000000000,
294.000000000000,-206.000000000000,
86.0000000000000,-778.000000000000,
-473.000000000000,-576.000000000000,
-209.000000000000,288.000000000000,
-587.000000000000,-498.000000000000,
-835.000000000000,-82.0000000000000,
328.000000000000,88.0000000000000,
1043.00000000000,862.000000000000,
-541.000000000000,1058.00000000000,
697.000000000000,238.000000000000,
882.000000000000,290.000000000000,
-817.000000000000,247.000000000000,
310.000000000000,394.000000000000,
-276.000000000000,-1021.00000000000,
-70.0000000000000,-880.000000000000,
183.000000000000,349.000000000000,
447.000000000000,-369.000000000000,
178.000000000000,-915.000000000000,
36.0000000000000,143.000000000000,
1330.00000000000,242.000000000000,
-118.000000000000,177.000000000000,
149.000000000000,1392.00000000000,
686.000000000000,-997.000000000000,
-665.000000000000,-846.000000000000,
-13.0000000000000,796.000000000000,
879.000000000000,-157.000000000000,
182.000000000000,724.000000000000,
-584.000000000000,1.00000000000000,
107.000000000000,-1031.00000000000,
-391.000000000000,-143.000000000000,
508.000000000000,801.000000000000,
-133.000000000000,453.000000000000,
-1708.00000000000,327.000000000000,
564.000000000000,-444.000000000000,
509.000000000000,-124.000000000000,
-270.000000000000,1815.00000000000,
-504.000000000000,48.0000000000000,
316.000000000000,-444.000000000000,
192.000000000000,180.000000000000,
-1089.00000000000,571.000000000000,
311.000000000000,-550.000000000000,
-184.000000000000,-757.000000000000,
202.000000000000,771.000000000000,
-61.0000000000000,92.0000000000000,
-776.000000000000,726.000000000000,
-149.000000000000,640.000000000000,
-1350.00000000000,48.0000000000000,
-118.000000000000,-456.000000000000,
192.000000000000,271.000000000000,
-436.000000000000,341.000000000000,
827.000000000000,-448.000000000000,
666.000000000000,125.000000000000,
132.000000000000,-1188.00000000000,
-307.000000000000,-513.000000000000,
-147.000000000000,142.000000000000,
414.000000000000,15.0000000000000,
597.000000000000,732.000000000000,
-713.000000000000,-336.000000000000,
274.000000000000,-544.000000000000,
1333.00000000000,-175.000000000000,
338.000000000000,-315.000000000000,
521.000000000000,-1010.00000000000,
498.000000000000,-702.000000000000,
-185.000000000000,339.000000000000,
-1042.00000000000,271.000000000000,
-189.000000000000,442.000000000000,
326.000000000000,514.000000000000,
-512.000000000000,260.000000000000,
-41.0000000000000,-991.000000000000,
53.0000000000000,-1320.00000000000,
9.00000000000000,-403.000000000000,
-6.00000000000000,-538.000000000000,
-50.0000000000000,-379.000000000000,
-301.000000000000,-312.000000000000,
-27.0000000000000,-538.000000000000,
-124.000000000000,-868.000000000000,
-583.000000000000,133.000000000000,
1204.00000000000,88.0000000000000,
48.0000000000000,-780.000000000000,
-450.000000000000,941.000000000000,
311.000000000000,1101.00000000000,
-1083.00000000000,261.000000000000,
-208.000000000000,-781.000000000000,
-294.000000000000,181.000000000000,
495.000000000000,603.000000000000,
1090.00000000000,33.0000000000000,
209.000000000000,157.000000000000,
110.000000000000,-293.000000000000,
333.000000000000,1083.00000000000,
403.000000000000,-717.000000000000,
194.000000000000,-809.000000000000,
118.000000000000,1017.00000000000,
-1041.00000000000,-514.000000000000,
437.000000000000,13.0000000000000,
202.000000000000,-13.0000000000000,
37.0000000000000,266.000000000000,
843.000000000000,830.000000000000,
-1297.00000000000,360.000000000000,
-356.000000000000,-371.000000000000,
977.000000000000,-1083.00000000000,
387.000000000000,482.000000000000,
-786.000000000000,456.000000000000,
-543.000000000000,843.000000000000,
-680.000000000000,268.000000000000,
-112.000000000000,-627.000000000000,
857.000000000000,722.000000000000,
155.000000000000,-269.000000000000,
1012.00000000000,155.000000000000,
-523.000000000000,86.0000000000000,
-393.000000000000,61.0000000000000,
-145.000000000000,682.000000000000,
281.000000000000,117.000000000000,
516.000000000000,902.000000000000,
-1376.00000000000,-72.0000000000000,
296.000000000000,-254.000000000000,
-1.00000000000000,614.000000000000,
-727.000000000000,999.000000000000,
-204.000000000000,-615.000000000000,
-286.000000000000,-1397.00000000000,
153.000000000000,154.000000000000,
-281.000000000000,590.000000000000,
456.000000000000,753.000000000000,
-284.000000000000,361.000000000000,
-1005.00000000000,491.000000000000,
71.0000000000000,-233.000000000000,
510.000000000000,-112.000000000000,
603.000000000000,707.000000000000,
103.000000000000,-277.000000000000,
415.000000000000,-662.000000000000,
562.000000000000,-340.000000000000,
655.000000000000,610.000000000000,
-235.000000000000,-756.000000000000,
70.0000000000000,0.00000000000000,
-36.0000000000000,1300.00000000000,
-599.000000000000,-455.000000000000,
1344.00000000000,286.000000000000,
-255.000000000000,381.000000000000,
-1294.00000000000,-166.000000000000,
-180.000000000000,110.000000000000,
-75.0000000000000,-595.000000000000,
247.000000000000,-776.000000000000,
-272.000000000000,-967.000000000000,
-52.0000000000000,-637.000000000000,
242.000000000000,757.000000000000,
-928.000000000000,358.000000000000,
-349.000000000000,-948.000000000000,
1079.00000000000,-48.0000000000000,
-37.0000000000000,649.000000000000,
-542.000000000000,918.000000000000,
504.000000000000,-51.0000000000000,
164.000000000000,-1023.00000000000,
-61.0000000000000,490.000000000000,
-136.000000000000,892.000000000000,
-869.000000000000,-505.000000000000,
743.000000000000,-548.000000000000,
1051.00000000000,202.000000000000,
-759.000000000000,559.000000000000,
300.000000000000,105.000000000000,
416.000000000000,-560.000000000000,
-503.000000000000,579.000000000000,
732.000000000000,862.000000000000,
618.000000000000,130.000000000000,
-61.0000000000000,846.000000000000,
45.0000000000000,263.000000000000,
-650.000000000000,-701.000000000000,
686.000000000000,-556.000000000000,
1084.00000000000,171.000000000000,
-550.000000000000,426.000000000000,
466.000000000000,-693.000000000000,
-243.000000000000,187.000000000000,
-926.000000000000,-183.000000000000,
424.000000000000,-1400.00000000000,
884.000000000000,52.0000000000000,
-155.000000000000,-632.000000000000,
-871.000000000000,122.000000000000,
-658.000000000000,119.000000000000,
-325.000000000000,-584.000000000000,
-42.0000000000000,538.000000000000,
-542.000000000000,-960.000000000000,
145.000000000000,-974.000000000000,
-329.000000000000,314.000000000000,
50.0000000000000,171.000000000000,
710.000000000000,23.0000000000000,
-977.000000000000,287.000000000000,
-938.000000000000,-192.000000000000,
-504.000000000000,-581.000000000000,
598.000000000000,-739.000000000000,
395.000000000000,-627.000000000000,
236.000000000000,715.000000000000,
823.000000000000,-147.000000000000,
-399.000000000000,-3.00000000000000,
295.000000000000,315.000000000000,
-270.000000000000,601.000000000000,
-630.000000000000,-38.0000000000000,
383.000000000000,-1778.00000000000,
140.000000000000,-292.000000000000,
211.000000000000,-502.000000000000,
-244.000000000000,-346.000000000000,
-141.000000000000,54.0000000000000,
-1096.00000000000,-450.000000000000,
-139.000000000000,-830.000000000000,
-173.000000000000,-1025.00000000000,
-930.000000000000,155.000000000000,
514.000000000000,-570.000000000000,
53.0000000000000,676.000000000000,
-168.000000000000,557.000000000000,
-915.000000000000,-626.000000000000,
315.000000000000,-700.000000000000,
67.0000000000000,-973.000000000000,
-194.000000000000,269.000000000000,
640.000000000000,-296.000000000000,
-993.000000000000,115.000000000000,
483.000000000000,-1341.00000000000,
-186.000000000000,100.000000000000,
258.000000000000,901.000000000000,
250.000000000000,-265.000000000000,
-282.000000000000,1741.00000000000,
522.000000000000,-473.000000000000,
-1529.00000000000,-154.000000000000,
-425.000000000000,-274.000000000000,
-457.000000000000,-1321.00000000000,
-11.0000000000000,-635.000000000000,
998.000000000000,-163.000000000000,
-195.000000000000,839.000000000000,
-307.000000000000,-695.000000000000,
-7.00000000000000,-1239.00000000000,
676.000000000000,-654.000000000000,
-207.000000000000,102.000000000000,
329.000000000000,-300.000000000000,
721.000000000000,410.000000000000,
352.000000000000,1065.00000000000,
470.000000000000,315.000000000000,
-895.000000000000,849.000000000000,
-1083.00000000000,-159.000000000000,
447.000000000000,-224.000000000000,
762.000000000000,603.000000000000,
-131.000000000000,594.000000000000,
297.000000000000,568.000000000000,
48.0000000000000,535.000000000000,
-978.000000000000,873.000000000000,
-698.000000000000,332.000000000000,
55.0000000000000,528.000000000000,
-25.0000000000000,351.000000000000,
-1121.00000000000,-473.000000000000,
-113.000000000000,811.000000000000,
670.000000000000,80.0000000000000,
686.000000000000,96.0000000000000,
-212.000000000000,750.000000000000,
-1302.00000000000,55.0000000000000,
-249.000000000000,471.000000000000,
-112.000000000000,-575.000000000000,
553.000000000000,25.0000000000000,
393.000000000000,784.000000000000,
-250.000000000000,-164.000000000000,
-306.000000000000,521.000000000000,
-188.000000000000,632.000000000000,
-59.0000000000000,-1149.00000000000,
-721.000000000000,-389.000000000000,
-260.000000000000,318.000000000000,
-1011.00000000000,-551.000000000000,
-1227.00000000000,-133.000000000000,
779.000000000000,-652.000000000000,
421.000000000000,623.000000000000,
749.000000000000,855.000000000000,
1074.00000000000,-233.000000000000,
306.000000000000,986.000000000000,
442.000000000000,478.000000000000,
97.0000000000000,-486.000000000000,
364.000000000000,464.000000000000,
-158.000000000000,252.000000000000,
-281.000000000000,-754.000000000000,
590.000000000000,592.000000000000,
1017.00000000000,-6.00000000000000,
-251.000000000000,-246.000000000000,
-416.000000000000,1101.00000000000,
551.000000000000,-845.000000000000,
248.000000000000,577.000000000000,
818.000000000000,662.000000000000,
125.000000000000,-281.000000000000,
149.000000000000,1093.00000000000,
-656.000000000000,-337.000000000000,
-300.000000000000,248.000000000000,
686.000000000000,-624.000000000000,
-408.000000000000,-1103.00000000000,
350.000000000000,-190.000000000000,
-315.000000000000,150.000000000000,
-158.000000000000,885.000000000000,
-858.000000000000,-55.0000000000000,
-383.000000000000,155.000000000000,
1240.00000000000,-17.0000000000000,
-414.000000000000,-66.0000000000000,
-329.000000000000,230.000000000000,
265.000000000000,556.000000000000,
-340.000000000000,60.0000000000000,
-323.000000000000,-74.0000000000000,
836.000000000000,778.000000000000,
-238.000000000000,-29.0000000000000,
-572.000000000000,986.000000000000,
1057.00000000000,-40.0000000000000,
-785.000000000000,-273.000000000000,
-64.0000000000000,1138.00000000000,
-222.000000000000,-31.0000000000000,
-1442.00000000000,-24.0000000000000,
-41.0000000000000,-837.000000000000,
652.000000000000,-229.000000000000,
-361.000000000000,397.000000000000,
-1341.00000000000,-203.000000000000,
-201.000000000000,-650.000000000000,
-530.000000000000,-958.000000000000,
-187.000000000000,1.00000000000000,
-500.000000000000,-75.0000000000000,
-1259.00000000000,-637.000000000000,
1224.00000000000,-572.000000000000,
985.000000000000,319.000000000000,
288.000000000000,-842.000000000000,
133.000000000000,-1150.00000000000,
-558.000000000000,500.000000000000,
-115.000000000000,45.0000000000000,
-618.000000000000,-74.0000000000000,
-201.000000000000,227.000000000000,
28.0000000000000,862.000000000000,
-18.0000000000000,475.000000000000,
-427.000000000000,395.000000000000,
-395.000000000000,-636.000000000000,
688.000000000000,-798.000000000000,
500.000000000000,1167.00000000000,
587.000000000000,-264.000000000000,
1013.00000000000,439.000000000000,
-67.0000000000000,1056.00000000000,
-1539.00000000000,-206.000000000000,
45.0000000000000,746.000000000000,
-224.000000000000,-37.0000000000000,
-722.000000000000,469.000000000000,
-202.000000000000,94.0000000000000,
-265.000000000000,-1074.00000000000,
1111.00000000000,-620.000000000000,
-398.000000000000,-751.000000000000,
-111.000000000000,-486.000000000000,
-273.000000000000,-429.000000000000,
-1059.00000000000,-55.0000000000000,
863.000000000000,-521.000000000000,
-478.000000000000,17.0000000000000,
-410.000000000000,-27.0000000000000,
828.000000000000,-617.000000000000,
642.000000000000,-41.0000000000000,
557.000000000000,491.000000000000,
140.000000000000,664.000000000000,
-304.000000000000,-175.000000000000,
-1140.00000000000,198.000000000000,
121.000000000000,-1264.00000000000,
361.000000000000,-1152.00000000000,
683.000000000000,-532.000000000000,
369.000000000000,-510.000000000000,
-482.000000000000,665.000000000000,
908.000000000000,-438.000000000000,
461.000000000000,507.000000000000,
-196.000000000000,84.0000000000000,
-1081.00000000000,-177.000000000000,
-2.00000000000000,-335.000000000000,
253.000000000000,-1302.00000000000,
643.000000000000,419.000000000000,
1036.00000000000,-27.0000000000000,
-825.000000000000,955.000000000000,
720.000000000000,1108.00000000000,
-367.000000000000,658.000000000000,
-913.000000000000,1014.00000000000,
-230.000000000000,-324.000000000000,
-1426.00000000000,242.000000000000,
-768.000000000000,-686.000000000000,
463.000000000000,-385.000000000000,
451.000000000000,613.000000000000,
-283.000000000000,-325.000000000000,
641.000000000000,-1042.00000000000,
212.000000000000,-215.000000000000,
-145.000000000000,878.000000000000,
53.0000000000000,684.000000000000,
-697.000000000000,592.000000000000,
-182.000000000000,501.000000000000,
-229.000000000000,717.000000000000,
949.000000000000,119.000000000000,
374.000000000000,975.000000000000,
-1040.00000000000,117.000000000000,
267.000000000000,-907.000000000000,
-193.000000000000,800.000000000000,
283.000000000000,-517.000000000000,
-77.0000000000000,455.000000000000,
-685.000000000000,420.000000000000,
232.000000000000,-1195.00000000000,
151.000000000000,367.000000000000,
-242.000000000000,-339.000000000000,
-558.000000000000,-810.000000000000,
164.000000000000,287.000000000000,
-310.000000000000,744.000000000000,
-367.000000000000,878.000000000000,
383.000000000000,446.000000000000,
-473.000000000000,-134.000000000000,
-817.000000000000,-423.000000000000,
698.000000000000,-886.000000000000,
93.0000000000000,90.0000000000000,
-1129.00000000000,1104.00000000000,
385.000000000000,-744.000000000000,
-262.000000000000,-551.000000000000,
178.000000000000,736.000000000000,
592.000000000000,429.000000000000,
-819.000000000000,1247.00000000000,
229.000000000000,96.0000000000000,
-284.000000000000,235.000000000000,
-126.000000000000,281.000000000000,
1048.00000000000,-233.000000000000,
479.000000000000,729.000000000000,
-1294.00000000000,-69.0000000000000,
-559.000000000000,-161.000000000000,
314.000000000000,-1067.00000000000,
-1379.00000000000,-10.0000000000000,
938.000000000000,31.0000000000000,
69.0000000000000,-326.000000000000,
257.000000000000,1138.00000000000,
573.000000000000,-471.000000000000,
-1706.00000000000,16.0000000000000,
360.000000000000,-543.000000000000,
964.000000000000,-433.000000000000,
-738.000000000000,-273.000000000000,
-781.000000000000,-588.000000000000,
513.000000000000,649.000000000000,
-890.000000000000,-39.0000000000000,
644.000000000000,123.000000000000,
1564.00000000000,72.0000000000000,
-625.000000000000,1149.00000000000,
-7.00000000000000,530.000000000000,
-893.000000000000,-259.000000000000,
-1001.00000000000,651.000000000000,
-1260.00000000000,-1209.00000000000,
265.000000000000,232.000000000000,
303.000000000000,9.00000000000000,
-1477.00000000000,-367.000000000000,
-250.000000000000,7.00000000000000,
-1176.00000000000,-1035.00000000000,
-17.0000000000000,53.0000000000000,
421.000000000000,-236.000000000000,
-387.000000000000,224.000000000000,
-398.000000000000,-538.000000000000,
422.000000000000,-690.000000000000,
1194.00000000000,-200.000000000000,
-932.000000000000,12.0000000000000,
29.0000000000000,319.000000000000,
333.000000000000,599.000000000000,
-1146.00000000000,718.000000000000,
-701.000000000000,17.0000000000000,
-936.000000000000,560.000000000000,
-888.000000000000,-532.000000000000,
-966.000000000000,-808.000000000000,
-209.000000000000,-568.000000000000,
528.000000000000,-500.000000000000,
532.000000000000,1043.00000000000,
-45.0000000000000,519.000000000000,
-719.000000000000,-22.0000000000000,
-516.000000000000,-530.000000000000,
-483.000000000000,-876.000000000000,
830.000000000000,-1394.00000000000,
349.000000000000,-234.000000000000,
-410.000000000000,851.000000000000,
16.0000000000000,-1359.00000000000,
428.000000000000,-125.000000000000,
810.000000000000,693.000000000000,
-727.000000000000,-243.000000000000,
739.000000000000,-178.000000000000,
188.000000000000,702.000000000000,
-529.000000000000,481.000000000000,
770.000000000000,89.0000000000000,
-1180.00000000000,651.000000000000,
-499.000000000000,-690.000000000000,
81.0000000000000,1173.00000000000,
-60.0000000000000,815.000000000000,
127.000000000000,-1076.00000000000,
761.000000000000,230.000000000000,
502.000000000000,436.000000000000,
-1044.00000000000,492.000000000000,
-664.000000000000,3.00000000000000,
-259.000000000000,1150.00000000000,
243.000000000000,136.000000000000,
130.000000000000,-1457.00000000000,
1004.00000000000,-64.0000000000000,
1020.00000000000,-311.000000000000,
404.000000000000,-341.000000000000,
1146.00000000000,258.000000000000,
-105.000000000000,816.000000000000,
254.000000000000,118.000000000000,
337.000000000000,141.000000000000,
-498.000000000000,1205.00000000000,
-677.000000000000,-471.000000000000,
213.000000000000,-1331.00000000000,
1437.00000000000,-375.000000000000,
605.000000000000,595.000000000000,
239.000000000000,343.000000000000,
365.000000000000,138.000000000000,
861.000000000000,176.000000000000,
489.000000000000,378.000000000000,
-149.000000000000,795.000000000000,
-956.000000000000,-605.000000000000,
-1032.00000000000,295.000000000000,
304.000000000000,-423.000000000000,
-586.000000000000,-1041.00000000000,
-268.000000000000,1026.00000000000,
102.000000000000,-676.000000000000,
672.000000000000,129.000000000000,
-22.0000000000000,813.000000000000,
-1206.00000000000,-292.000000000000,
838.000000000000,0.00000000000000,
-467.000000000000,-52.0000000000000,
-270.000000000000,-469.000000000000,
199.000000000000,-914.000000000000,
-728.000000000000,322.000000000000,
-22.0000000000000,222.000000000000,
218.000000000000,796.000000000000,
-130.000000000000,-180.000000000000,
377.000000000000,-935.000000000000,
841.000000000000,591.000000000000,
-978.000000000000,-458.000000000000,
-330.000000000000,79.0000000000000,
115.000000000000,-244.000000000000,
-196.000000000000,-548.000000000000,
471.000000000000,777.000000000000,
694.000000000000,127.000000000000,
-171.000000000000,705.000000000000,
-739.000000000000,-356.000000000000,
826.000000000000,-401.000000000000,
-118.000000000000,1532.00000000000,
12.0000000000000,-519.000000000000,
829.000000000000,-1404.00000000000,
-601.000000000000,556.000000000000,
39.0000000000000,-606.000000000000,
182.000000000000,-599.000000000000,
175.000000000000,958.000000000000,
371.000000000000,-440.000000000000,
-732.000000000000,-184.000000000000,
915.000000000000,-228.000000000000,
210.000000000000,899.000000000000,
-465.000000000000,1251.00000000000,
-435.000000000000,242.000000000000,
-276.000000000000,-336.000000000000,
260.000000000000,-1357.00000000000,
-457.000000000000,486.000000000000,
479.000000000000,160.000000000000,
-441.000000000000,234.000000000000,
127.000000000000,-43.0000000000000,
415.000000000000,-542.000000000000,
-1368.00000000000,698.000000000000,
-632.000000000000,-783.000000000000,
607.000000000000,-87.0000000000000,
-633.000000000000,194.000000000000,
-420.000000000000,-765.000000000000,
976.000000000000,775.000000000000,
-550.000000000000,281.000000000000,
-129.000000000000,-809.000000000000,
563.000000000000,-1048.00000000000,
483.000000000000,-696.000000000000,
869.000000000000,432.000000000000,
71.0000000000000,225.000000000000,
-260.000000000000,-328.000000000000,
90.0000000000000,248.000000000000,
495.000000000000,142.000000000000,
-285.000000000000,246.000000000000,
-341.000000000000,382.000000000000,
569.000000000000,-853.000000000000,
-566.000000000000,9.00000000000000,
-656.000000000000,-35.0000000000000,
-282.000000000000,43.0000000000000,
-685.000000000000,299.000000000000,
-303.000000000000,-1315.00000000000,
900.000000000000,-657.000000000000,
748.000000000000,-1067.00000000000,
747.000000000000,-622.000000000000,
1690.00000000000,653.000000000000,
40.0000000000000,-546.000000000000,
-355.000000000000,442.000000000000,
5.00000000000000,861.000000000000,
-189.000000000000,345.000000000000,
-3.00000000000000,260.000000000000,
-72.0000000000000,-677.000000000000,
771.000000000000,-759.000000000000,
755.000000000000,782.000000000000,
196.000000000000,599.000000000000,
-585.000000000000,-481.000000000000,
-241.000000000000,-314.000000000000,
410.000000000000,-160.000000000000,
445.000000000000,796.000000000000,
589.000000000000,-340.000000000000,
-608.000000000000,-558.000000000000,
95.0000000000000,1201.00000000000,
567.000000000000,486.000000000000,
-732.000000000000,373.000000000000,
-123.000000000000,440.000000000000,
-121.000000000000,-356.000000000000,
-664.000000000000,-63.0000000000000,
144.000000000000,-234.000000000000,
-394.000000000000,-676.000000000000,
-768.000000000000,191.000000000000,
-205.000000000000,318.000000000000,
-1063.00000000000,-417.000000000000,
-95.0000000000000,-417.000000000000,
895.000000000000,418.000000000000,
418.000000000000,586.000000000000,
487.000000000000,-783.000000000000,
308.000000000000,-1259.00000000000,
869.000000000000,241.000000000000,
948.000000000000,-125.000000000000,
-191.000000000000,-802.000000000000,
-270.000000000000,131.000000000000,
39.0000000000000,-9.00000000000000,
400.000000000000,-478.000000000000,
585.000000000000,-989.000000000000,
256.000000000000,-771.000000000000,
265.000000000000,117.000000000000,
28.0000000000000,272.000000000000,
-660.000000000000,-375.000000000000,
569.000000000000,92.0000000000000,
1194.00000000000,329.000000000000,
-60.0000000000000,-590.000000000000,
1356.00000000000,161.000000000000,
881.000000000000,395.000000000000,
-619.000000000000,171.000000000000,
59.0000000000000,-1240.00000000000,
-106.000000000000,-288.000000000000,
-493.000000000000,1496.00000000000,
-638.000000000000,-1181.00000000000,
408.000000000000,-229.000000000000,
-586.000000000000,546.000000000000,
-678.000000000000,-594.000000000000,
414.000000000000,-854.000000000000,
567.000000000000,-165.000000000000,
1017.00000000000,957.000000000000,
-992.000000000000,600.000000000000,
-375.000000000000,-288.000000000000,
205.000000000000,-1337.00000000000,
-377.000000000000,712.000000000000,
142.000000000000,381.000000000000,
-927.000000000000,18.0000000000000,
-40.0000000000000,455.000000000000,
-1100.00000000000,-520.000000000000,
-832.000000000000,126.000000000000,
222.000000000000,-474.000000000000,
-446.000000000000,-416.000000000000,
330.000000000000,-818.000000000000,
-429.000000000000,299.000000000000,
-374.000000000000,813.000000000000,
-533.000000000000,706.000000000000,
212.000000000000,186.000000000000,
613.000000000000,-1105.00000000000,
1096.00000000000,312.000000000000,
1182.00000000000,81.0000000000000,
-860.000000000000,1190.00000000000,
472.000000000000,180.000000000000,
60.0000000000000,-727.000000000000,
-56.0000000000000,860.000000000000,
120.000000000000,581.000000000000,
-90.0000000000000,965.000000000000,
1019.00000000000,260.000000000000,
-567.000000000000,-288.000000000000,
220.000000000000,-676.000000000000,
281.000000000000,555.000000000000,
-587.000000000000,1141.00000000000,
17.0000000000000,-95.0000000000000,
363.000000000000,-305.000000000000,
535.000000000000,-1141.00000000000,
-295.000000000000,-420.000000000000,
158.000000000000,29.0000000000000,
364.000000000000,506.000000000000,
-313.000000000000,1251.00000000000,
-283.000000000000,75.0000000000000,
592.000000000000,-378.000000000000,
750.000000000000,25.0000000000000,
635.000000000000,1193.00000000000,
-234.000000000000,805.000000000000,
-166.000000000000,-1053.00000000000,
552.000000000000,-218.000000000000,
-278.000000000000,453.000000000000,
255.000000000000,206.000000000000,
-234.000000000000,-600.000000000000,
408.000000000000,-447.000000000000,
531.000000000000,705.000000000000,
-944.000000000000,205.000000000000,
424.000000000000,180.000000000000,
-37.0000000000000,636.000000000000,
-577.000000000000,-49.0000000000000,
562.000000000000,-919.000000000000,
-142.000000000000,-324.000000000000,
-389.000000000000,-106.000000000000,
18.0000000000000,-740.000000000000,
884.000000000000,-928.000000000000,
401.000000000000,611.000000000000,
-534.000000000000,203.000000000000,
267.000000000000,-1873.00000000000,
934.000000000000,73.0000000000000,
877.000000000000,-65.0000000000000,
245.000000000000,-305.000000000000,
688.000000000000,1226.00000000000,
-531.000000000000,270.000000000000,
-1249.00000000000,205.000000000000,
-394.000000000000,-369.000000000000,
57.0000000000000,-137.000000000000,
-182.000000000000,-154.000000000000,
-263.000000000000,-1081.00000000000,
688.000000000000,-916.000000000000,
343.000000000000,187.000000000000,
602.000000000000,896.000000000000,
-554.000000000000,-286.000000000000,
-1480.00000000000,-402.000000000000,
607.000000000000,251.000000000000,
-75.0000000000000,300.000000000000,
-826.000000000000,-77.0000000000000,
-45.0000000000000,-447.000000000000,
-178.000000000000,-737.000000000000,
143.000000000000,177.000000000000,
572.000000000000,154.000000000000,
636.000000000000,-976.000000000000,
443.000000000000,706.000000000000,
545.000000000000,-133.000000000000,
435.000000000000,-1013.00000000000,
1158.00000000000,449.000000000000,
641.000000000000,30.0000000000000,
-671.000000000000,158.000000000000,
500.000000000000,322.000000000000,
574.000000000000,-199.000000000000,
-551.000000000000,-72.0000000000000,
-40.0000000000000,-492.000000000000,
367.000000000000,-89.0000000000000,
-306.000000000000,833.000000000000,
336.000000000000,1056.00000000000,
272.000000000000,219.000000000000,
-205.000000000000,113.000000000000,
-299.000000000000,706.000000000000,
-110.000000000000,585.000000000000,
-34.0000000000000,927.000000000000,
-310.000000000000,-411.000000000000,
450.000000000000,-509.000000000000,
-280.000000000000,871.000000000000,
238.000000000000,-470.000000000000,
1092.00000000000,-466.000000000000,
300.000000000000,880.000000000000,
663.000000000000,593.000000000000,
408.000000000000,-5.00000000000000,
857.000000000000,186.000000000000,
714.000000000000,-164.000000000000,
-1132.00000000000,450.000000000000,
-52.0000000000000,135.000000000000,
983.000000000000,-406.000000000000,
-378.000000000000,853.000000000000,
-230.000000000000,-324.000000000000,
27.0000000000000,-760.000000000000,
-437.000000000000,-98.0000000000000,
694.000000000000,-43.0000000000000,
580.000000000000,605.000000000000,
113.000000000000,-44.0000000000000,
17.0000000000000,-5.00000000000000,
-734.000000000000,702.000000000000,
-64.0000000000000,-353.000000000000,
505.000000000000,117.000000000000,
-565.000000000000,125.000000000000,
-599.000000000000,-318.000000000000,
-31.0000000000000,768.000000000000,
-86.0000000000000,797.000000000000,
251.000000000000,379.000000000000,
387.000000000000,-257.000000000000,
695.000000000000,394.000000000000,
-175.000000000000,22.0000000000000,
360.000000000000,-1114.00000000000,
447.000000000000,508.000000000000,
274.000000000000,293.000000000000,
-121.000000000000,-117.000000000000,
-278.000000000000,-556.000000000000,
1013.00000000000,-647.000000000000,
-116.000000000000,676.000000000000,
289.000000000000,-590.000000000000,
258.000000000000,-122.000000000000,
-901.000000000000,-84.0000000000000,
-268.000000000000,-739.000000000000,
620.000000000000,879.000000000000,
292.000000000000,146.000000000000,
321.000000000000,-260.000000000000,
391.000000000000,191.000000000000,
-853.000000000000,-15.0000000000000,
387.000000000000,-151.000000000000,
340.000000000000,9.00000000000000,
24.0000000000000,104.000000000000,
325.000000000000,-302.000000000000,
-583.000000000000,-122.000000000000,
-349.000000000000,-53.0000000000000,
-211.000000000000,449.000000000000,
61.0000000000000,-44.0000000000000,
-719.000000000000,-667.000000000000,
-341.000000000000,-614.000000000000,
593.000000000000,-202.000000000000,
706.000000000000,1585.00000000000,
548.000000000000,-614.000000000000,
120.000000000000,-405.000000000000,
86.0000000000000,1427.00000000000,
-768.000000000000,-761.000000000000,
379.000000000000,-801.000000000000,
-483.000000000000,-208.000000000000,
-913.000000000000,-162.000000000000,
353.000000000000,-499.000000000000,
-997.000000000000,-117.000000000000,
-307.000000000000,358.000000000000,
-501.000000000000,-448.000000000000,
-909.000000000000,-309.000000000000,
464.000000000000,202.000000000000,
-36.0000000000000,-652.000000000000,
81.0000000000000,-155.000000000000,
730.000000000000,42.0000000000000,
261.000000000000,-1083.00000000000,
237.000000000000,1074.00000000000,
414.000000000000,655.000000000000,
-368.000000000000,-659.000000000000,
124.000000000000,-609.000000000000,
870.000000000000,-1094.00000000000,
-884.000000000000,289.000000000000,
188.000000000000,-49.0000000000000,
749.000000000000,-162.000000000000,
316.000000000000,742.000000000000,
-259.000000000000,651.000000000000,
-1078.00000000000,26.0000000000000,
371.000000000000,-1667.00000000000,
141.000000000000,-549.000000000000,
-398.000000000000,798.000000000000,
552.000000000000,190.000000000000,
-38.0000000000000,699.000000000000,
-679.000000000000,321.000000000000,
-53.0000000000000,37.0000000000000,
-501.000000000000,768.000000000000,
232.000000000000,717.000000000000,
970.000000000000,-182.000000000000,
578.000000000000,108.000000000000,
202.000000000000,1129.00000000000,
-942.000000000000,-537.000000000000,
535.000000000000,-1124.00000000000,
684.000000000000,-412.000000000000,
-304.000000000000,609.000000000000,
-598.000000000000,59.0000000000000,
-1092.00000000000,117.000000000000,
-199.000000000000,696.000000000000,
-125.000000000000,-956.000000000000,
383.000000000000,876.000000000000,
-695.000000000000,-234.000000000000,
-326.000000000000,-230.000000000000,
520.000000000000,713.000000000000,
-713.000000000000,-410.000000000000,
-211.000000000000,546.000000000000,
-542.000000000000,-1045.00000000000,
199.000000000000,-672.000000000000,
-160.000000000000,-116.000000000000,
-453.000000000000,-40.0000000000000,
306.000000000000,-118.000000000000,
536.000000000000,-314.000000000000,
39.0000000000000,1174.00000000000,
-476.000000000000,237.000000000000,
226.000000000000,-907.000000000000,
-414.000000000000,-667.000000000000,
-197.000000000000,-671.000000000000,
349.000000000000,-1059.00000000000,
-99.0000000000000,-1080.00000000000,
646.000000000000,-213.000000000000,
974.000000000000,654.000000000000,
703.000000000000,25.0000000000000,
998.000000000000,136.000000000000,
68.0000000000000,768.000000000000,
-522.000000000000,-56.0000000000000,
-51.0000000000000,-261.000000000000,
426.000000000000,36.0000000000000,
23.0000000000000,319.000000000000,
-11.0000000000000,-283.000000000000,
-67.0000000000000,-356.000000000000,
-129.000000000000,568.000000000000,
194.000000000000,-1415.00000000000,
568.000000000000,-426.000000000000,
779.000000000000,928.000000000000,
-998.000000000000,421.000000000000,
-357.000000000000,1268.00000000000,
-678.000000000000,289.000000000000,
-705.000000000000,948.000000000000,
1008.00000000000,-641.000000000000,
837.000000000000,-547.000000000000,
1132.00000000000,1211.00000000000,
612.000000000000,-647.000000000000,
-545.000000000000,-122.000000000000,
-451.000000000000,-344.000000000000,
769.000000000000,-66.0000000000000,
-668.000000000000,142.000000000000,
-150.000000000000,-973.000000000000,
592.000000000000,756.000000000000,
-1328.00000000000,774.000000000000,
-491.000000000000,-541.000000000000,
1067.00000000000,-122.000000000000,
410.000000000000,535.000000000000,
-173.000000000000,734.000000000000,
878.000000000000,541.000000000000,
865.000000000000,779.000000000000,
-380.000000000000,1122.00000000000,
-582.000000000000,-384.000000000000,
90.0000000000000,-832.000000000000,
1296.00000000000,231.000000000000,
1209.00000000000,534.000000000000,
-33.0000000000000,193.000000000000,
571.000000000000,-785.000000000000,
-313.000000000000,146.000000000000,
73.0000000000000,-264.000000000000,
587.000000000000,-277.000000000000,
-238.000000000000,1549.00000000000,
-55.0000000000000,648.000000000000,
-1094.00000000000,533.000000000000,
-429.000000000000,-2.00000000000000,
66.0000000000000,-822.000000000000,
596.000000000000,-694.000000000000,
292.000000000000,132.000000000000,
-668.000000000000,629.000000000000,
-547.000000000000,431.000000000000,
-714.000000000000,-38.0000000000000,
674.000000000000,-394.000000000000,
-100.000000000000,1134.00000000000,
-78.0000000000000,714.000000000000,
1139.00000000000,-184.000000000000,
160.000000000000,619.000000000000,
-470.000000000000,976.000000000000,
-1340.00000000000,-328.000000000000,
-613.000000000000,-510.000000000000,
-161.000000000000,62.0000000000000,
-163.000000000000,-832.000000000000,
802.000000000000,259.000000000000,
-188.000000000000,-302.000000000000,
-272.000000000000,-11.0000000000000,
18.0000000000000,1190.00000000000,
-1073.00000000000,-814.000000000000,
188.000000000000,-617.000000000000,
1501.00000000000,186.000000000000,
-151.000000000000,-765.000000000000,
-53.0000000000000,23.0000000000000,
570.000000000000,467.000000000000,
84.0000000000000,71.0000000000000,
466.000000000000,-629.000000000000,
278.000000000000,-348.000000000000,
679.000000000000,613.000000000000,
-349.000000000000,475.000000000000,
-1218.00000000000,713.000000000000,
-490.000000000000,-957.000000000000,
302.000000000000,-1193.00000000000,
319.000000000000,-230.000000000000,
805.000000000000,-181.000000000000,
28.0000000000000,446.000000000000,
-554.000000000000,-488.000000000000,
19.0000000000000,-832.000000000000,
-94.0000000000000,-565.000000000000,
1121.00000000000,-219.000000000000,
47.0000000000000,74.0000000000000,
-598.000000000000,607.000000000000,
426.000000000000,342.000000000000,
692.000000000000,-952.000000000000,
192.000000000000,804.000000000000,
-182.000000000000,395.000000000000,
774.000000000000,219.000000000000,
-320.000000000000,1714.00000000000,
-975.000000000000,257.000000000000,
-529.000000000000,-380.000000000000,
-383.000000000000,-495.000000000000,
500.000000000000,-645.000000000000,
83.0000000000000,479.000000000000,
640.000000000000,-22.0000000000000,
842.000000000000,-349.000000000000,
-680.000000000000,963.000000000000,
524.000000000000,-1175.00000000000,
-697.000000000000,-602.000000000000,
86.0000000000000,-190.000000000000,
611.000000000000,-1067.00000000000,
-1284.00000000000,653.000000000000,
-323.000000000000,-624.000000000000,
-977.000000000000,-450.000000000000,
336.000000000000,-505.000000000000,
132.000000000000,-618.000000000000,
-684.000000000000,651.000000000000,
-78.0000000000000,639.000000000000,
-686.000000000000,8.00000000000000,
-50.0000000000000,-1700.00000000000,
642.000000000000,-645.000000000000,
227.000000000000,-378.000000000000,
643.000000000000,-554.000000000000,
537.000000000000,1289.00000000000,
-333.000000000000,376.000000000000,
520.000000000000,577.000000000000,
-310.000000000000,-103.000000000000,
-385.000000000000,-1366.00000000000,
-292.000000000000,-262.000000000000,
-519.000000000000,-1238.00000000000,
1109.00000000000,-1012.00000000000,
325.000000000000,757.000000000000,
-1330.00000000000,189.000000000000,
-400.000000000000,220.000000000000,
1104.00000000000,406.000000000000,
189.000000000000,-252.000000000000,
-1185.00000000000,102.000000000000,
167.000000000000,-393.000000000000,
89.0000000000000,490.000000000000,
-560.000000000000,357.000000000000,
-39.0000000000000,-1619.00000000000,
103.000000000000,319.000000000000,
1375.00000000000,161.000000000000,
170.000000000000,-523.000000000000,
310.000000000000,341.000000000000,
200.000000000000,252.000000000000,
-483.000000000000,-348.000000000000,
293.000000000000,-1596.00000000000,
352.000000000000,-39.0000000000000,
-221.000000000000,589.000000000000,
-883.000000000000,168.000000000000,
1319.00000000000,625.000000000000,
-207.000000000000,1000.00000000000,
-784.000000000000,-429.000000000000,
596.000000000000,-824.000000000000,
-1182.00000000000,193.000000000000,
-377.000000000000,-458.000000000000,
-487.000000000000,222.000000000000,
-962.000000000000,-902.000000000000,
431.000000000000,-1319.00000000000,
653.000000000000,311.000000000000,
255.000000000000,-474.000000000000,
493.000000000000,-270.000000000000,
-235.000000000000,574.000000000000,
-876.000000000000,898.000000000000,
-858.000000000000,-88.0000000000000,
-1128.00000000000,-1007.00000000000,
-80.0000000000000,309.000000000000,
397.000000000000,-70.0000000000000,
693.000000000000,676.000000000000,
-66.0000000000000,1095.00000000000,
-536.000000000000,-207.000000000000,
952.000000000000,-44.0000000000000,
836.000000000000,458.000000000000,
859.000000000000,543.000000000000,
416.000000000000,-275.000000000000,
145.000000000000,-418.000000000000,
-304.000000000000,-1013.00000000000,
-596.000000000000,173.000000000000,
-70.0000000000000,-260.000000000000,
136.000000000000,-1133.00000000000,
1208.00000000000,584.000000000000,
-651.000000000000,-182.000000000000,
-576.000000000000,804.000000000000,
369.000000000000,-853.000000000000,
-7.00000000000000,-535.000000000000,
629.000000000000,1119.00000000000,
304.000000000000,78.0000000000000,
63.0000000000000,1242.00000000000,
-764.000000000000,-296.000000000000,
986.000000000000,-322.000000000000,
-175.000000000000,-543.000000000000,
-936.000000000000,211.000000000000,
1158.00000000000,188.000000000000,
-1704.00000000000,-863.000000000000,
-594.000000000000,-257.000000000000,
-457.000000000000,-471.000000000000,
-589.000000000000,553.000000000000,
1129.00000000000,226.000000000000,
-120.000000000000,695.000000000000,
717.000000000000,525.000000000000,
-96.0000000000000,757.000000000000,
-626.000000000000,-90.0000000000000,
-22.0000000000000,-535.000000000000,
140.000000000000,73.0000000000000,
382.000000000000,-1524.00000000000,
314.000000000000,126.000000000000,
479.000000000000,646.000000000000,
-562.000000000000,894.000000000000,
135.000000000000,1024.00000000000,
-543.000000000000,48.0000000000000,
353.000000000000,576.000000000000,
611.000000000000,-48.0000000000000,
-1150.00000000000,75.0000000000000,
90.0000000000000,-700.000000000000,
161.000000000000,-250.000000000000,
44.0000000000000,622.000000000000,
-348.000000000000,-943.000000000000,
513.000000000000,-947.000000000000,
1459.00000000000,445.000000000000,
-248.000000000000,499.000000000000,
-215.000000000000,-329.000000000000,
855.000000000000,468.000000000000,
1023.00000000000,673.000000000000,
391.000000000000,728.000000000000,
-357.000000000000,-169.000000000000,
-110.000000000000,-596.000000000000,
1129.00000000000,863.000000000000,
276.000000000000,79.0000000000000,
-1243.00000000000,19.0000000000000,
169.000000000000,824.000000000000,
458.000000000000,286.000000000000,
426.000000000000,394.000000000000,
61.0000000000000,814.000000000000,
-1239.00000000000,-162.000000000000,
388.000000000000,-756.000000000000,
399.000000000000,-743.000000000000,
-370.000000000000,-313.000000000000,
117.000000000000,759.000000000000,
-344.000000000000,462.000000000000,
-227.000000000000,787.000000000000,
4.00000000000000,-447.000000000000,
615.000000000000,-179.000000000000,
-94.0000000000000,721.000000000000,
-711.000000000000,-714.000000000000,
1175.00000000000,360.000000000000,
578.000000000000,978.000000000000,
-96.0000000000000,-229.000000000000,
428.000000000000,-511.000000000000,
163.000000000000,229.000000000000,
35.0000000000000,41.0000000000000,
-834.000000000000,-56.0000000000000,
-595.000000000000,-66.0000000000000,
-392.000000000000,-67.0000000000000,
-592.000000000000,-284.000000000000,
994.000000000000,-586.000000000000,
503.000000000000,685.000000000000,
-626.000000000000,947.000000000000,
694.000000000000,-663.000000000000,
-588.000000000000,-562.000000000000,
-340.000000000000,-683.000000000000,
728.000000000000,-1684.00000000000,
897.000000000000,162.000000000000,
1302.00000000000,-175.000000000000,
48.0000000000000,-144.000000000000,
-29.0000000000000,-397.000000000000,
-837.000000000000,19.0000000000000,
-246.000000000000,645.000000000000,
188.000000000000,-1080.00000000000,
694.000000000000,-429.000000000000,
1063.00000000000,-442.000000000000,
-102.000000000000,-33.0000000000000,
269.000000000000,544.000000000000,
-693.000000000000,875.000000000000,
-575.000000000000,353.000000000000,
-900.000000000000,-742.000000000000,
-150.000000000000,566.000000000000,
216.000000000000,-635.000000000000,
-940.000000000000,-497.000000000000,
-489.000000000000,-724.000000000000,
-1105.00000000000,-809.000000000000,
736.000000000000,-411.000000000000,
738.000000000000,-909.000000000000,
393.000000000000,1068.00000000000,
551.000000000000,-277.000000000000,
-446.000000000000,-505.000000000000,
51.0000000000000,-88.0000000000000,
574.000000000000,-508.000000000000,
421.000000000000,540.000000000000,
-1117.00000000000,232.000000000000,
-876.000000000000,261.000000000000,
-900.000000000000,-430.000000000000,
-581.000000000000,431.000000000000,
256.000000000000,329.000000000000,
-82.0000000000000,-711.000000000000,
231.000000000000,370.000000000000,
-194.000000000000,373.000000000000,
493.000000000000,-348.000000000000,
831.000000000000,-10.0000000000000,
-263.000000000000,96.0000000000000,
-728.000000000000,-988.000000000000,
107.000000000000,-72.0000000000000,
521.000000000000,460.000000000000,
-834.000000000000,51.0000000000000,
-571.000000000000,295.000000000000,
242.000000000000,-613.000000000000,
861.000000000000,-142.000000000000,
1027.00000000000,-301.000000000000,
-191.000000000000,-544.000000000000,
-34.0000000000000,161.000000000000,
-787.000000000000,-422.000000000000,
-1441.00000000000,-405.000000000000,
186.000000000000,316.000000000000,
475.000000000000,-629.000000000000,
-12.0000000000000,106.000000000000,
209.000000000000,1214.00000000000,
738.000000000000,-268.000000000000,
186.000000000000,834.000000000000,
792.000000000000,878.000000000000,
26.0000000000000,-747.000000000000,
-930.000000000000,-7.00000000000000,
987.000000000000,-508.000000000000,
443.000000000000,-21.0000000000000,
163.000000000000,-874.000000000000,
1111.00000000000,-1287.00000000000,
200.000000000000,342.000000000000,
-697.000000000000,-746.000000000000,
813.000000000000,265.000000000000,
98.0000000000000,1074.00000000000,
-812.000000000000,1203.00000000000,
29.0000000000000,716.000000000000,
-490.000000000000,-1386.00000000000,
1017.00000000000,-355.000000000000,
1252.00000000000,-229.000000000000,
697.000000000000,266.000000000000,
350.000000000000,1016.00000000000,
-1062.00000000000,29.0000000000000,
-997.000000000000,-36.0000000000000,
-746.000000000000,274.000000000000,
-766.000000000000,401.000000000000,
-236.000000000000,60.0000000000000,
-66.0000000000000,140.000000000000,
-692.000000000000,-119.000000000000,
288.000000000000,-537.000000000000,
1029.00000000000,-1442.00000000000,
-343.000000000000,-115.000000000000,
328.000000000000,207.000000000000,
-120.000000000000,-826.000000000000,
-315.000000000000,611.000000000000,
62.0000000000000,-164.000000000000,
-512.000000000000,17.0000000000000,
79.0000000000000,765.000000000000,
-829.000000000000,475.000000000000,
-478.000000000000,-120.000000000000,
20.0000000000000,-798.000000000000,
178.000000000000,571.000000000000,
-36.0000000000000,-112.000000000000,
-660.000000000000,73.0000000000000,
-282.000000000000,126.000000000000,
-135.000000000000,242.000000000000,
847.000000000000,710.000000000000,
962.000000000000,-375.000000000000,
445.000000000000,886.000000000000,
-819.000000000000,13.0000000000000,
300.000000000000,-1064.00000000000,
1180.00000000000,-765.000000000000,
-640.000000000000,-323.000000000000,
775.000000000000,-55.0000000000000,
-433.000000000000,498.000000000000,
-405.000000000000,737.000000000000,
910.000000000000,-211.000000000000,
-351.000000000000,1526.00000000000,
-448.000000000000,-290.000000000000,
-819.000000000000,-872.000000000000,
181.000000000000,316.000000000000,
-233.000000000000,-190.000000000000,
-574.000000000000,581.000000000000,
309.000000000000,-626.000000000000,
849.000000000000,264.000000000000,
813.000000000000,1034.00000000000,
-483.000000000000,332.000000000000,
-193.000000000000,831.000000000000,
19.0000000000000,101.000000000000,
230.000000000000,-486.000000000000,
64.0000000000000,225.000000000000,
153.000000000000,487.000000000000,
386.000000000000,483.000000000000,
-774.000000000000,677.000000000000,
-275.000000000000,-1013.00000000000,
-248.000000000000,181.000000000000,
-451.000000000000,1458.00000000000,
-971.000000000000,-332.000000000000,
-671.000000000000,1110.00000000000,
149.000000000000,-432.000000000000,
206.000000000000,-1354.00000000000,
600.000000000000,-381.000000000000,
160.000000000000,-855.000000000000,
795.000000000000,457.000000000000,
-39.0000000000000,-247.000000000000,
288.000000000000,248.000000000000,
680.000000000000,1067.00000000000,
-319.000000000000,534.000000000000,
914.000000000000,860.000000000000,
435.000000000000,295.000000000000,
-495.000000000000,-113.000000000000,
554.000000000000,-74.0000000000000,
-98.0000000000000,-756.000000000000,
-629.000000000000,317.000000000000,
-132.000000000000,223.000000000000,
-120.000000000000,-233.000000000000,
-450.000000000000,1225.00000000000,
-1036.00000000000,-383.000000000000,
491.000000000000,-614.000000000000,
924.000000000000,816.000000000000,
-413.000000000000,-252.000000000000,
643.000000000000,-607.000000000000,
660.000000000000,670.000000000000,
-1088.00000000000,697.000000000000,
-456.000000000000,120.000000000000,
385.000000000000,-246.000000000000,
-93.0000000000000,-496.000000000000,
-260.000000000000,626.000000000000,
-427.000000000000,533.000000000000,
267.000000000000,-890.000000000000,
37.0000000000000,395.000000000000,
-775.000000000000,1065.00000000000,
56.0000000000000,2.00000000000000,
413.000000000000,778.000000000000,
-951.000000000000,372.000000000000,
-901.000000000000,179.000000000000,
-203.000000000000,-171.000000000000,
-229.000000000000,47.0000000000000,
686.000000000000,328.000000000000,
189.000000000000,-1265.00000000000,
1212.00000000000,389.000000000000,
1226.00000000000,539.000000000000,
-211.000000000000,-99.0000000000000,
127.000000000000,193.000000000000,
-635.000000000000,1181.00000000000,
62.0000000000000,653.000000000000,
-863.000000000000,-599.000000000000,
220.000000000000,359.000000000000,
737.000000000000,-729.000000000000,
-775.000000000000,229.000000000000,
1169.00000000000,-437.000000000000,
-147.000000000000,208.000000000000,
-495.000000000000,1570.00000000000,
279.000000000000,-339.000000000000,
174.000000000000,763.000000000000,
-589.000000000000,1222.00000000000,
-959.000000000000,29.0000000000000,
-412.000000000000,-841.000000000000,
-473.000000000000,576.000000000000,
776.000000000000,-60.0000000000000,
288.000000000000,-1286.00000000000,
529.000000000000,-105.000000000000,
548.000000000000,-598.000000000000,
118.000000000000,-777.000000000000,
1087.00000000000,-2.00000000000000,
-391.000000000000,226.000000000000,
274.000000000000,-235.000000000000,
318.000000000000,588.000000000000,
473.000000000000,27.0000000000000,
235.000000000000,-71.0000000000000,
-508.000000000000,901.000000000000,
987.000000000000,158.000000000000,
-911.000000000000,963.000000000000,
223.000000000000,-983.000000000000,
-10.0000000000000,-445.000000000000,
-823.000000000000,20.0000000000000,
-653.000000000000,-1213.00000000000,
-339.000000000000,660.000000000000,
1380.00000000000,-18.0000000000000,
-862.000000000000,375.000000000000,
636.000000000000,-454.000000000000,
-229.000000000000,-610.000000000000,
242.000000000000,-356.000000000000,
987.000000000000,100.000000000000,
-720.000000000000,1686.00000000000,
792.000000000000,-754.000000000000,
-452.000000000000,-86.0000000000000,
-704.000000000000,109.000000000000,
-666.000000000000,-525.000000000000,
665.000000000000,358.000000000000,
1204.00000000000,-386.000000000000,
417.000000000000,662.000000000000,
86.0000000000000,1172.00000000000,
-1077.00000000000,207.000000000000,
-478.000000000000,-412.000000000000,
-71.0000000000000,-208.000000000000,
269.000000000000,-106.000000000000,
475.000000000000,158.000000000000,
-65.0000000000000,357.000000000000,
381.000000000000,113.000000000000,
600.000000000000,163.000000000000,
-570.000000000000,-238.000000000000,
325.000000000000,-255.000000000000,
297.000000000000,193.000000000000,
-599.000000000000,241.000000000000,
867.000000000000,130.000000000000,
239.000000000000,100.000000000000,
-116.000000000000,-110.000000000000,
739.000000000000,-639.000000000000,
158.000000000000,-1243.00000000000,
738.000000000000,-265.000000000000,
166.000000000000,1053.00000000000,
-838.000000000000,-176.000000000000,
422.000000000000,-354.000000000000,
380.000000000000,-240.000000000000,
487.000000000000,-226.000000000000,
-730.000000000000,410.000000000000,
88.0000000000000,-950.000000000000,
1299.00000000000,77.0000000000000,
-396.000000000000,1104.00000000000,
-104.000000000000,493.000000000000,
-798.000000000000,11.0000000000000,
-802.000000000000,-314.000000000000,
176.000000000000,964.000000000000,
-492.000000000000,115.000000000000,
-683.000000000000,-272.000000000000,
357.000000000000,-41.0000000000000,
-419.000000000000,-1221.00000000000,
-183.000000000000,465.000000000000,
651.000000000000,332.000000000000,
-522.000000000000,211.000000000000,
-3.00000000000000,928.000000000000,
-389.000000000000,-814.000000000000,
302.000000000000,486.000000000000,
1076.00000000000,239.000000000000,
124.000000000000,-14.0000000000000,
-507.000000000000,440.000000000000,
-610.000000000000,107.000000000000,
1010.00000000000,378.000000000000,
-364.000000000000,297.000000000000,
-433.000000000000,490.000000000000,
55.0000000000000,502.000000000000,
-1274.00000000000,367.000000000000,
-494.000000000000,-1344.00000000000,
-323.000000000000,-161.000000000000,
77.0000000000000,860.000000000000,
-487.000000000000,69.0000000000000,
-550.000000000000,39.0000000000000,
-612.000000000000,-741.000000000000,
-22.0000000000000,-310.000000000000,
1318.00000000000,-168.000000000000,
658.000000000000,998.000000000000,
469.000000000000,687.000000000000,
-1120.00000000000,290.000000000000,
-422.000000000000,150.000000000000,
7.00000000000000,-1084.00000000000,
494.000000000000,704.000000000000,
1052.00000000000,-161.000000000000,
-878.000000000000,363.000000000000,
-578.000000000000,356.000000000000,
-470.000000000000,-1368.00000000000,
399.000000000000,920.000000000000,
-249.000000000000,-94.0000000000000,
-936.000000000000,-648.000000000000,
277.000000000000,-213.000000000000,
512.000000000000,110.000000000000,
-150.000000000000,-159.000000000000,
60.0000000000000,-815.000000000000,
386.000000000000,880.000000000000,
-544.000000000000,233.000000000000,
438.000000000000,-591.000000000000,
125.000000000000,-274.000000000000,
-563.000000000000,786.000000000000,
-422.000000000000,48.0000000000000,
-30.0000000000000,-1002.00000000000,
749.000000000000,168.000000000000,
-477.000000000000,-220.000000000000,
-756.000000000000,-550.000000000000,
-583.000000000000,-183.000000000000,
63.0000000000000,307.000000000000,
582.000000000000,868.000000000000,
-826.000000000000,474.000000000000,
-642.000000000000,-41.0000000000000,
-309.000000000000,372.000000000000,
-1176.00000000000,-207.000000000000,
-439.000000000000,-136.000000000000,
158.000000000000,779.000000000000,
99.0000000000000,-587.000000000000,
-627.000000000000,-513.000000000000,
-425.000000000000,-550.000000000000,
315.000000000000,-969.000000000000,
390.000000000000,440.000000000000,
-334.000000000000,-648.000000000000,
62.0000000000000,-1000.00000000000,
843.000000000000,-677.000000000000,
-49.0000000000000,-611.000000000000,
140.000000000000,-549.000000000000,
-147.000000000000,-877.000000000000,
365.000000000000,429.000000000000,
819.000000000000,163.000000000000,
106.000000000000,33.0000000000000,
403.000000000000,967.000000000000,
218.000000000000,-106.000000000000,
44.0000000000000,-212.000000000000,
287.000000000000,744.000000000000,
-752.000000000000,-56.0000000000000,
-606.000000000000,-348.000000000000,
754.000000000000,-425.000000000000,
271.000000000000,412.000000000000,
-498.000000000000,954.000000000000,
360.000000000000,-53.0000000000000,
370.000000000000,442.000000000000,
420.000000000000,-259.000000000000,
701.000000000000,-417.000000000000,
-665.000000000000,197.000000000000,
-416.000000000000,-1011.00000000000,
211.000000000000,-987.000000000000,
912.000000000000,-581.000000000000,
-600.000000000000,270.000000000000,
-93.0000000000000,-454.000000000000,
723.000000000000,-730.000000000000,
-845.000000000000,143.000000000000,
347.000000000000,-685.000000000000,
-928.000000000000,-10.0000000000000,
641.000000000000,352.000000000000,
1159.00000000000,-76.0000000000000,
-558.000000000000,-133.000000000000,
445.000000000000,290.000000000000,
223.000000000000,-28.0000000000000,
235.000000000000,-396.000000000000,
548.000000000000,1109.00000000000,
231.000000000000,-377.000000000000,
-1062.00000000000,-106.000000000000,
-128.000000000000,1189.00000000000,
-720.000000000000,-414.000000000000,
-734.000000000000,-620.000000000000,
562.000000000000,-415.000000000000,
-643.000000000000,461.000000000000,
795.000000000000,-220.000000000000,
97.0000000000000,-176.000000000000,
247.000000000000,1169.00000000000,
556.000000000000,-61.0000000000000,
-233.000000000000,-37.0000000000000,
251.000000000000,354.000000000000,
-491.000000000000,-454.000000000000,
1079.00000000000,-287.000000000000,
128.000000000000,765.000000000000,
-928.000000000000,-399.000000000000,
275.000000000000,351.000000000000,
-417.000000000000,27.0000000000000,
-518.000000000000,-1450.00000000000,
-103.000000000000,578.000000000000,
-21.0000000000000,492.000000000000,
-498.000000000000,351.000000000000,
669.000000000000,850.000000000000,
435.000000000000,374.000000000000,
-458.000000000000,697.000000000000,
344.000000000000,391.000000000000,
280.000000000000,-331.000000000000,
368.000000000000,-1085.00000000000,
291.000000000000,-5.00000000000000,
149.000000000000,1112.00000000000,
-1111.00000000000,446.000000000000,
-336.000000000000,592.000000000000,
265.000000000000,627.000000000000,
-1231.00000000000,1107.00000000000,
-335.000000000000,611.000000000000,
169.000000000000,-531.000000000000,
-267.000000000000,-181.000000000000,
-1195.00000000000,-17.0000000000000,
-686.000000000000,-1059.00000000000,
864.000000000000,-425.000000000000,
333.000000000000,276.000000000000,
60.0000000000000,-747.000000000000,
-147.000000000000,314.000000000000,
-411.000000000000,277.000000000000,
-363.000000000000,-904.000000000000,
847.000000000000,-262.000000000000,
696.000000000000,679.000000000000,
-857.000000000000,797.000000000000,
-774.000000000000,-506.000000000000,
-744.000000000000,-295.000000000000,
645.000000000000,-34.0000000000000,
299.000000000000,-121.000000000000,
437.000000000000,698.000000000000,
775.000000000000,591.000000000000,
-1756.00000000000,6.00000000000000,
-816.000000000000,-120.000000000000,
2.00000000000000,-62.0000000000000,
-405.000000000000,-184.000000000000,
509.000000000000,273.000000000000,
-128.000000000000,170.000000000000,
-665.000000000000,-609.000000000000,
662.000000000000,-692.000000000000,
391.000000000000,-1130.00000000000,
-75.0000000000000,-313.000000000000,
515.000000000000,-127.000000000000,
870.000000000000,-158.000000000000,
336.000000000000,950.000000000000,
-1484.00000000000,-119.000000000000,
-65.0000000000000,-61.0000000000000,
979.000000000000,79.0000000000000,
-648.000000000000,-26.0000000000000,
-109.000000000000,935.000000000000,
-1255.00000000000,103.000000000000,
-211.000000000000,-694.000000000000,
215.000000000000,-61.0000000000000,
-1150.00000000000,-298.000000000000,
1196.00000000000,-382.000000000000,
499.000000000000,520.000000000000,
159.000000000000,-549.000000000000,
754.000000000000,297.000000000000,
795.000000000000,805.000000000000,
294.000000000000,9.00000000000000,
-450.000000000000,137.000000000000,
713.000000000000,-420.000000000000,
216.000000000000,666.000000000000,
-203.000000000000,701.000000000000,
-395.000000000000,589.000000000000,
93.0000000000000,685.000000000000,
-394.000000000000,-163.000000000000,
-545.000000000000,-486.000000000000,
815.000000000000,-860.000000000000,
253.000000000000,501.000000000000,
-787.000000000000,457.000000000000,
30.0000000000000,-400.000000000000,
498.000000000000,766.000000000000,
-359.000000000000,96.0000000000000,
322.000000000000,83.0000000000000,
-916.000000000000,35.0000000000000,
-952.000000000000,-262.000000000000,
855.000000000000,-553.000000000000,
-591.000000000000,-424.000000000000,
-627.000000000000,435.000000000000,
-38.0000000000000,60.0000000000000,
-413.000000000000,157.000000000000,
281.000000000000,-752.000000000000,
463.000000000000,238.000000000000,
-329.000000000000,817.000000000000,
423.000000000000,13.0000000000000,
160.000000000000,1120.00000000000,
-905.000000000000,594.000000000000,
787.000000000000,170.000000000000,
31.0000000000000,-814.000000000000,
-257.000000000000,-141.000000000000,
591.000000000000,163.000000000000,
229.000000000000,94.0000000000000,
1526.00000000000,479.000000000000,
-709.000000000000,407.000000000000,
-348.000000000000,816.000000000000,
837.000000000000,-184.000000000000,
-431.000000000000,879.000000000000,
1109.00000000000,133.000000000000,
-179.000000000000,228.000000000000,
-231.000000000000,1042.00000000000,
269.000000000000,-226.000000000000,
261.000000000000,780.000000000000,
48.0000000000000,974.000000000000,
-517.000000000000,164.000000000000,
1062.00000000000,-54.0000000000000,
-647.000000000000,514.000000000000,
-1162.00000000000,-368.000000000000,
-489.000000000000,-112.000000000000,
-673.000000000000,-265.000000000000,
-942.000000000000,-904.000000000000,
-418.000000000000,-177.000000000000,
774.000000000000,-914.000000000000,
-999.000000000000,-526.000000000000,
-416.000000000000,-320.000000000000,
-467.000000000000,-157.000000000000,
-1025.00000000000,-30.0000000000000,
-210.000000000000,-312.000000000000,
-487.000000000000,-77.0000000000000,
441.000000000000,-243.000000000000,
754.000000000000,71.0000000000000,
-415.000000000000,-488.000000000000,
-1179.00000000000,-689.000000000000,
277.000000000000,-609.000000000000,
1015.00000000000,-100.000000000000,
850.000000000000,1028.00000000000,
556.000000000000,142.000000000000,
-733.000000000000,-1.00000000000000,
-768.000000000000,-718.000000000000,
-410.000000000000,-802.000000000000,
423.000000000000,748.000000000000,
71.0000000000000,-557.000000000000,
-211.000000000000,200.000000000000,
21.0000000000000,1323.00000000000,
-386.000000000000,120.000000000000,
247.000000000000,196.000000000000,
664.000000000000,453.000000000000,
-409.000000000000,111.000000000000,
-697.000000000000,-608.000000000000,
263.000000000000,134.000000000000,
-161.000000000000,1013.00000000000,
-606.000000000000,107.000000000000,
-564.000000000000,-497.000000000000,
80.0000000000000,-544.000000000000,
-128.000000000000,-805.000000000000,
297.000000000000,-270.000000000000,
780.000000000000,548.000000000000,
-832.000000000000,1166.00000000000,
-333.000000000000,922.000000000000,
246.000000000000,430.000000000000,
-448.000000000000,-526.000000000000,
444.000000000000,-507.000000000000,
1013.00000000000,543.000000000000,
368.000000000000,-37.0000000000000,
731.000000000000,558.000000000000,
-502.000000000000,294.000000000000,
-570.000000000000,-842.000000000000,
743.000000000000,-452.000000000000,
49.0000000000000,-835.000000000000,
-433.000000000000,-671.000000000000,
658.000000000000,-842.000000000000,
330.000000000000,326.000000000000,
-1093.00000000000,282.000000000000,
888.000000000000,-703.000000000000,
-209.000000000000,483.000000000000,
-1060.00000000000,35.0000000000000,
500.000000000000,-256.000000000000,
-861.000000000000,-88.0000000000000,
-497.000000000000,-613.000000000000,
437.000000000000,-980.000000000000,
346.000000000000,-538.000000000000,
485.000000000000,174.000000000000,
-459.000000000000,-239.000000000000,
72.0000000000000,-764.000000000000,
844.000000000000,-245.000000000000,
654.000000000000,257.000000000000,
411.000000000000,199.000000000000,
-219.000000000000,1172.00000000000,
232.000000000000,-344.000000000000,
487.000000000000,-528.000000000000,
240.000000000000,984.000000000000,
164.000000000000,-872.000000000000,
-228.000000000000,-321.000000000000,
-700.000000000000,915.000000000000,
-626.000000000000,747.000000000000,
-973.000000000000,30.0000000000000,
183.000000000000,-1024.00000000000,
-21.0000000000000,-206.000000000000,
-1139.00000000000,-221.000000000000,
233.000000000000,272.000000000000,
-208.000000000000,49.0000000000000,
136.000000000000,-1456.00000000000,
1098.00000000000,-614.000000000000,
-141.000000000000,646.000000000000,
-62.0000000000000,812.000000000000,
9.00000000000000,417.000000000000,
-1532.00000000000,-393.000000000000,
-465.000000000000,234.000000000000,
867.000000000000,-186.000000000000,
71.0000000000000,-389.000000000000,
-218.000000000000,891.000000000000,
141.000000000000,509.000000000000,
-125.000000000000,183.000000000000,
-1171.00000000000,-803.000000000000,
-682.000000000000,-24.0000000000000,
-644.000000000000,-74.0000000000000,
43.0000000000000,-874.000000000000,
1430.00000000000,-341.000000000000,
-484.000000000000,111.000000000000,
-108.000000000000,467.000000000000,
34.0000000000000,-247.000000000000,
-1045.00000000000,193.000000000000,
-5.00000000000000,-774.000000000000,
355.000000000000,-798.000000000000,
651.000000000000,458.000000000000,
-159.000000000000,892.000000000000,
-612.000000000000,671.000000000000,
-211.000000000000,-24.0000000000000,
968.000000000000,84.0000000000000,
752.000000000000,-406.000000000000,
-843.000000000000,732.000000000000,
-198.000000000000,997.000000000000,
-347.000000000000,387.000000000000,
-602.000000000000,782.000000000000,
-22.0000000000000,-204.000000000000,
-138.000000000000,-804.000000000000,
218.000000000000,-695.000000000000,
1161.00000000000,226.000000000000,
-16.0000000000000,-128.000000000000,
-186.000000000000,-337.000000000000,
1518.00000000000,727.000000000000,
-399.000000000000,238.000000000000,
-510.000000000000,-444.000000000000,
862.000000000000,-859.000000000000,
253.000000000000,860.000000000000,
1019.00000000000,854.000000000000,
849.000000000000,166.000000000000,
-414.000000000000,532.000000000000,
-411.000000000000,-1026.00000000000,
832.000000000000,-897.000000000000,
-150.000000000000,-603.000000000000,
-421.000000000000,-78.0000000000000,
878.000000000000,-370.000000000000,
-798.000000000000,268.000000000000,
-1020.00000000000,287.000000000000,
-567.000000000000,-1208.00000000000,
428.000000000000,206.000000000000,
340.000000000000,-404.000000000000,
-155.000000000000,-1198.00000000000,
866.000000000000,165.000000000000,
-885.000000000000,496.000000000000,
-297.000000000000,-440.000000000000,
851.000000000000,472.000000000000,
-529.000000000000,-25.0000000000000,
-75.0000000000000,-1479.00000000000,
691.000000000000,734.000000000000,
-211.000000000000,458.000000000000,
194.000000000000,-357.000000000000,
855.000000000000,402.000000000000,
-790.000000000000,30.0000000000000,
-253.000000000000,802.000000000000,
-647.000000000000,445.000000000000,
-908.000000000000,-200.000000000000,
976.000000000000,-1094.00000000000,
7.00000000000000,-137.000000000000,
-676.000000000000,116.000000000000,
306.000000000000,-1269.00000000000,
1017.00000000000,995.000000000000,
386.000000000000,675.000000000000,
-24.0000000000000,-424.000000000000,
-239.000000000000,229.000000000000,
-51.0000000000000,1209.00000000000,
253.000000000000,-122.000000000000,
420.000000000000,-1110.00000000000,
761.000000000000,714.000000000000,
-958.000000000000,-598.000000000000,
-161.000000000000,-926.000000000000,
703.000000000000,-192.000000000000,
-199.000000000000,87.0000000000000,
756.000000000000,-524.000000000000,
-230.000000000000,-645.000000000000,
419.000000000000,545.000000000000,
-171.000000000000,588.000000000000,
-1013.00000000000,255.000000000000,
365.000000000000,-1449.00000000000,
-715.000000000000,-11.0000000000000,
-188.000000000000,590.000000000000,
-343.000000000000,-676.000000000000,
902.000000000000,-459.000000000000,
637.000000000000,30.0000000000000,
-953.000000000000,347.000000000000,
544.000000000000,-1510.00000000000,
518.000000000000,-396.000000000000,
707.000000000000,-792.000000000000,
293.000000000000,-667.000000000000,
-117.000000000000,913.000000000000,
-497.000000000000,-983.000000000000,
722.000000000000,877.000000000000,
314.000000000000,-123.000000000000,
17.0000000000000,-292.000000000000,
448.000000000000,148.000000000000,
-901.000000000000,-763.000000000000,
468.000000000000,1095.00000000000,
-808.000000000000,320.000000000000,
-422.000000000000,544.000000000000,
904.000000000000,808.000000000000,
-747.000000000000,-20.0000000000000,
284.000000000000,-305.000000000000,
106.000000000000,828.000000000000,
-1058.00000000000,202.000000000000,
-450.000000000000,-879.000000000000,
969.000000000000,340.000000000000,
127.000000000000,-518.000000000000,
-399.000000000000,-56.0000000000000,
753.000000000000,556.000000000000,
-501.000000000000,397.000000000000,
-306.000000000000,173.000000000000,
93.0000000000000,309.000000000000,
-394.000000000000,968.000000000000,
-861.000000000000,-644.000000000000,
-455.000000000000,726.000000000000,
-189.000000000000,289.000000000000,
-438.000000000000,-150.000000000000,
995.000000000000,849.000000000000,
-192.000000000000,-141.000000000000,
442.000000000000,700.000000000000,
737.000000000000,-689.000000000000,
-387.000000000000,-367.000000000000,
221.000000000000,230.000000000000,
362.000000000000,-560.000000000000,
340.000000000000,-58.0000000000000,
-752.000000000000,206.000000000000,
-681.000000000000,947.000000000000,
41.0000000000000,531.000000000000,
246.000000000000,551.000000000000,
-30.0000000000000,-262.000000000000,
-317.000000000000,-110.000000000000,
914.000000000000,623.000000000000,
655.000000000000,523.000000000000,
622.000000000000,1060.00000000000,
621.000000000000,771.000000000000,
24.0000000000000,232.000000000000,
-785.000000000000,238.000000000000,
-1406.00000000000,35.0000000000000,
628.000000000000,-658.000000000000,
-624.000000000000,133.000000000000,
-701.000000000000,-193.000000000000,
-8.00000000000000,-205.000000000000,
-1047.00000000000,78.0000000000000,
552.000000000000,-794.000000000000,
115.000000000000,1047.00000000000,
311.000000000000,-60.0000000000000,
-92.0000000000000,-415.000000000000,
-206.000000000000,1204.00000000000,
21.0000000000000,232.000000000000,
-422.000000000000,874.000000000000,
582.000000000000,722.000000000000,
-116.000000000000,446.000000000000,
-313.000000000000,695.000000000000,
167.000000000000,158.000000000000,
129.000000000000,831.000000000000,
-507.000000000000,725.000000000000,
50.0000000000000,653.000000000000,
-356.000000000000,132.000000000000,
-684.000000000000,541.000000000000,
192.000000000000,-213.000000000000,
-258.000000000000,-1265.00000000000,
1065.00000000000,-937.000000000000,
-85.0000000000000,-1053.00000000000,
27.0000000000000,17.0000000000000,
700.000000000000,-1337.00000000000,
-841.000000000000,731.000000000000,
-139.000000000000,840.000000000000,
-852.000000000000,-164.000000000000,
59.0000000000000,1003.00000000000,
-318.000000000000,-1144.00000000000,
-465.000000000000,525.000000000000,
-439.000000000000,166.000000000000,
-869.000000000000,49.0000000000000,
66.0000000000000,-341.000000000000,
-611.000000000000,-931.000000000000,
313.000000000000,1301.00000000000,
265.000000000000,310.000000000000,
-421.000000000000,204.000000000000,
-403.000000000000,-994.000000000000,
720.000000000000,-755.000000000000,
1214.00000000000,-524.000000000000,
111.000000000000,-115.000000000000,
592.000000000000,1135.00000000000,
-138.000000000000,-41.0000000000000,
221.000000000000,565.000000000000,
719.000000000000,-226.000000000000,
527.000000000000,-122.000000000000,
333.000000000000,59.0000000000000,
-145.000000000000,396.000000000000,
-316.000000000000,814.000000000000,
21.0000000000000,-1292.00000000000,
343.000000000000,157.000000000000,
-654.000000000000,328.000000000000,
5.00000000000000,-1111.00000000000,
-37.0000000000000,191.000000000000,
-841.000000000000,1020.00000000000,
-504.000000000000,-761.000000000000,
-179.000000000000,-924.000000000000,
114.000000000000,780.000000000000,
-713.000000000000,-174.000000000000,
287.000000000000,147.000000000000,
984.000000000000,177.000000000000,
-430.000000000000,361.000000000000,
-243.000000000000,507.000000000000,
-145.000000000000,-1207.00000000000,
364.000000000000,-95.0000000000000,
369.000000000000,-126.000000000000,
-305.000000000000,-455.000000000000,
-258.000000000000,-717.000000000000,
-327.000000000000,-150.000000000000,
-336.000000000000,312.000000000000,
60.0000000000000,-878.000000000000,
51.0000000000000,-236.000000000000,
-450.000000000000,591.000000000000,
129.000000000000,1314.00000000000,
-881.000000000000,-335.000000000000,
-306.000000000000,-602.000000000000,
1591.00000000000,931.000000000000,
404.000000000000,572.000000000000,
177.000000000000,678.000000000000,
94.0000000000000,224.000000000000,
-915.000000000000,111.000000000000,
-672.000000000000,452.000000000000,
53.0000000000000,446.000000000000,
259.000000000000,566.000000000000,
-1046.00000000000,91.0000000000000,
-64.0000000000000,-658.000000000000,
688.000000000000,-363.000000000000,
347.000000000000,291.000000000000,
1196.00000000000,26.0000000000000,
84.0000000000000,348.000000000000,
41.0000000000000,-833.000000000000,
179.000000000000,-121.000000000000,
378.000000000000,489.000000000000,
-24.0000000000000,-679.000000000000,
721.000000000000,1014.00000000000,
351.000000000000,-74.0000000000000,
-1367.00000000000,-119.000000000000,
147.000000000000,-39.0000000000000,
-925.000000000000,135.000000000000,
-314.000000000000,1094.00000000000,
258.000000000000,-1267.00000000000,
396.000000000000,-654.000000000000,
858.000000000000,33.0000000000000,
-75.0000000000000,766.000000000000,
261.000000000000,902.000000000000,
-989.000000000000,61.0000000000000,
-277.000000000000,-298.000000000000,
-75.0000000000000,-591.000000000000,
-259.000000000000,651.000000000000,
-129.000000000000,-688.000000000000,
-978.000000000000,-676.000000000000,
164.000000000000,368.000000000000,
93.0000000000000,258.000000000000,
411.000000000000,-932.000000000000,
729.000000000000,-1105.00000000000,
35.0000000000000,836.000000000000,
-115.000000000000,36.0000000000000,
701.000000000000,376.000000000000,
-8.00000000000000,658.000000000000,
-986.000000000000,-308.000000000000,
171.000000000000,328.000000000000,
406.000000000000,249.000000000000,
-285.000000000000,800.000000000000,
-617.000000000000,762.000000000000,
-340.000000000000,872.000000000000,
-560.000000000000,590.000000000000,
159.000000000000,-239.000000000000,
992.000000000000,-92.0000000000000,
-327.000000000000,683.000000000000,
390.000000000000,1050.00000000000,
-346.000000000000,-114.000000000000,
-735.000000000000,619.000000000000,
31.0000000000000,-942.000000000000,
-1147.00000000000,-302.000000000000,
536.000000000000,484.000000000000,
91.0000000000000,-1268.00000000000,
-716.000000000000,1271.00000000000,
-396.000000000000,152.000000000000,
-992.000000000000,-294.000000000000,
-209.000000000000,-5.00000000000000,
179.000000000000,-1181.00000000000,
721.000000000000,-54.0000000000000,
644.000000000000,672.000000000000,
789.000000000000,-600.000000000000,
194.000000000000,-1041.00000000000,
85.0000000000000,426.000000000000,
198.000000000000,-517.000000000000,
331.000000000000,-128.000000000000,
496.000000000000,1169.00000000000,
-1035.00000000000,654.000000000000,
115.000000000000,178.000000000000,
662.000000000000,347.000000000000,
-606.000000000000,1599.00000000000,
-747.000000000000,-404.000000000000,
-863.000000000000,-892.000000000000,
757.000000000000,289.000000000000,
-458.000000000000,188.000000000000,
-713.000000000000,444.000000000000,
346.000000000000,-163.000000000000,
-46.0000000000000,-282.000000000000,
-231.000000000000,-711.000000000000,
-1075.00000000000,-608.000000000000,
-173.000000000000,-1240.00000000000,
-599.000000000000,-404.000000000000,
191.000000000000,344.000000000000,
-135.000000000000,-637.000000000000,
-620.000000000000,228.000000000000,
821.000000000000,-192.000000000000,
77.0000000000000,-355.000000000000,
581.000000000000,21.0000000000000,
131.000000000000,-109.000000000000,
348.000000000000,-779.000000000000,
24.0000000000000,-689.000000000000,
-289.000000000000,-302.000000000000,
991.000000000000,81.0000000000000,
-617.000000000000,1448.00000000000,
-674.000000000000,1129.00000000000,
-551.000000000000,-16.0000000000000,
70.0000000000000,-305.000000000000,
275.000000000000,640.000000000000,
-684.000000000000,-519.000000000000,
-394.000000000000,-78.0000000000000,
-765.000000000000,766.000000000000,
-184.000000000000,-927.000000000000,
212.000000000000,-342.000000000000,
774.000000000000,491.000000000000,
279.000000000000,666.000000000000,
-855.000000000000,231.000000000000,
-26.0000000000000,-667.000000000000,
408.000000000000,-693.000000000000,
110.000000000000,-1002.00000000000,
-532.000000000000,69.0000000000000,
-261.000000000000,84.0000000000000,
-412.000000000000,-710.000000000000,
151.000000000000,780.000000000000,
-453.000000000000,-447.000000000000,
17.0000000000000,-726.000000000000,
1057.00000000000,-999.000000000000,
-769.000000000000,-165.000000000000,
178.000000000000,431.000000000000,
-416.000000000000,-1061.00000000000,
278.000000000000,802.000000000000,
1072.00000000000,-898.000000000000,
463.000000000000,-593.000000000000,
1510.00000000000,-109.000000000000,
-353.000000000000,-544.000000000000,
-731.000000000000,276.000000000000,
-503.000000000000,-1426.00000000000,
504.000000000000,-525.000000000000,
807.000000000000,561.000000000000,
-404.000000000000,-19.0000000000000,
-226.000000000000,16.0000000000000,
-486.000000000000,1191.00000000000,
602.000000000000,-475.000000000000,
-510.000000000000,-609.000000000000,
368.000000000000,903.000000000000,
1110.00000000000,-193.000000000000,
-613.000000000000,27.0000000000000,
-122.000000000000,544.000000000000,
-1122.00000000000,243.000000000000,
-470.000000000000,-1112.00000000000,
434.000000000000,230.000000000000,
648.000000000000,906.000000000000,
243.000000000000,-776.000000000000,
472.000000000000,467.000000000000,
1105.00000000000,268.000000000000,
-901.000000000000,623.000000000000,
-631.000000000000,45.0000000000000,
-837.000000000000,-1219.00000000000,
-907.000000000000,568.000000000000,
-310.000000000000,125.000000000000,
-459.000000000000,254.000000000000,
-661.000000000000,-141.000000000000,
-281.000000000000,-648.000000000000,
53.0000000000000,-316.000000000000,
-955.000000000000,-626.000000000000,
411.000000000000,-158.000000000000,
1149.00000000000,-296.000000000000,
426.000000000000,700.000000000000,
-368.000000000000,926.000000000000,
-801.000000000000,477.000000000000,
-616.000000000000,-423.000000000000,
-243.000000000000,46.0000000000000,
-77.0000000000000,337.000000000000,
9.00000000000000,-1294.00000000000,
1145.00000000000,368.000000000000,
671.000000000000,359.000000000000,
141.000000000000,286.000000000000,
-26.0000000000000,504.000000000000,
366.000000000000,-1406.00000000000,
255.000000000000,-90.0000000000000,
519.000000000000,602.000000000000,
318.000000000000,436.000000000000,
-1239.00000000000,-325.000000000000,
-211.000000000000,-766.000000000000,
-60.0000000000000,355.000000000000,
565.000000000000,-380.000000000000,
-152.000000000000,-134.000000000000,
22.0000000000000,632.000000000000,
710.000000000000,789.000000000000,
-1477.00000000000,326.000000000000,
-389.000000000000,52.0000000000000,
42.0000000000000,492.000000000000,
-901.000000000000,443.000000000000,
240.000000000000,343.000000000000,
420.000000000000,428.000000000000,
-736.000000000000,892.000000000000,
-774.000000000000,-526.000000000000,
775.000000000000,-562.000000000000,
1157.00000000000,-146.000000000000,
470.000000000000,-262.000000000000,
663.000000000000,-554.000000000000,
134.000000000000,-848.000000000000,
587.000000000000,744.000000000000,
-134.000000000000,-235.000000000000,
-839.000000000000,-898.000000000000,
918.000000000000,-246.000000000000,
-57.0000000000000,1047.00000000000,
527.000000000000,1013.00000000000,
-131.000000000000,-479.000000000000,
297.000000000000,-49.0000000000000,
669.000000000000,68.0000000000000,
-929.000000000000,1048.00000000000,
1072.00000000000,12.0000000000000,
8.00000000000000,407.000000000000,
4.00000000000000,428.000000000000,
519.000000000000,-841.000000000000,
200.000000000000,112.000000000000,
814.000000000000,-1061.00000000000,
330.000000000000,-866.000000000000,
-371.000000000000,791.000000000000,
-409.000000000000,523.000000000000,
441.000000000000,-126.000000000000,
-1045.00000000000,380.000000000000,
-349.000000000000,-392.000000000000,
948.000000000000,-844.000000000000,
298.000000000000,-434.000000000000,
966.000000000000,-288.000000000000,
686.000000000000,219.000000000000,
681.000000000000,-657.000000000000,
638.000000000000,-418.000000000000,
293.000000000000,-249.000000000000,
-41.0000000000000,-1044.00000000000,
-312.000000000000,888.000000000000,
25.0000000000000,890.000000000000,
159.000000000000,94.0000000000000,
-35.0000000000000,-629.000000000000,
-525.000000000000,-404.000000000000,
-110.000000000000,1179.00000000000,
-539.000000000000,-354.000000000000,
-735.000000000000,1008.00000000000,
-669.000000000000,-153.000000000000,
354.000000000000,-984.000000000000,
-115.000000000000,147.000000000000,
-697.000000000000,-1208.00000000000,
1231.00000000000,6.00000000000000,
130.000000000000,85.0000000000000,
-99.0000000000000,362.000000000000,
168.000000000000,-480.000000000000,
-592.000000000000,-329.000000000000,
93.0000000000000,557.000000000000,
504.000000000000,-414.000000000000,
-301.000000000000,550.000000000000,
135.000000000000,424.000000000000,
458.000000000000,-16.0000000000000,
-1106.00000000000,232.000000000000,
-776.000000000000,-112.000000000000,
362.000000000000,-1250.00000000000,
821.000000000000,-580.000000000000,
146.000000000000,867.000000000000,
-481.000000000000,-136.000000000000,
395.000000000000,-545.000000000000,
742.000000000000,-641.000000000000,
883.000000000000,100.000000000000,
751.000000000000,1100.00000000000,
51.0000000000000,641.000000000000,
-677.000000000000,253.000000000000,
-1157.00000000000,-201.000000000000,
-1016.00000000000,326.000000000000,
-124.000000000000,190.000000000000,
673.000000000000,-153.000000000000,
-346.000000000000,43.0000000000000,
-155.000000000000,600.000000000000,
-104.000000000000,362.000000000000,
-350.000000000000,-1147.00000000000,
-205.000000000000,-720.000000000000,
-515.000000000000,-440.000000000000,
-198.000000000000,-783.000000000000,
-218.000000000000,-369.000000000000,
-533.000000000000,-468.000000000000,
-234.000000000000,-178.000000000000,
-482.000000000000,515.000000000000,
821.000000000000,795.000000000000,
801.000000000000,644.000000000000,
-1015.00000000000,788.000000000000,
-32.0000000000000,-57.0000000000000,
378.000000000000,84.0000000000000,
1021.00000000000,441.000000000000,
-794.000000000000,605.000000000000,
-334.000000000000,127.000000000000,
758.000000000000,-382.000000000000,
-718.000000000000,633.000000000000,
346.000000000000,398.000000000000,
-1282.00000000000,508.000000000000,
-148.000000000000,-671.000000000000,
-7.00000000000000,-695.000000000000,
-252.000000000000,-329.000000000000,
824.000000000000,-1254.00000000000,
-324.000000000000,254.000000000000,
449.000000000000,717.000000000000,
-78.0000000000000,775.000000000000,
101.000000000000,-96.0000000000000,
343.000000000000,-1124.00000000000,
-451.000000000000,699.000000000000,
-248.000000000000,190.000000000000,
467.000000000000,-258.000000000000,
627.000000000000,403.000000000000,
688.000000000000,1041.00000000000,
-83.0000000000000,463.000000000000,
-52.0000000000000,-867.000000000000,
852.000000000000,-481.000000000000,
-829.000000000000,-763.000000000000,
276.000000000000,-678.000000000000,
891.000000000000,-1155.00000000000,
-763.000000000000,552.000000000000,
-262.000000000000,779.000000000000,
-692.000000000000,-921.000000000000,
-318.000000000000,1198.00000000000,
102.000000000000,563.000000000000,
-442.000000000000,-588.000000000000,
-588.000000000000,260.000000000000,
-968.000000000000,123.000000000000,
-521.000000000000,-1091.00000000000,
224.000000000000,-437.000000000000,
737.000000000000,95.0000000000000,
-190.000000000000,-922.000000000000,
-352.000000000000,-483.000000000000,
521.000000000000,158.000000000000,
627.000000000000,843.000000000000,
665.000000000000,769.000000000000,
-723.000000000000,385.000000000000,
849.000000000000,83.0000000000000,
-111.000000000000,405.000000000000,
-741.000000000000,-74.0000000000000,
865.000000000000,-1255.00000000000,
-874.000000000000,803.000000000000,
343.000000000000,228.000000000000,
-686.000000000000,-1076.00000000000,
738.000000000000,-584.000000000000,
566.000000000000,242.000000000000,
-678.000000000000,554.000000000000,
931.000000000000,-357.000000000000,
-1155.00000000000,876.000000000000,
-559.000000000000,-460.000000000000,
-602.000000000000,-316.000000000000,
616.000000000000,841.000000000000,
-289.000000000000,337.000000000000,
-319.000000000000,17.0000000000000,
722.000000000000,-976.000000000000,
-882.000000000000,-288.000000000000,
970.000000000000,-684.000000000000,
222.000000000000,-1056.00000000000,
707.000000000000,-107.000000000000,
1282.00000000000,160.000000000000,
-247.000000000000,-165.000000000000,
182.000000000000,-218.000000000000,
-430.000000000000,26.0000000000000,
-747.000000000000,-781.000000000000,
226.000000000000,-709.000000000000,
1109.00000000000,-482.000000000000,
551.000000000000,-2.00000000000000,
204.000000000000,196.000000000000,
-213.000000000000,-760.000000000000,
-201.000000000000,-672.000000000000,
41.0000000000000,-672.000000000000,
1.00000000000000,-658.000000000000,
69.0000000000000,-104.000000000000,
-914.000000000000,35.0000000000000,
144.000000000000,-55.0000000000000,
48.0000000000000,-249.000000000000,
13.0000000000000,-409.000000000000,
1324.00000000000,-653.000000000000,
-631.000000000000,646.000000000000,
-558.000000000000,201.000000000000,
-881.000000000000,-324.000000000000,
-594.000000000000,519.000000000000,
8.00000000000000,138.000000000000,
-758.000000000000,443.000000000000,
787.000000000000,-661.000000000000,
866.000000000000,-430.000000000000,
330.000000000000,-52.0000000000000,
-233.000000000000,-798.000000000000,
393.000000000000,-32.0000000000000,
-489.000000000000,-729.000000000000,
-861.000000000000,-402.000000000000,
767.000000000000,-518.000000000000,
116.000000000000,702.000000000000,
-474.000000000000,1247.00000000000,
-340.000000000000,-389.000000000000,
443.000000000000,-328.000000000000,
172.000000000000,-319.000000000000,
148.000000000000,582.000000000000,
-556.000000000000,672.000000000000,
-1346.00000000000,-156.000000000000,
651.000000000000,-923.000000000000,
1163.00000000000,-1176.00000000000,
85.0000000000000,-360.000000000000,
-38.0000000000000,28.0000000000000,
-91.0000000000000,370.000000000000,
-1.00000000000000,152.000000000000,
123.000000000000,331.000000000000,
-647.000000000000,-226.000000000000,
373.000000000000,-241.000000000000,
970.000000000000,226.000000000000,
-245.000000000000,-444.000000000000,
586.000000000000,780.000000000000,
19.0000000000000,-174.000000000000,
-441.000000000000,89.0000000000000,
582.000000000000,594.000000000000,
-842.000000000000,-894.000000000000,
-636.000000000000,-353.000000000000,
-5.00000000000000,-433.000000000000,
-25.0000000000000,-639.000000000000,
-68.0000000000000,-664.000000000000,
-182.000000000000,-820.000000000000,
918.000000000000,430.000000000000,
227.000000000000,625.000000000000,
-469.000000000000,-495.000000000000,
335.000000000000,358.000000000000,
223.000000000000,465.000000000000,
-2.00000000000000,304.000000000000,
362.000000000000,1262.00000000000,
238.000000000000,235.000000000000,
282.000000000000,391.000000000000,
841.000000000000,666.000000000000,
-95.0000000000000,-773.000000000000,
-474.000000000000,-435.000000000000,
78.0000000000000,182.000000000000,
-200.000000000000,1221.00000000000,
-942.000000000000,127.000000000000,
-1206.00000000000,-1029.00000000000,
-407.000000000000,17.0000000000000,
-16.0000000000000,-596.000000000000,
610.000000000000,658.000000000000,
363.000000000000,760.000000000000,
-161.000000000000,537.000000000000,
418.000000000000,92.0000000000000,
716.000000000000,572.000000000000,
-423.000000000000,1010.00000000000,
-776.000000000000,-391.000000000000,
343.000000000000,651.000000000000,
-732.000000000000,-635.000000000000,
-248.000000000000,-245.000000000000,
759.000000000000,659.000000000000,
91.0000000000000,503.000000000000,
919.000000000000,188.000000000000,
210.000000000000,-63.0000000000000,
226.000000000000,1150.00000000000,
114.000000000000,-5.00000000000000,
-387.000000000000,456.000000000000,
-49.0000000000000,952.000000000000,
-1065.00000000000,277.000000000000,
-305.000000000000,-124.000000000000,
195.000000000000,-446.000000000000,
137.000000000000,66.0000000000000,
-680.000000000000,-483.000000000000,
-835.000000000000,0.00000000000000,
478.000000000000,214.000000000000,
-601.000000000000,-130.000000000000,
555.000000000000,-211.000000000000,
967.000000000000,686.000000000000,
755.000000000000,413.000000000000,
384.000000000000,-95.0000000000000,
-286.000000000000,1086.00000000000,
-211.000000000000,-606.000000000000,
-559.000000000000,-808.000000000000,
635.000000000000,290.000000000000,
-625.000000000000,781.000000000000,
-510.000000000000,580.000000000000,
-469.000000000000,-815.000000000000,
-1009.00000000000,45.0000000000000,
387.000000000000,-339.000000000000,
147.000000000000,-29.0000000000000,
16.0000000000000,1020.00000000000,
-590.000000000000,-92.0000000000000,
-699.000000000000,-592.000000000000,
-107.000000000000,-147.000000000000,
31.0000000000000,712.000000000000,
-175.000000000000,730.000000000000,
303.000000000000,312.000000000000,
958.000000000000,-812.000000000000,
-154.000000000000,-544.000000000000,
554.000000000000,63.0000000000000,
1099.00000000000,87.0000000000000,
240.000000000000,1283.00000000000,
-655.000000000000,-377.000000000000,
-504.000000000000,-554.000000000000,
208.000000000000,174.000000000000,
-1074.00000000000,129.000000000000,
-301.000000000000,449.000000000000,
-328.000000000000,-36.0000000000000,
649.000000000000,729.000000000000,
544.000000000000,-256.000000000000,
-1233.00000000000,-16.0000000000000,
488.000000000000,-308.000000000000,
-810.000000000000,-336.000000000000,
211.000000000000,-524.000000000000,
1113.00000000000,-1126.00000000000,
363.000000000000,875.000000000000,
-126.000000000000,-735.000000000000,
-566.000000000000,-303.000000000000,
829.000000000000,-810.000000000000,
178.000000000000,-524.000000000000,
1303.00000000000,1292.00000000000,
63.0000000000000,-83.0000000000000,
-125.000000000000,714.000000000000,
-60.0000000000000,-680.000000000000,
-541.000000000000,306.000000000000,
987.000000000000,226.000000000000,
-1009.00000000000,-694.000000000000,
831.000000000000,-107.000000000000,
706.000000000000,-145.000000000000,
130.000000000000,997.000000000000,
125.000000000000,-732.000000000000,
-1194.00000000000,423.000000000000,
199.000000000000,190.000000000000,
-329.000000000000,-350.000000000000,
794.000000000000,-248.000000000000,
213.000000000000,-214.000000000000,
-7.00000000000000,1190.00000000000,
28.0000000000000,-966.000000000000,
-300.000000000000,-701.000000000000,
450.000000000000,-977.000000000000,
-859.000000000000,-256.000000000000,
42.0000000000000,-234.000000000000,
487.000000000000,-1112.00000000000,
1354.00000000000,1091.00000000000,
537.000000000000,-671.000000000000,
-134.000000000000,292.000000000000,
-86.0000000000000,503.000000000000,
-1219.00000000000,-719.000000000000,
899.000000000000,-644.000000000000,
-552.000000000000,-962.000000000000,
214.000000000000,185.000000000000,
563.000000000000,544.000000000000,
-737.000000000000,463.000000000000,
649.000000000000,-996.000000000000,
-673.000000000000,-289.000000000000,
110.000000000000,-817.000000000000,
372.000000000000,-831.000000000000,
1199.00000000000,622.000000000000,
217.000000000000,170.000000000000,
-1262.00000000000,906.000000000000,
231.000000000000,-942.000000000000,
-63.0000000000000,-788.000000000000,
-23.0000000000000,368.000000000000,
-779.000000000000,104.000000000000,
-379.000000000000,152.000000000000,
-210.000000000000,-718.000000000000,
740.000000000000,604.000000000000,
503.000000000000,-209.000000000000,
-605.000000000000,150.000000000000,
1058.00000000000,677.000000000000,
-793.000000000000,-162.000000000000,
-336.000000000000,-731.000000000000,
112.000000000000,-1450.00000000000,
111.000000000000,816.000000000000,
422.000000000000,774.000000000000,
-820.000000000000,339.000000000000,
1120.00000000000,93.0000000000000,
-226.000000000000,808.000000000000,
-511.000000000000,1168.00000000000,
-756.000000000000,-645.000000000000,
-566.000000000000,-180.000000000000,
1186.00000000000,-44.0000000000000,
187.000000000000,1033.00000000000,
637.000000000000,451.000000000000,
580.000000000000,-254.000000000000,
866.000000000000,-372.000000000000,
599.000000000000,-556.000000000000,
582.000000000000,1060.00000000000,
72.0000000000000,-808.000000000000,
-739.000000000000,64.0000000000000,
-251.000000000000,394.000000000000,
-495.000000000000,-311.000000000000,
374.000000000000,1373.00000000000,
-340.000000000000,650.000000000000,
-380.000000000000,950.000000000000,
-1134.00000000000,-49.0000000000000,
-831.000000000000,146.000000000000,
1120.00000000000,262.000000000000,
-251.000000000000,450.000000000000,
529.000000000000,132.000000000000,
157.000000000000,-176.000000000000,
-400.000000000000,1396.00000000000,
608.000000000000,-1220.00000000000,
352.000000000000,34.0000000000000,
196.000000000000,648.000000000000,
348.000000000000,-763.000000000000,
127.000000000000,-157.000000000000,
-637.000000000000,-994.000000000000,
120.000000000000,-410.000000000000,
281.000000000000,-219.000000000000,
-17.0000000000000,832.000000000000,
-697.000000000000,-105.000000000000,
-438.000000000000,-940.000000000000,
630.000000000000,820.000000000000,
-1251.00000000000,767.000000000000,
-308.000000000000,-165.000000000000,
-299.000000000000,-78.0000000000000,
-745.000000000000,327.000000000000,
1109.00000000000,-149.000000000000,
-588.000000000000,1061.00000000000,
886.000000000000,-189.000000000000,
-414.000000000000,-385.000000000000,
-98.0000000000000,970.000000000000,
854.000000000000,-96.0000000000000,
-1402.00000000000,719.000000000000,
246.000000000000,-120.000000000000,
155.000000000000,31.0000000000000,
742.000000000000,1017.00000000000,
305.000000000000,596.000000000000,
-34.0000000000000,-40.0000000000000,
-206.000000000000,-1121.00000000000,
-863.000000000000,-745.000000000000,
137.000000000000,-724.000000000000,
440.000000000000,735.000000000000,
391.000000000000,737.000000000000,
-537.000000000000,889.000000000000,
-7.00000000000000,1061.00000000000,
-670.000000000000,-1151.00000000000,
-786.000000000000,643.000000000000,
-451.000000000000,62.0000000000000,
72.0000000000000,-776.000000000000,
1295.00000000000,172.000000000000,
-758.000000000000,697.000000000000,
484.000000000000,892.000000000000,
-102.000000000000,-874.000000000000,
-884.000000000000,441.000000000000,
723.000000000000,381.000000000000,
-937.000000000000,587.000000000000,
179.000000000000,190.000000000000,
161.000000000000,160.000000000000,
-1055.00000000000,1090.00000000000,
24.0000000000000,207.000000000000,
613.000000000000,1149.00000000000,
-714.000000000000,-443.000000000000,
-1046.00000000000,205.000000000000,
-728.000000000000,675.000000000000,
-567.000000000000,-706.000000000000,
-134.000000000000,412.000000000000,
-517.000000000000,-619.000000000000,
368.000000000000,-875.000000000000,
120.000000000000,-569.000000000000,
-474.000000000000,74.0000000000000,
-401.000000000000,933.000000000000,
101.000000000000,-283.000000000000,
897.000000000000,-597.000000000000,
839.000000000000,450.000000000000,
234.000000000000,137.000000000000,
-747.000000000000,563.000000000000,
-879.000000000000,583.000000000000,
152.000000000000,-189.000000000000,
-107.000000000000,825.000000000000,
-522.000000000000,475.000000000000,
-1539.00000000000,-52.0000000000000,
43.0000000000000,273.000000000000,
688.000000000000,116.000000000000,
-1261.00000000000,747.000000000000,
441.000000000000,-1110.00000000000,
608.000000000000,-822.000000000000,
384.000000000000,876.000000000000,
258.000000000000,372.000000000000,
48.0000000000000,1115.00000000000,
120.000000000000,117.000000000000,
-399.000000000000,-945.000000000000,
-565.000000000000,-299.000000000000,
-1136.00000000000,-823.000000000000,
641.000000000000,-736.000000000000,
1029.00000000000,725.000000000000,
428.000000000000,130.000000000000,
439.000000000000,32.0000000000000,
186.000000000000,-358.000000000000,
672.000000000000,-401.000000000000,
192.000000000000,375.000000000000,
573.000000000000,-60.0000000000000,
-311.000000000000,675.000000000000,
-865.000000000000,-115.000000000000,
-225.000000000000,-907.000000000000,
-764.000000000000,-125.000000000000,
32.0000000000000,-1053.00000000000,
104.000000000000,-654.000000000000,
-347.000000000000,343.000000000000,
-841.000000000000,-234.000000000000,
132.000000000000,-633.000000000000,
791.000000000000,-1052.00000000000,
-49.0000000000000,-159.000000000000,
-394.000000000000,540.000000000000,
-351.000000000000,-416.000000000000,
199.000000000000,81.0000000000000,
173.000000000000,661.000000000000,
59.0000000000000,-780.000000000000,
-396.000000000000,-911.000000000000,
-359.000000000000,865.000000000000,
528.000000000000,365.000000000000,
390.000000000000,398.000000000000,
65.0000000000000,974.000000000000,
372.000000000000,317.000000000000,
355.000000000000,582.000000000000,
-608.000000000000,740.000000000000,
-776.000000000000,397.000000000000,
-990.000000000000,-929.000000000000,
-611.000000000000,220.000000000000,
693.000000000000,75.0000000000000,
-292.000000000000,-942.000000000000,
-59.0000000000000,160.000000000000,
-14.0000000000000,-1019.00000000000,
87.0000000000000,706.000000000000,
1008.00000000000,991.000000000000,
33.0000000000000,-27.0000000000000,
-303.000000000000,-513.000000000000,
-154.000000000000,-492.000000000000,
-343.000000000000,363.000000000000,
-697.000000000000,-297.000000000000,
173.000000000000,5.00000000000000,
466.000000000000,-874.000000000000,
270.000000000000,-216.000000000000,
-126.000000000000,-15.0000000000000,
-1077.00000000000,-1266.00000000000,
420.000000000000,-667.000000000000,
-89.0000000000000,-549.000000000000,
-313.000000000000,-598.000000000000,
1329.00000000000,-1137.00000000000,
937.000000000000,888.000000000000,
345.000000000000,613.000000000000,
-533.000000000000,-128.000000000000,
-412.000000000000,943.000000000000,
-542.000000000000,-440.000000000000,
184.000000000000,-34.0000000000000,
-8.00000000000000,-422.000000000000,
-185.000000000000,-553.000000000000,
1301.00000000000,-899.000000000000,
-363.000000000000,289.000000000000,
-957.000000000000,310.000000000000,
-146.000000000000,-1319.00000000000,
934.000000000000,1064.00000000000,
-92.0000000000000,601.000000000000,
-513.000000000000,-797.000000000000,
1321.00000000000,-539.000000000000,
-12.0000000000000,-468.000000000000,
570.000000000000,-560.000000000000,
1281.00000000000,-368.000000000000,
-254.000000000000,558.000000000000,
-592.000000000000,567.000000000000,
176.000000000000,-427.000000000000,
822.000000000000,-291.000000000000,
717.000000000000,252.000000000000,
1336.00000000000,235.000000000000,
-285.000000000000,1068.00000000000,
-200.000000000000,-373.000000000000,
389.000000000000,-735.000000000000,
-1270.00000000000,1241.00000000000,
-253.000000000000,-78.0000000000000,
699.000000000000,597.000000000000,
551.000000000000,833.000000000000,
231.000000000000,-677.000000000000,
568.000000000000,895.000000000000,
-672.000000000000,301.000000000000,
-1026.00000000000,-72.0000000000000,
136.000000000000,-891.000000000000,
-325.000000000000,-247.000000000000,
-21.0000000000000,1039.00000000000,
-1405.00000000000,-953.000000000000,
470.000000000000,-805.000000000000,
888.000000000000,340.000000000000,
-905.000000000000,402.000000000000,
915.000000000000,-476.000000000000,
130.000000000000,-687.000000000000,
-283.000000000000,-224.000000000000,
-50.0000000000000,279.000000000000,
567.000000000000,-391.000000000000,
767.000000000000,-263.000000000000,
1144.00000000000,983.000000000000,
632.000000000000,595.000000000000,
-1428.00000000000,448.000000000000,
-7.00000000000000,295.000000000000,
-441.000000000000,591.000000000000,
-5.00000000000000,-151.000000000000,
337.000000000000,-765.000000000000,
-217.000000000000,341.000000000000,
908.000000000000,-136.000000000000,
236.000000000000,278.000000000000,
763.000000000000,1188.00000000000,
513.000000000000,366.000000000000,
369.000000000000,329.000000000000,
259.000000000000,779.000000000000,
-130.000000000000,150.000000000000,
629.000000000000,-875.000000000000,
497.000000000000,-35.0000000000000,
-81.0000000000000,558.000000000000,
-911.000000000000,594.000000000000,
-941.000000000000,-497.000000000000,
-377.000000000000,-611.000000000000,
1024.00000000000,989.000000000000,
-53.0000000000000,21.0000000000000,
-458.000000000000,141.000000000000,
1255.00000000000,1097.00000000000,
-1265.00000000000,525.000000000000,
117.000000000000,208.000000000000,
502.000000000000,413.000000000000,
-1363.00000000000,1094.00000000000,
-573.000000000000,446.000000000000,
-881.000000000000,-998.000000000000,
321.000000000000,-171.000000000000,
-228.000000000000,472.000000000000,
930.000000000000,-1158.00000000000,
146.000000000000,243.000000000000,
265.000000000000,994.000000000000,
558.000000000000,376.000000000000,
-1594.00000000000,-65.0000000000000,
881.000000000000,-252.000000000000,
-545.000000000000,647.000000000000,
-1174.00000000000,-383.000000000000,
-501.000000000000,-312.000000000000,
-449.000000000000,-288.000000000000,
904.000000000000,-724.000000000000,
103.000000000000,150.000000000000,
-648.000000000000,-582.000000000000,
-653.000000000000,379.000000000000,
253.000000000000,662.000000000000,
323.000000000000,-1039.00000000000,
95.0000000000000,-247.000000000000,
-143.000000000000,-482.000000000000,
749.000000000000,467.000000000000,
694.000000000000,124.000000000000,
-649.000000000000,-718.000000000000,
836.000000000000,299.000000000000,
342.000000000000,126.000000000000,
13.0000000000000,134.000000000000,
-237.000000000000,-234.000000000000,
-373.000000000000,723.000000000000,
889.000000000000,-686.000000000000,
578.000000000000,-271.000000000000,
731.000000000000,181.000000000000,
-970.000000000000,-993.000000000000,
259.000000000000,952.000000000000,
456.000000000000,644.000000000000,
-715.000000000000,-24.0000000000000,
147.000000000000,-13.0000000000000,
-1138.00000000000,639.000000000000,
550.000000000000,-54.0000000000000,
581.000000000000,-942.000000000000,
1008.00000000000,-178.000000000000,
381.000000000000,440.000000000000,
-496.000000000000,1223.00000000000,
616.000000000000,-364.000000000000,
-1291.00000000000,-77.0000000000000,
-62.0000000000000,352.000000000000,
357.000000000000,220.000000000000,
531.000000000000,184.000000000000,
610.000000000000,-1125.00000000000,
379.000000000000,286.000000000000,
200.000000000000,-745.000000000000,
-787.000000000000,-401.000000000000,
1112.00000000000,-95.0000000000000,
497.000000000000,-488.000000000000,
-365.000000000000,106.000000000000,
-341.000000000000,-870.000000000000,
-685.000000000000,1048.00000000000,
-533.000000000000,-635.000000000000,
742.000000000000,-177.000000000000,
1201.00000000000,1234.00000000000,
-754.000000000000,-174.000000000000,
-681.000000000000,-263.000000000000,
-446.000000000000,-1169.00000000000,
458.000000000000,636.000000000000,
804.000000000000,-336.000000000000,
705.000000000000,-794.000000000000,
758.000000000000,-386.000000000000,
-878.000000000000,-443.000000000000,
-349.000000000000,737.000000000000,
154.000000000000,225.000000000000,
330.000000000000,460.000000000000,
-124.000000000000,56.0000000000000,
-338.000000000000,131.000000000000,
807.000000000000,-462.000000000000,
-778.000000000000,-420.000000000000,
-239.000000000000,165.000000000000,
516.000000000000,-205.000000000000,
506.000000000000,443.000000000000,
445.000000000000,511.000000000000,
-616.000000000000,1133.00000000000,
-626.000000000000,551.000000000000,
-1166.00000000000,-350.000000000000,
508.000000000000,4.00000000000000,
-691.000000000000,-83.0000000000000,
-283.000000000000,-854.000000000000,
1376.00000000000,-378.000000000000,
137.000000000000,346.000000000000,
967.000000000000,-184.000000000000,
-219.000000000000,252.000000000000,
542.000000000000,20.0000000000000,
910.000000000000,608.000000000000,
-867.000000000000,631.000000000000,
-810.000000000000,-985.000000000000,
-623.000000000000,160.000000000000,
-579.000000000000,713.000000000000,
-559.000000000000,-594.000000000000,
290.000000000000,-273.000000000000,
1225.00000000000,746.000000000000,
-278.000000000000,704.000000000000,
-373.000000000000,72.0000000000000,
633.000000000000,537.000000000000,
-961.000000000000,-150.000000000000,
-365.000000000000,-171.000000000000,
122.000000000000,74.0000000000000,
-183.000000000000,-118.000000000000,
839.000000000000,915.000000000000,
326.000000000000,-344.000000000000,
-320.000000000000,554.000000000000,
-675.000000000000,786.000000000000,
-55.0000000000000,374.000000000000,
354.000000000000,53.0000000000000,
15.0000000000000,-849.000000000000,
-48.0000000000000,747.000000000000,
-273.000000000000,151.000000000000,
-208.000000000000,153.000000000000,
-250.000000000000,-356.000000000000,
-98.0000000000000,226.000000000000,
-571.000000000000,862.000000000000,
-944.000000000000,-696.000000000000,
-188.000000000000,188.000000000000,
-874.000000000000,58.0000000000000,
-532.000000000000,-740.000000000000,
286.000000000000,-862.000000000000,
-789.000000000000,97.0000000000000,
-626.000000000000,-392.000000000000,
-579.000000000000,-1305.00000000000,
87.0000000000000,-333.000000000000,
6.00000000000000,-142.000000000000,
148.000000000000,162.000000000000,
1137.00000000000,266.000000000000,
46.0000000000000,237.000000000000,
-78.0000000000000,-704.000000000000,
-614.000000000000,-841.000000000000,
-855.000000000000,-332.000000000000,
111.000000000000,-886.000000000000,
1051.00000000000,-591.000000000000,
97.0000000000000,-42.0000000000000,
-632.000000000000,388.000000000000,
986.000000000000,-950.000000000000,
187.000000000000,-24.0000000000000,
-18.0000000000000,859.000000000000,
510.000000000000,-768.000000000000,
-77.0000000000000,798.000000000000,
-533.000000000000,632.000000000000,
-276.000000000000,222.000000000000,
435.000000000000,-254.000000000000,
-203.000000000000,-585.000000000000,
-209.000000000000,645.000000000000,
-907.000000000000,48.0000000000000,
-53.0000000000000,-38.0000000000000,
518.000000000000,-1099.00000000000,
-604.000000000000,-69.0000000000000,
785.000000000000,484.000000000000,
729.000000000000,264.000000000000,
270.000000000000,460.000000000000,
254.000000000000,-454.000000000000,
-54.0000000000000,976.000000000000,
-323.000000000000,881.000000000000,
333.000000000000,-319.000000000000,
1097.00000000000,-938.000000000000,
609.000000000000,186.000000000000,
794.000000000000,886.000000000000,
423.000000000000,570.000000000000,
545.000000000000,1098.00000000000,
-340.000000000000,-263.000000000000,
-630.000000000000,-199.000000000000,
427.000000000000,-612.000000000000,
-673.000000000000,-526.000000000000,
195.000000000000,383.000000000000,
822.000000000000,406.000000000000,
63.0000000000000,1213.00000000000,
-608.000000000000,-560.000000000000,
-952.000000000000,-782.000000000000,
-183.000000000000,-550.000000000000,
-291.000000000000,435.000000000000,
-392.000000000000,715.000000000000,
-1179.00000000000,-1468.00000000000,
431.000000000000,-619.000000000000,
728.000000000000,549.000000000000,
-627.000000000000,331.000000000000,
140.000000000000,-977.000000000000,
67.0000000000000,-847.000000000000,
188.000000000000,-282.000000000000,
118.000000000000,-340.000000000000,
-355.000000000000,-191.000000000000,
-76.0000000000000,-832.000000000000,
976.000000000000,-190.000000000000,
765.000000000000,337.000000000000,
-783.000000000000,726.000000000000,
-614.000000000000,289.000000000000,
-266.000000000000,459.000000000000,
-387.000000000000,716.000000000000,
-648.000000000000,-1219.00000000000,
304.000000000000,-358.000000000000,
818.000000000000,-224.000000000000,
405.000000000000,-884.000000000000,
1321.00000000000,315.000000000000,
602.000000000000,884.000000000000,
-733.000000000000,785.000000000000,
-1210.00000000000,332.000000000000,
-1109.00000000000,-52.0000000000000,
83.0000000000000,-1219.00000000000,
991.000000000000,-845.000000000000,
709.000000000000,114.000000000000,
194.000000000000,793.000000000000,
224.000000000000,762.000000000000,
-504.000000000000,12.0000000000000,
-1296.00000000000,509.000000000000,
-391.000000000000,-1323.00000000000,
691.000000000000,-344.000000000000,
-398.000000000000,404.000000000000,
385.000000000000,-1046.00000000000,
102.000000000000,682.000000000000,
-1127.00000000000,519.000000000000,
-515.000000000000,-169.000000000000,
-134.000000000000,-545.000000000000,
438.000000000000,413.000000000000,
-200.000000000000,164.000000000000,
-29.0000000000000,-756.000000000000,
771.000000000000,430.000000000000,
-564.000000000000,267.000000000000,
-922.000000000000,899.000000000000,
-330.000000000000,-24.0000000000000,
738.000000000000,-3.00000000000000,
905.000000000000,925.000000000000,
-756.000000000000,642.000000000000,
385.000000000000,684.000000000000,
-376.000000000000,12.0000000000000,
-1287.00000000000,-336.000000000000,
98.0000000000000,-125.000000000000,
-595.000000000000,77.0000000000000,
-461.000000000000,-111.000000000000,
-660.000000000000,386.000000000000,
-920.000000000000,80.0000000000000,
202.000000000000,-675.000000000000,
386.000000000000,-291.000000000000,
-57.0000000000000,324.000000000000,
346.000000000000,585.000000000000,
51.0000000000000,866.000000000000,
-734.000000000000,325.000000000000,
-532.000000000000,-1083.00000000000,
523.000000000000,-910.000000000000,
551.000000000000,538.000000000000,
-114.000000000000,210.000000000000,
25.0000000000000,-215.000000000000,
501.000000000000,94.0000000000000,
555.000000000000,740.000000000000,
-642.000000000000,385.000000000000,
-709.000000000000,-724.000000000000,
932.000000000000,124.000000000000,
492.000000000000,1000.00000000000,
-1022.00000000000,503.000000000000,
-182.000000000000,-908.000000000000,
695.000000000000,-1324.00000000000,
-345.000000000000,-83.0000000000000,
333.000000000000,31.0000000000000,
676.000000000000,-516.000000000000,
-723.000000000000,-291.000000000000,
-753.000000000000,-25.0000000000000,
-827.000000000000,-378.000000000000,
-727.000000000000,-78.0000000000000,
-57.0000000000000,248.000000000000,
-106.000000000000,11.0000000000000,
389.000000000000,-649.000000000000,
226.000000000000,-885.000000000000,
-473.000000000000,622.000000000000,
-782.000000000000,-96.0000000000000,
-883.000000000000,-376.000000000000,
674.000000000000,6.00000000000000,
-206.000000000000,75.0000000000000,
-490.000000000000,660.000000000000,
-244.000000000000,-1030.00000000000,
128.000000000000,-440.000000000000,
1182.00000000000,-620.000000000000,
544.000000000000,-922.000000000000,
357.000000000000,202.000000000000,
-1213.00000000000,-250.000000000000,
421.000000000000,-697.000000000000,
765.000000000000,-388.000000000000,
-116.000000000000,281.000000000000,
886.000000000000,104.000000000000,
-898.000000000000,-347.000000000000,
-550.000000000000,-481.000000000000,
-462.000000000000,806.000000000000,
-1136.00000000000,75.0000000000000,
308.000000000000,-1126.00000000000,
177.000000000000,697.000000000000,
80.0000000000000,-721.000000000000,
918.000000000000,317.000000000000,
-217.000000000000,763.000000000000,
499.000000000000,-869.000000000000,
70.0000000000000,535.000000000000,
-372.000000000000,-578.000000000000,
851.000000000000,819.000000000000,
-306.000000000000,853.000000000000,
-427.000000000000,-364.000000000000,
49.0000000000000,-724.000000000000,
351.000000000000,-540.000000000000,
-96.0000000000000,852.000000000000,
-248.000000000000,574.000000000000,
778.000000000000,904.000000000000,
229.000000000000,-425.000000000000,
234.000000000000,-574.000000000000,
285.000000000000,-603.000000000000,
-426.000000000000,-472.000000000000,
96.0000000000000,855.000000000000,
-165.000000000000,105.000000000000,
-66.0000000000000,446.000000000000,
-291.000000000000,540.000000000000,
-570.000000000000,-151.000000000000,
931.000000000000,-764.000000000000,
-427.000000000000,-35.0000000000000,
132.000000000000,175.000000000000,
218.000000000000,-178.000000000000,
-474.000000000000,435.000000000000,
-671.000000000000,-624.000000000000,
-627.000000000000,-839.000000000000,
748.000000000000,-275.000000000000,
-615.000000000000,-461.000000000000,
262.000000000000,-71.0000000000000,
-717.000000000000,253.000000000000,
-52.0000000000000,-742.000000000000,
1182.00000000000,171.000000000000,
64.0000000000000,1572.00000000000,
644.000000000000,119.000000000000,
-1146.00000000000,-216.000000000000,
659.000000000000,-31.0000000000000,
1044.00000000000,-649.000000000000,
-718.000000000000,-518.000000000000,
815.000000000000,-87.0000000000000,
14.0000000000000,-614.000000000000,
-289.000000000000,504.000000000000,
448.000000000000,451.000000000000,
-847.000000000000,-749.000000000000,
313.000000000000,-481.000000000000,
225.000000000000,-157.000000000000,
-716.000000000000,703.000000000000,
1126.00000000000,-212.000000000000,
695.000000000000,-414.000000000000,
577.000000000000,98.0000000000000,
826.000000000000,329.000000000000,
-876.000000000000,592.000000000000,
292.000000000000,-682.000000000000,
218.000000000000,14.0000000000000,
-589.000000000000,934.000000000000,
44.0000000000000,-393.000000000000,
-1018.00000000000,-669.000000000000,
831.000000000000,703.000000000000,
348.000000000000,235.000000000000,
-64.0000000000000,-533.000000000000,
-82.0000000000000,446.000000000000,
-522.000000000000,-82.0000000000000,
800.000000000000,-795.000000000000,
-792.000000000000,-403.000000000000,
-422.000000000000,-508.000000000000,
-72.0000000000000,-160.000000000000,
851.000000000000,168.000000000000,
690.000000000000,95.0000000000000,
270.000000000000,111.000000000000,
654.000000000000,-953.000000000000,
-688.000000000000,10.0000000000000,
445.000000000000,24.0000000000000,
-49.0000000000000,-373.000000000000,
179.000000000000,272.000000000000,
447.000000000000,-686.000000000000,
808.000000000000,-338.000000000000,
796.000000000000,-1023.00000000000,
-350.000000000000,497.000000000000,
327.000000000000,843.000000000000,
-121.000000000000,19.0000000000000,
522.000000000000,971.000000000000,
569.000000000000,-329.000000000000,
-555.000000000000,-135.000000000000,
-388.000000000000,-307.000000000000,
-664.000000000000,-365.000000000000,
-553.000000000000,-150.000000000000,
568.000000000000,-385.000000000000,
978.000000000000,58.0000000000000,
960.000000000000,675.000000000000,
-29.0000000000000,1416.00000000000,
-1033.00000000000,-68.0000000000000,
-745.000000000000,282.000000000000,
-790.000000000000,-163.000000000000,
251.000000000000,-1539.00000000000,
-265.000000000000,-267.000000000000,
292.000000000000,-657.000000000000,
1022.00000000000,-558.000000000000,
-432.000000000000,799.000000000000,
368.000000000000,160.000000000000,
678.000000000000,584.000000000000,
-235.000000000000,490.000000000000,
-443.000000000000,-889.000000000000,
-187.000000000000,-673.000000000000,
1242.00000000000,-698.000000000000,
693.000000000000,610.000000000000,
-688.000000000000,319.000000000000,
-384.000000000000,-809.000000000000,
-970.000000000000,315.000000000000,
316.000000000000,37.0000000000000,
642.000000000000,-759.000000000000,
897.000000000000,-316.000000000000,
932.000000000000,455.000000000000,
-1620.00000000000,1274.00000000000,
-862.000000000000,-91.0000000000000,
465.000000000000,238.000000000000,
633.000000000000,611.000000000000,
653.000000000000,-244.000000000000,
948.000000000000,736.000000000000,
688.000000000000,-336.000000000000,
551.000000000000,1007.00000000000,
77.0000000000000,839.000000000000,
-959.000000000000,-783.000000000000,
-48.0000000000000,-6.00000000000000,
440.000000000000,-10.0000000000000,
110.000000000000,-319.000000000000,
366.000000000000,-488.000000000000,
-114.000000000000,802.000000000000,
-714.000000000000,-338.000000000000,
-367.000000000000,-344.000000000000,
-585.000000000000,1287.00000000000,
264.000000000000,316.000000000000,
-211.000000000000,650.000000000000,
-606.000000000000,520.000000000000,
788.000000000000,-843.000000000000,
379.000000000000,-111.000000000000,
56.0000000000000,1142.00000000000,
128.000000000000,437.000000000000,
-322.000000000000,-446.000000000000,
-922.000000000000,-679.000000000000,
291.000000000000,-1236.00000000000,
276.000000000000,-381.000000000000,
-443.000000000000,152.000000000000,
660.000000000000,-596.000000000000,
-361.000000000000,-713.000000000000,
-212.000000000000,-391.000000000000,
529.000000000000,-773.000000000000,
326.000000000000,-176.000000000000,
-52.0000000000000,1208.00000000000,
-649.000000000000,465.000000000000,
420.000000000000,64.0000000000000,
975.000000000000,-40.0000000000000,
343.000000000000,-920.000000000000,
-424.000000000000,80.0000000000000,
-147.000000000000,318.000000000000,
617.000000000000,-457.000000000000,
659.000000000000,475.000000000000,
85.0000000000000,1609.00000000000,
-666.000000000000,-239.000000000000,
-207.000000000000,-799.000000000000,
1085.00000000000,803.000000000000,
-303.000000000000,111.000000000000,
-982.000000000000,-476.000000000000,
-543.000000000000,-1274.00000000000,
-833.000000000000,-375.000000000000,
839.000000000000,179.000000000000,
291.000000000000,514.000000000000,
-399.000000000000,349.000000000000,
-259.000000000000,-303.000000000000,
-654.000000000000,967.000000000000,
-858.000000000000,-887.000000000000,
-92.0000000000000,5.00000000000000,
611.000000000000,1132.00000000000,
-441.000000000000,-154.000000000000,
-217.000000000000,276.000000000000,
-147.000000000000,-222.000000000000,
-131.000000000000,-721.000000000000,
763.000000000000,-543.000000000000,
372.000000000000,545.000000000000,
-231.000000000000,-91.0000000000000,
572.000000000000,-597.000000000000,
859.000000000000,-180.000000000000,
705.000000000000,-691.000000000000,
18.0000000000000,195.000000000000,
-490.000000000000,478.000000000000,
207.000000000000,86.0000000000000,
-29.0000000000000,646.000000000000,
-76.0000000000000,1032.00000000000,
663.000000000000,296.000000000000,
404.000000000000,298.000000000000,
172.000000000000,255.000000000000,
347.000000000000,-914.000000000000,
108.000000000000,82.0000000000000,
-803.000000000000,-181.000000000000,
-1143.00000000000,-925.000000000000,
-418.000000000000,-71.0000000000000,
-244.000000000000,-669.000000000000,
463.000000000000,-655.000000000000,
476.000000000000,293.000000000000,
213.000000000000,-200.000000000000,
187.000000000000,-43.0000000000000,
-1112.00000000000,1368.00000000000,
-791.000000000000,-512.000000000000,
-493.000000000000,-1000.00000000000,
-521.000000000000,446.000000000000,
643.000000000000,-1220.00000000000,
376.000000000000,-221.000000000000,
-225.000000000000,-604.000000000000,
465.000000000000,-708.000000000000,
330.000000000000,623.000000000000,
38.0000000000000,-330.000000000000,
1226.00000000000,-6.00000000000000,
164.000000000000,-644.000000000000,
21.0000000000000,-638.000000000000,
1054.00000000000,378.000000000000,
-567.000000000000,215.000000000000,
-631.000000000000,-421.000000000000,
398.000000000000,-148.000000000000,
921.000000000000,1054.00000000000,
-878.000000000000,1047.00000000000,
-739.000000000000,-292.000000000000,
1233.00000000000,167.000000000000,
-165.000000000000,500.000000000000,
32.0000000000000,-823.000000000000,
515.000000000000,332.000000000000,
538.000000000000,403.000000000000,
-257.000000000000,-870.000000000000,
-523.000000000000,91.0000000000000,
322.000000000000,-1062.00000000000,
245.000000000000,-447.000000000000,
1187.00000000000,906.000000000000,
537.000000000000,660.000000000000,
3.00000000000000,535.000000000000,
143.000000000000,-698.000000000000,
1047.00000000000,-192.000000000000,
374.000000000000,-510.000000000000,
-263.000000000000,-477.000000000000,
797.000000000000,-480.000000000000,
-984.000000000000,-839.000000000000,
582.000000000000,-136.000000000000,
494.000000000000,0.00000000000000,
-780.000000000000,238.000000000000,
-476.000000000000,78.0000000000000,
-923.000000000000,-29.0000000000000,
1201.00000000000,-914.000000000000,
706.000000000000,79.0000000000000,
436.000000000000,1103.00000000000,
892.000000000000,345.000000000000,
-110.000000000000,680.000000000000,
-308.000000000000,22.0000000000000,
829.000000000000,-512.000000000000,
584.000000000000,-726.000000000000,
-899.000000000000,-540.000000000000,
1027.00000000000,-994.000000000000,
427.000000000000,-401.000000000000,
-422.000000000000,1570.00000000000,
162.000000000000,-438.000000000000,
-392.000000000000,60.0000000000000,
-242.000000000000,346.000000000000,
-461.000000000000,-119.000000000000,
394.000000000000,1139.00000000000,
330.000000000000,350.000000000000,
874.000000000000,-221.000000000000,
-118.000000000000,-90.0000000000000,
-628.000000000000,241.000000000000,
1189.00000000000,-6.00000000000000,
-335.000000000000,1281.00000000000,
-102.000000000000,683.000000000000,
526.000000000000,-996.000000000000,
-599.000000000000,-263.000000000000,
253.000000000000,-991.000000000000,
590.000000000000,391.000000000000,
-993.000000000000,772.000000000000,
-287.000000000000,380.000000000000,
834.000000000000,1213.00000000000,
-1028.00000000000,663.000000000000,
-1246.00000000000,-72.0000000000000,
90.0000000000000,56.0000000000000,
397.000000000000,1275.00000000000,
324.000000000000,-209.000000000000,
533.000000000000,46.0000000000000,
-164.000000000000,636.000000000000,
-607.000000000000,-1199.00000000000,
972.000000000000,-492.000000000000,
216.000000000000,294.000000000000,
-1024.00000000000,892.000000000000,
-383.000000000000,638.000000000000,
-921.000000000000,-550.000000000000,
64.0000000000000,-484.000000000000,
1102.00000000000,603.000000000000,
-535.000000000000,32.0000000000000,
201.000000000000,-902.000000000000,
1137.00000000000,-621.000000000000,
-362.000000000000,-138.000000000000,
-484.000000000000,459.000000000000,
-865.000000000000,619.000000000000,
-586.000000000000,520.000000000000,
531.000000000000,554.000000000000,
434.000000000000,548.000000000000,
774.000000000000,-142.000000000000,
194.000000000000,-493.000000000000,
-901.000000000000,213.000000000000,
-546.000000000000,136.000000000000,
-692.000000000000,286.000000000000,
-463.000000000000,217.000000000000,
309.000000000000,-511.000000000000,
-159.000000000000,266.000000000000,
-559.000000000000,-806.000000000000,
18.0000000000000,-1521.00000000000,
888.000000000000,195.000000000000,
-79.0000000000000,622.000000000000,
-328.000000000000,-109.000000000000,
-70.0000000000000,-41.0000000000000,
-964.000000000000,1233.00000000000,
-292.000000000000,464.000000000000,
196.000000000000,-138.000000000000,
-341.000000000000,-1170.00000000000,
916.000000000000,-690.000000000000,
1135.00000000000,360.000000000000,
364.000000000000,-318.000000000000,
897.000000000000,808.000000000000,
-568.000000000000,778.000000000000,
-1266.00000000000,144.000000000000,
-47.0000000000000,-288.000000000000,
-403.000000000000,-1106.00000000000,
-27.0000000000000,-191.000000000000,
-132.000000000000,86.0000000000000,
263.000000000000,30.0000000000000,
-339.000000000000,397.000000000000,
-632.000000000000,379.000000000000,
890.000000000000,427.000000000000,
-1100.00000000000,383.000000000000,
1031.00000000000,-1189.00000000000,
429.000000000000,-750.000000000000,
3.00000000000000,533.000000000000,
1159.00000000000,-1008.00000000000,
-315.000000000000,-706.000000000000,
822.000000000000,-411.000000000000,
51.0000000000000,593.000000000000,
542.000000000000,563.000000000000,
-805.000000000000,-280.000000000000,
-312.000000000000,604.000000000000,
25.0000000000000,-1012.00000000000,
-661.000000000000,-190.000000000000,
1024.00000000000,-461.000000000000,
-908.000000000000,-914.000000000000,
325.000000000000,-586.000000000000,
433.000000000000,-942.000000000000,
-344.000000000000,530.000000000000,
-355.000000000000,53.0000000000000,
-555.000000000000,327.000000000000,
454.000000000000,116.000000000000,
-79.0000000000000,-621.000000000000,
-205.000000000000,-111.000000000000,
-1035.00000000000,439.000000000000,
-431.000000000000,161.000000000000,
904.000000000000,-1177.00000000000,
611.000000000000,78.0000000000000,
-482.000000000000,689.000000000000,
-483.000000000000,306.000000000000,
706.000000000000,-890.000000000000,
-384.000000000000,-587.000000000000,
645.000000000000,760.000000000000,
563.000000000000,-517.000000000000,
-80.0000000000000,-154.000000000000,
415.000000000000,305.000000000000,
-298.000000000000,441.000000000000,
698.000000000000,432.000000000000,
3.00000000000000,72.0000000000000,
697.000000000000,-20.0000000000000,
872.000000000000,149.000000000000,
35.0000000000000,1234.00000000000,
-367.000000000000,-362.000000000000,
-1076.00000000000,-139.000000000000,
830.000000000000,-166.000000000000,
-138.000000000000,-915.000000000000,
-200.000000000000,432.000000000000,
-290.000000000000,-61.0000000000000,
-1373.00000000000,306.000000000000,
-153.000000000000,-204.000000000000,
245.000000000000,-1040.00000000000,
493.000000000000,69.0000000000000,
429.000000000000,923.000000000000,
-243.000000000000,497.000000000000,
-1196.00000000000,63.0000000000000,
570.000000000000,531.000000000000,
238.000000000000,652.000000000000,
-1009.00000000000,-404.000000000000,
463.000000000000,-805.000000000000,
-683.000000000000,349.000000000000,
150.000000000000,-336.000000000000,
672.000000000000,-320.000000000000,
-547.000000000000,741.000000000000,
-120.000000000000,-659.000000000000,
137.000000000000,-988.000000000000,
1119.00000000000,83.0000000000000,
714.000000000000,212.000000000000,
391.000000000000,-593.000000000000,
-270.000000000000,-586.000000000000,
-192.000000000000,1078.00000000000,
-898.000000000000,488.000000000000,
-1157.00000000000,445.000000000000,
879.000000000000,-606.000000000000,
7.00000000000000,-533.000000000000,
-411.000000000000,1004.00000000000,
-573.000000000000,176.000000000000,
-802.000000000000,299.000000000000,
303.000000000000,115.000000000000,
-351.000000000000,481.000000000000,
-636.000000000000,658.000000000000,
621.000000000000,171.000000000000,
-142.000000000000,-528.000000000000,
-539.000000000000,-782.000000000000,
-119.000000000000,217.000000000000,
385.000000000000,-255.000000000000,
492.000000000000,55.0000000000000,
-836.000000000000,117.000000000000,
148.000000000000,-119.000000000000,
31.0000000000000,-416.000000000000,
-1038.00000000000,-1139.00000000000,
465.000000000000,-707.000000000000,
976.000000000000,-936.000000000000,
269.000000000000,42.0000000000000,
-373.000000000000,796.000000000000,
-1153.00000000000,-263.000000000000,
-30.0000000000000,-752.000000000000,
596.000000000000,-442.000000000000,
350.000000000000,-332.000000000000,
-229.000000000000,198.000000000000,
-273.000000000000,683.000000000000,
-58.0000000000000,258.000000000000,
-1218.00000000000,-408.000000000000,
-526.000000000000,-341.000000000000,
-241.000000000000,42.0000000000000,
-94.0000000000000,474.000000000000,
-316.000000000000,556.000000000000,
-149.000000000000,-607.000000000000,
1250.00000000000,-274.000000000000,
640.000000000000,1225.00000000000,
349.000000000000,-23.0000000000000,
549.000000000000,-954.000000000000,
1347.00000000000,731.000000000000,
-1.00000000000000,1133.00000000000,
-120.000000000000,-373.000000000000,
928.000000000000,-554.000000000000,
-660.000000000000,885.000000000000,
513.000000000000,747.000000000000,
-221.000000000000,-404.000000000000,
-831.000000000000,539.000000000000,
-538.000000000000,391.000000000000,
47.0000000000000,-798.000000000000,
888.000000000000,286.000000000000,
251.000000000000,-44.0000000000000,
430.000000000000,-89.0000000000000,
-789.000000000000,580.000000000000,
-411.000000000000,-302.000000000000,
44.0000000000000,602.000000000000,
-792.000000000000,-162.000000000000,
-259.000000000000,-1320.00000000000,
722.000000000000,-719.000000000000,
595.000000000000,287.000000000000,
-601.000000000000,899.000000000000,
-16.0000000000000,-338.000000000000,
807.000000000000,4.00000000000000,
-210.000000000000,1359.00000000000,
-160.000000000000,-847.000000000000,
708.000000000000,-327.000000000000,
336.000000000000,173.000000000000,
-96.0000000000000,-400.000000000000,
-314.000000000000,321.000000000000,
522.000000000000,50.0000000000000,
-54.0000000000000,1320.00000000000,
-38.0000000000000,-402.000000000000,
495.000000000000,418.000000000000,
-958.000000000000,953.000000000000,
-2.00000000000000,373.000000000000,
-123.000000000000,199.000000000000,
-517.000000000000,-1262.00000000000,
549.000000000000,726.000000000000,
-585.000000000000,242.000000000000,
-1209.00000000000,284.000000000000,
-679.000000000000,-146.000000000000,
251.000000000000,-1059.00000000000,
576.000000000000,144.000000000000,
-33.0000000000000,-689.000000000000,
-339.000000000000,-356.000000000000,
200.000000000000,481.000000000000,
376.000000000000,-195.000000000000,
846.000000000000,235.000000000000,
750.000000000000,446.000000000000,
-716.000000000000,-91.0000000000000,
-30.0000000000000,559.000000000000,
148.000000000000,59.0000000000000,
-280.000000000000,-314.000000000000,
1003.00000000000,-443.000000000000,
997.000000000000,-377.000000000000,
165.000000000000,845.000000000000,
318.000000000000,1178.00000000000,
472.000000000000,-72.0000000000000,
-351.000000000000,-176.000000000000,
-301.000000000000,464.000000000000,
590.000000000000,-633.000000000000,
-384.000000000000,317.000000000000,
-1064.00000000000,555.000000000000,
758.000000000000,-332.000000000000,
-130.000000000000,674.000000000000,
-1090.00000000000,175.000000000000,
-132.000000000000,-562.000000000000,
878.000000000000,-501.000000000000,
876.000000000000,-471.000000000000,
-282.000000000000,-562.000000000000,
1217.00000000000,-548.000000000000,
-76.0000000000000,170.000000000000,
-584.000000000000,-7.00000000000000,
-735.000000000000,-315.000000000000,
-726.000000000000,977.000000000000,
264.000000000000,-673.000000000000,
-957.000000000000,-1036.00000000000,
1110.00000000000,-109.000000000000,
761.000000000000,-80.0000000000000,
628.000000000000,1402.00000000000,
-58.0000000000000,579.000000000000,
-1159.00000000000,-459.000000000000,
192.000000000000,-905.000000000000,
-691.000000000000,-536.000000000000,
216.000000000000,-1258.00000000000,
929.000000000000,-151.000000000000,
-177.000000000000,831.000000000000,
390.000000000000,-1021.00000000000,
478.000000000000,702.000000000000,
-490.000000000000,-234.000000000000,
384.000000000000,-223.000000000000,
467.000000000000,1049.00000000000,
-121.000000000000,-371.000000000000,
437.000000000000,-105.000000000000,
367.000000000000,288.000000000000,
-339.000000000000,1087.00000000000,
-562.000000000000,108.000000000000,
-421.000000000000,-921.000000000000,
104.000000000000,-215.000000000000,
513.000000000000,775.000000000000,
-470.000000000000,-120.000000000000,
-762.000000000000,-876.000000000000,
958.000000000000,727.000000000000,
17.0000000000000,392.000000000000,
-809.000000000000,157.000000000000,
1081.00000000000,-683.000000000000,
802.000000000000,-598.000000000000,
961.000000000000,750.000000000000,
717.000000000000,135.000000000000,
230.000000000000,-385.000000000000,
24.0000000000000,-786.000000000000,
-751.000000000000,625.000000000000,
-238.000000000000,704.000000000000,
-158.000000000000,-240.000000000000,
1216.00000000000,-231.000000000000,
444.000000000000,-571.000000000000,
29.0000000000000,145.000000000000,
-5.00000000000000,-752.000000000000,
-727.000000000000,-427.000000000000,
903.000000000000,-278.000000000000,
532.000000000000,353.000000000000,
773.000000000000,960.000000000000,
41.0000000000000,489.000000000000,
505.000000000000,885.000000000000,
-28.0000000000000,-194.000000000000,
-978.000000000000,30.0000000000000,
918.000000000000,-145.000000000000,
-172.000000000000,758.000000000000,
236.000000000000,1088.00000000000,
-297.000000000000,399.000000000000,
-1075.00000000000,906.000000000000,
-713.000000000000,-1032.00000000000,
-450.000000000000,-145.000000000000,
848.000000000000,-783.000000000000,
520.000000000000,-772.000000000000,
1272.00000000000,295.000000000000,
691.000000000000,-14.0000000000000,
88.0000000000000,1416.00000000000,
-1102.00000000000,-97.0000000000000,
-270.000000000000,-127.000000000000,
1269.00000000000,-1022.00000000000,
-238.000000000000,439.000000000000,
957.000000000000,556.000000000000,
-200.000000000000,-409.000000000000,
-94.0000000000000,1593.00000000000,
409.000000000000,-426.000000000000,
-499.000000000000,959.000000000000,
840.000000000000,640.000000000000,
-159.000000000000,715.000000000000,
-1121.00000000000,1081.00000000000,
-716.000000000000,-477.000000000000,
-349.000000000000,-308.000000000000,
464.000000000000,-1240.00000000000,
445.000000000000,352.000000000000,
-872.000000000000,367.000000000000,
-198.000000000000,-590.000000000000,
223.000000000000,-143.000000000000,
-848.000000000000,-114.000000000000,
-701.000000000000,3.00000000000000,
-700.000000000000,-612.000000000000,
-705.000000000000,-895.000000000000,
-243.000000000000,132.000000000000,
-117.000000000000,-213.000000000000,
-306.000000000000,-442.000000000000,
8.00000000000000,702.000000000000,
30.0000000000000,-367.000000000000,
-168.000000000000,-21.0000000000000,
532.000000000000,696.000000000000,
-209.000000000000,-505.000000000000,
-525.000000000000,824.000000000000,
830.000000000000,-83.0000000000000,
518.000000000000,-822.000000000000,
1092.00000000000,60.0000000000000,
1157.00000000000,-414.000000000000,
119.000000000000,1432.00000000000,
-990.000000000000,-320.000000000000,
-947.000000000000,-351.000000000000,
785.000000000000,3.00000000000000,
9.00000000000000,-857.000000000000,
627.000000000000,-58.0000000000000,
469.000000000000,-828.000000000000,
-963.000000000000,-89.0000000000000,
510.000000000000,-491.000000000000,
292.000000000000,818.000000000000,
-904.000000000000,846.000000000000,
-299.000000000000,638.000000000000,
451.000000000000,943.000000000000,
187.000000000000,-469.000000000000,
613.000000000000,483.000000000000,
-837.000000000000,-326.000000000000,
-642.000000000000,-772.000000000000,
879.000000000000,660.000000000000,
-548.000000000000,9.00000000000000,
526.000000000000,-384.000000000000,
1246.00000000000,779.000000000000,
-296.000000000000,590.000000000000,
-306.000000000000,346.000000000000,
-249.000000000000,-123.000000000000,
151.000000000000,-675.000000000000,
560.000000000000,782.000000000000,
-444.000000000000,1028.00000000000,
-738.000000000000,-186.000000000000,
-388.000000000000,-787.000000000000,
-48.0000000000000,-273.000000000000,
-438.000000000000,748.000000000000,
-480.000000000000,-752.000000000000,
515.000000000000,-539.000000000000,
-597.000000000000,893.000000000000,
-800.000000000000,140.000000000000,
-390.000000000000,506.000000000000,
-194.000000000000,496.000000000000,
330.000000000000,851.000000000000,
-375.000000000000,478.000000000000,
469.000000000000,-632.000000000000,
631.000000000000,122.000000000000,
-740.000000000000,661.000000000000,
-276.000000000000,-998.000000000000,
-529.000000000000,-1039.00000000000,
-212.000000000000,918.000000000000,
557.000000000000,-173.000000000000,
-1161.00000000000,-185.000000000000,
-55.0000000000000,-502.000000000000,
645.000000000000,-918.000000000000,
-203.000000000000,1128.00000000000,
-708.000000000000,-94.0000000000000,
233.000000000000,-767.000000000000,
881.000000000000,-396.000000000000,
-639.000000000000,-90.0000000000000,
212.000000000000,-507.000000000000,
475.000000000000,-414.000000000000,
565.000000000000,1342.00000000000,
215.000000000000,773.000000000000,
-649.000000000000,1075.00000000000,
-148.000000000000,572.000000000000,
215.000000000000,-256.000000000000,
280.000000000000,-908.000000000000,
-660.000000000000,-911.000000000000,
-204.000000000000,-353.000000000000,
376.000000000000,-430.000000000000,
523.000000000000,362.000000000000,
1068.00000000000,-422.000000000000,
731.000000000000,-54.0000000000000,
-541.000000000000,1026.00000000000,
-1190.00000000000,-868.000000000000,
25.0000000000000,-607.000000000000,
-275.000000000000,602.000000000000,
-133.000000000000,-365.000000000000,
193.000000000000,728.000000000000,
-62.0000000000000,-29.0000000000000,
283.000000000000,-262.000000000000,
-869.000000000000,1005.00000000000,
-40.0000000000000,-702.000000000000,
-297.000000000000,-442.000000000000,
-7.00000000000000,104.000000000000,
950.000000000000,-826.000000000000,
-604.000000000000,-697.000000000000,
159.000000000000,-356.000000000000,
-112.000000000000,491.000000000000,
-534.000000000000,263.000000000000,
-173.000000000000,-482.000000000000,
-376.000000000000,783.000000000000,
-704.000000000000,-501.000000000000,
-784.000000000000,-1004.00000000000,
210.000000000000,-1137.00000000000,
717.000000000000,-976.000000000000,
1013.00000000000,426.000000000000,
394.000000000000,468.000000000000,
-807.000000000000,667.000000000000,
-143.000000000000,-136.000000000000,
551.000000000000,528.000000000000,
-89.0000000000000,-56.0000000000000,
-101.000000000000,517.000000000000,
140.000000000000,377.000000000000,
-260.000000000000,-1227.00000000000,
537.000000000000,562.000000000000,
504.000000000000,-619.000000000000,
791.000000000000,-318.000000000000,
1024.00000000000,-164.000000000000,
-7.00000000000000,-232.000000000000,
1074.00000000000,546.000000000000,
-730.000000000000,27.0000000000000,
-286.000000000000,479.000000000000,
124.000000000000,-915.000000000000,
-1091.00000000000,374.000000000000,
563.000000000000,930.000000000000,
-342.000000000000,436.000000000000,
278.000000000000,519.000000000000,
-750.000000000000,117.000000000000,
-596.000000000000,608.000000000000,
-271.000000000000,-154.000000000000,
-428.000000000000,-437.000000000000,
984.000000000000,-687.000000000000,
-441.000000000000,556.000000000000,
260.000000000000,749.000000000000,
574.000000000000,-645.000000000000,
-191.000000000000,-451.000000000000,
-567.000000000000,-800.000000000000,
-823.000000000000,-302.000000000000,
-423.000000000000,117.000000000000,
309.000000000000,-280.000000000000,
916.000000000000,-3.00000000000000,
639.000000000000,146.000000000000,
1135.00000000000,-99.0000000000000,
-265.000000000000,893.000000000000,
-832.000000000000,640.000000000000,
-171.000000000000,-851.000000000000,
-683.000000000000,343.000000000000,
74.0000000000000,966.000000000000,
-1184.00000000000,43.0000000000000,
-726.000000000000,-743.000000000000,
606.000000000000,-1222.00000000000,
-483.000000000000,591.000000000000,
-79.0000000000000,-159.000000000000,
918.000000000000,-843.000000000000,
856.000000000000,267.000000000000,
-286.000000000000,1388.00000000000,
40.0000000000000,273.000000000000,
1065.00000000000,-840.000000000000,
161.000000000000,1080.00000000000,
-420.000000000000,-749.000000000000,
177.000000000000,-948.000000000000,
455.000000000000,-287.000000000000,
754.000000000000,-181.000000000000,
75.0000000000000,1375.00000000000,
-777.000000000000,-437.000000000000,
172.000000000000,-13.0000000000000,
-128.000000000000,710.000000000000,
-12.0000000000000,-158.000000000000,
807.000000000000,219.000000000000,
-535.000000000000,497.000000000000,
283.000000000000,-434.000000000000,
927.000000000000,-301.000000000000,
-560.000000000000,594.000000000000,
403.000000000000,-502.000000000000,
576.000000000000,312.000000000000,
-376.000000000000,620.000000000000,
-304.000000000000,921.000000000000,
-467.000000000000,585.000000000000,
151.000000000000,-375.000000000000,
227.000000000000,278.000000000000,
-145.000000000000,-1119.00000000000,
453.000000000000,-541.000000000000,
-86.0000000000000,-135.000000000000,
242.000000000000,-589.000000000000,
1009.00000000000,-11.0000000000000,
407.000000000000,-793.000000000000,
1039.00000000000,-263.000000000000,
140.000000000000,38.0000000000000,
-324.000000000000,552.000000000000,
787.000000000000,778.000000000000,
-1542.00000000000,778.000000000000,
-1036.00000000000,-279.000000000000,
-186.000000000000,-845.000000000000,
263.000000000000,163.000000000000,
435.000000000000,-504.000000000000,
-516.000000000000,612.000000000000,
736.000000000000,-23.0000000000000,
286.000000000000,-275.000000000000,
-63.0000000000000,248.000000000000,
-546.000000000000,-327.000000000000,
543.000000000000,617.000000000000,
673.000000000000,-172.000000000000,
-124.000000000000,588.000000000000,
1149.00000000000,-379.000000000000,
448.000000000000,-290.000000000000,
174.000000000000,230.000000000000,
319.000000000000,-102.000000000000,
-451.000000000000,663.000000000000,
-205.000000000000,-1094.00000000000,
643.000000000000,-578.000000000000,
394.000000000000,-192.000000000000,
-159.000000000000,465.000000000000,
-543.000000000000,722.000000000000,
-992.000000000000,187.000000000000,
236.000000000000,1116.00000000000,
690.000000000000,520.000000000000,
-67.0000000000000,1080.00000000000,
-84.0000000000000,-66.0000000000000,
306.000000000000,-89.0000000000000,
999.000000000000,121.000000000000,
645.000000000000,177.000000000000,
656.000000000000,380.000000000000,
743.000000000000,-794.000000000000,
-339.000000000000,725.000000000000,
-449.000000000000,-20.0000000000000,
613.000000000000,-178.000000000000,
271.000000000000,263.000000000000,
-605.000000000000,-578.000000000000,
-236.000000000000,805.000000000000,
-1168.00000000000,250.000000000000,
-571.000000000000,-969.000000000000,
855.000000000000,539.000000000000,
193.000000000000,1338.00000000000,
-144.000000000000,446.000000000000,
-585.000000000000,135.000000000000,
194.000000000000,93.0000000000000,
-925.000000000000,-823.000000000000,
-31.0000000000000,-876.000000000000,
549.000000000000,414.000000000000,
-858.000000000000,-111.000000000000,
1443.00000000000,-760.000000000000,
-28.0000000000000,747.000000000000,
226.000000000000,486.000000000000,
-198.000000000000,-308.000000000000,
-642.000000000000,694.000000000000,
510.000000000000,191.000000000000,
-646.000000000000,61.0000000000000,
-427.000000000000,-854.000000000000,
-961.000000000000,-904.000000000000,
1189.00000000000,-481.000000000000,
732.000000000000,-661.000000000000,
756.000000000000,1402.00000000000,
367.000000000000,-190.000000000000,
-1108.00000000000,-115.000000000000,
1261.00000000000,-28.0000000000000,
-432.000000000000,-448.000000000000,
578.000000000000,734.000000000000,
269.000000000000,-128.000000000000,
-1198.00000000000,-91.0000000000000,
164.000000000000,-990.000000000000,
423.000000000000,-515.000000000000,
909.000000000000,-154.000000000000,
-492.000000000000,353.000000000000,
-879.000000000000,633.000000000000,
-214.000000000000,-397.000000000000,
142.000000000000,-314.000000000000,
203.000000000000,61.0000000000000,
567.000000000000,1391.00000000000,
-357.000000000000,222.000000000000,
-907.000000000000,118.000000000000,
478.000000000000,1059.00000000000,
-605.000000000000,-289.000000000000,
-926.000000000000,-691.000000000000,
473.000000000000,77.0000000000000,
308.000000000000,819.000000000000,
-655.000000000000,650.000000000000,
29.0000000000000,193.000000000000,
1052.00000000000,-187.000000000000,
-3.00000000000000,-310.000000000000,
865.000000000000,242.000000000000,
152.000000000000,310.000000000000,
-950.000000000000,-411.000000000000,
392.000000000000,-1314.00000000000,
-6.00000000000000,-169.000000000000,
665.000000000000,182.000000000000,
-162.000000000000,-921.000000000000,
664.000000000000,-234.000000000000,
849.000000000000,106.000000000000,
-384.000000000000,629.000000000000,
143.000000000000,-276.000000000000,
-128.000000000000,15.0000000000000,
724.000000000000,-113.000000000000,
-261.000000000000,-417.000000000000,
-438.000000000000,1229.00000000000,
-907.000000000000,261.000000000000,
-1191.00000000000,-506.000000000000,
-107.000000000000,-422.000000000000,
-698.000000000000,-763.000000000000,
-40.0000000000000,-752.000000000000,
671.000000000000,320.000000000000,
-621.000000000000,1144.00000000000,
-376.000000000000,489.000000000000,
720.000000000000,98.0000000000000,
293.000000000000,629.000000000000,
212.000000000000,-92.0000000000000,
182.000000000000,-453.000000000000,
134.000000000000,-41.0000000000000,
-165.000000000000,-1012.00000000000,
-774.000000000000,-974.000000000000,
-508.000000000000,-415.000000000000,
-445.000000000000,-462.000000000000,
-1046.00000000000,466.000000000000,
-798.000000000000,683.000000000000,
141.000000000000,-445.000000000000,
80.0000000000000,-408.000000000000,
-775.000000000000,-357.000000000000,
134.000000000000,-1128.00000000000,
1183.00000000000,-923.000000000000,
354.000000000000,-44.0000000000000,
787.000000000000,10.0000000000000,
906.000000000000,202.000000000000,
-404.000000000000,-237.000000000000,
-191.000000000000,-1228.00000000000,
174.000000000000,-38.0000000000000,
-70.0000000000000,786.000000000000,
-41.0000000000000,-247.000000000000,
-517.000000000000,-1121.00000000000,
-506.000000000000,-560.000000000000,
-94.0000000000000,-589.000000000000,
-112.000000000000,-872.000000000000,
1210.00000000000,398.000000000000,
147.000000000000,83.0000000000000,
-546.000000000000,-15.0000000000000,
1121.00000000000,566.000000000000,
-90.0000000000000,-386.000000000000,
714.000000000000,63.0000000000000,
536.000000000000,1037.00000000000,
77.0000000000000,415.000000000000,
-36.0000000000000,-733.000000000000,
-938.000000000000,-156.000000000000,
219.000000000000,72.0000000000000,
-184.000000000000,-520.000000000000,
1016.00000000000,-318.000000000000,
1034.00000000000,200.000000000000,
-227.000000000000,938.000000000000,
198.000000000000,671.000000000000,
-68.0000000000000,-497.000000000000,
-595.000000000000,-253.000000000000,
471.000000000000,1365.00000000000,
927.000000000000,433.000000000000,
-921.000000000000,-654.000000000000,
67.0000000000000,-174.000000000000,
432.000000000000,-411.000000000000,
-209.000000000000,352.000000000000,
82.0000000000000,-222.000000000000,
-830.000000000000,-705.000000000000,
413.000000000000,348.000000000000,
61.0000000000000,-127.000000000000,
-672.000000000000,-834.000000000000,
342.000000000000,-1225.00000000000,
938.000000000000,-173.000000000000,
644.000000000000,135.000000000000,
58.0000000000000,-10.0000000000000,
808.000000000000,33.0000000000000,
-880.000000000000,242.000000000000,
-845.000000000000,783.000000000000,
739.000000000000,342.000000000000,
-128.000000000000,1168.00000000000,
-882.000000000000,581.000000000000,
-918.000000000000,-695.000000000000,
-119.000000000000,-1331.00000000000,
324.000000000000,-498.000000000000,
-232.000000000000,990.000000000000,
-149.000000000000,-199.000000000000,
1246.00000000000,-164.000000000000,
461.000000000000,1042.00000000000,
-1137.00000000000,-244.000000000000,
-221.000000000000,-1339.00000000000,
427.000000000000,33.0000000000000,
397.000000000000,-208.000000000000,
-123.000000000000,-674.000000000000,
-252.000000000000,985.000000000000,
-390.000000000000,-514.000000000000,
-137.000000000000,-1053.00000000000,
1235.00000000000,1239.00000000000,
257.000000000000,233.000000000000,
-305.000000000000,-439.000000000000,
-484.000000000000,130.000000000000,
-743.000000000000,-1019.00000000000,
-673.000000000000,-459.000000000000,
-612.000000000000,708.000000000000,
43.0000000000000,-918.000000000000,
-839.000000000000,-344.000000000000,
479.000000000000,220.000000000000,
752.000000000000,-1040.00000000000,
961.000000000000,105.000000000000,
910.000000000000,-747.000000000000,
-559.000000000000,-524.000000000000,
594.000000000000,-76.0000000000000,
-60.0000000000000,445.000000000000,
-37.0000000000000,853.000000000000,
391.000000000000,-470.000000000000,
95.0000000000000,134.000000000000,
503.000000000000,-717.000000000000,
117.000000000000,-12.0000000000000,
305.000000000000,564.000000000000,
48.0000000000000,-453.000000000000,
-189.000000000000,-675.000000000000,
651.000000000000,-927.000000000000,
1177.00000000000,-226.000000000000,
-341.000000000000,-651.000000000000,
435.000000000000,-436.000000000000,
1245.00000000000,-718.000000000000,
-762.000000000000,-90.0000000000000,
1055.00000000000,268.000000000000,
-106.000000000000,-695.000000000000,
-124.000000000000,134.000000000000,
1462.00000000000,-198.000000000000,
81.0000000000000,1107.00000000000,
990.000000000000,576.000000000000,
128.000000000000,409.000000000000,
-497.000000000000,934.000000000000,
-658.000000000000,-3.00000000000000,
489.000000000000,654.000000000000,
179.000000000000,-762.000000000000,
-236.000000000000,-187.000000000000,
1123.00000000000,1023.00000000000,
171.000000000000,312.000000000000,
110.000000000000,-353.000000000000,
-1131.00000000000,-657.000000000000,
598.000000000000,317.000000000000,
280.000000000000,289.000000000000,
-535.000000000000,561.000000000000,
615.000000000000,750.000000000000,
-1602.00000000000,243.000000000000,
525.000000000000,-702.000000000000,
681.000000000000,333.000000000000,
-504.000000000000,1017.00000000000,
331.000000000000,-157.000000000000,
66.0000000000000,956.000000000000,
644.000000000000,-13.0000000000000,
-107.000000000000,686.000000000000,
-848.000000000000,-52.0000000000000,
-256.000000000000,-594.000000000000,
939.000000000000,1315.00000000000,
-340.000000000000,-1211.00000000000,
-794.000000000000,-227.000000000000,
438.000000000000,-258.000000000000,
336.000000000000,198.000000000000,
465.000000000000,816.000000000000,
122.000000000000,-1199.00000000000,
337.000000000000,-105.000000000000,
-869.000000000000,615.000000000000,
-494.000000000000,270.000000000000,
1091.00000000000,-299.000000000000,
144.000000000000,825.000000000000,
894.000000000000,-33.0000000000000,
444.000000000000,204.000000000000,
-331.000000000000,1217.00000000000,
473.000000000000,-777.000000000000,
686.000000000000,-79.0000000000000,
611.000000000000,572.000000000000,
49.0000000000000,702.000000000000,
-99.0000000000000,577.000000000000,
10.0000000000000,704.000000000000,
-705.000000000000,508.000000000000,
-521.000000000000,-162.000000000000,
374.000000000000,774.000000000000,
-304.000000000000,-594.000000000000,
-1023.00000000000,-730.000000000000,
-490.000000000000,-199.000000000000,
378.000000000000,123.000000000000,
169.000000000000,-35.0000000000000,
312.000000000000,-89.0000000000000,
351.000000000000,1029.00000000000,
91.0000000000000,47.0000000000000,
815.000000000000,496.000000000000,
427.000000000000,594.000000000000,
-877.000000000000,220.000000000000,
-345.000000000000,-181.000000000000,
-532.000000000000,-414.000000000000,
-1053.00000000000,746.000000000000,
-533.000000000000,-1362.00000000000,
-270.000000000000,-366.000000000000,
-354.000000000000,-109.000000000000,
-731.000000000000,-1256.00000000000,
1124.00000000000,-239.000000000000,
5.00000000000000,-328.000000000000,
-612.000000000000,97.0000000000000,
1001.00000000000,-77.0000000000000,
277.000000000000,1133.00000000000,
772.000000000000,141.000000000000,
340.000000000000,-424.000000000000,
-189.000000000000,78.0000000000000,
280.000000000000,-420.000000000000,
580.000000000000,531.000000000000,
-309.000000000000,158.000000000000,
-289.000000000000,1061.00000000000,
445.000000000000,224.000000000000,
210.000000000000,-971.000000000000,
910.000000000000,306.000000000000,
388.000000000000,889.000000000000,
372.000000000000,796.000000000000,
162.000000000000,-53.0000000000000,
-126.000000000000,-611.000000000000,
-647.000000000000,-171.000000000000,
-1354.00000000000,427.000000000000,
408.000000000000,21.0000000000000,
-709.000000000000,-1165.00000000000,
841.000000000000,-452.000000000000,
584.000000000000,822.000000000000,
-389.000000000000,67.0000000000000,
1068.00000000000,-564.000000000000,
-1228.00000000000,601.000000000000,
-176.000000000000,-555.000000000000,
-201.000000000000,-1006.00000000000,
288.000000000000,701.000000000000,
123.000000000000,113.000000000000,
-908.000000000000,546.000000000000,
664.000000000000,-273.000000000000,
-259.000000000000,-644.000000000000,
-267.000000000000,60.0000000000000,
-278.000000000000,243.000000000000,
205.000000000000,236.000000000000,
662.000000000000,-331.000000000000,
529.000000000000,1550.00000000000,
55.0000000000000,700.000000000000,
-885.000000000000,-542.000000000000,
-31.0000000000000,-1364.00000000000,
1057.00000000000,-502.000000000000,
5.00000000000000,803.000000000000,
-1141.00000000000,-658.000000000000,
-535.000000000000,-579.000000000000,
-47.0000000000000,-906.000000000000,
569.000000000000,-173.000000000000,
894.000000000000,-168.000000000000,
772.000000000000,-382.000000000000,
1043.00000000000,430.000000000000,
-588.000000000000,-498.000000000000,
-619.000000000000,-334.000000000000,
979.000000000000,-978.000000000000,
-359.000000000000,-464.000000000000,
-548.000000000000,617.000000000000,
468.000000000000,650.000000000000,
-210.000000000000,1089.00000000000,
-501.000000000000,599.000000000000,
-669.000000000000,-683.000000000000,
310.000000000000,-942.000000000000,
1133.00000000000,-287.000000000000,
258.000000000000,-267.000000000000,
535.000000000000,408.000000000000,
-790.000000000000,651.000000000000,
-498.000000000000,152.000000000000,
796.000000000000,349.000000000000,
332.000000000000,813.000000000000,
687.000000000000,378.000000000000,
214.000000000000,750.000000000000,
-220.000000000000,1073.00000000000,
-920.000000000000,197.000000000000,
-846.000000000000,-962.000000000000,
-499.000000000000,-884.000000000000,
-401.000000000000,179.000000000000,
36.0000000000000,-487.000000000000,
464.000000000000,-950.000000000000,
571.000000000000,-170.000000000000,
45.0000000000000,-1115.00000000000,
-302.000000000000,-943.000000000000,
1136.00000000000,280.000000000000,
165.000000000000,-845.000000000000,
-336.000000000000,49.0000000000000,
987.000000000000,471.000000000000,
-207.000000000000,195.000000000000,
795.000000000000,-207.000000000000,
-193.000000000000,-754.000000000000,
26.0000000000000,1313.00000000000,
523.000000000000,445.000000000000,
-982.000000000000,-322.000000000000,
922.000000000000,-865.000000000000,
429.000000000000,-124.000000000000,
-51.0000000000000,71.0000000000000,
85.0000000000000,-764.000000000000,
479.000000000000,1432.00000000000,
553.000000000000,1000.00000000000,
-6.00000000000000,-37.0000000000000,
-269.000000000000,-110.000000000000,
-504.000000000000,109.000000000000,
556.000000000000,-595.000000000000,
-580.000000000000,-778.000000000000,
-773.000000000000,81.0000000000000,
-439.000000000000,-368.000000000000,
-789.000000000000,878.000000000000,
-603.000000000000,-687.000000000000,
-705.000000000000,-919.000000000000,
918.000000000000,-408.000000000000,
73.0000000000000,-1171.00000000000,
-55.0000000000000,-446.000000000000,
963.000000000000,-175.000000000000,
17.0000000000000,1151.00000000000,
-285.000000000000,-326.000000000000,
892.000000000000,-382.000000000000,
1281.00000000000,-126.000000000000,
-282.000000000000,-921.000000000000,
-206.000000000000,-106.000000000000,
-89.0000000000000,-796.000000000000,
707.000000000000,-422.000000000000,
748.000000000000,-623.000000000000,
-766.000000000000,-74.0000000000000,
405.000000000000,624.000000000000,
390.000000000000,534.000000000000,
-20.0000000000000,1253.00000000000,
155.000000000000,-51.0000000000000,
-353.000000000000,-920.000000000000,
124.000000000000,271.000000000000,
699.000000000000,101.000000000000,
236.000000000000,170.000000000000,
-225.000000000000,184.000000000000,
40.0000000000000,-576.000000000000,
58.0000000000000,937.000000000000,
-571.000000000000,784.000000000000,
-25.0000000000000,-950.000000000000,
651.000000000000,1067.00000000000,
-47.0000000000000,587.000000000000,
35.0000000000000,-900.000000000000,
582.000000000000,-816.000000000000,
833.000000000000,-797.000000000000,
-157.000000000000,856.000000000000,
-214.000000000000,133.000000000000,
220.000000000000,-301.000000000000,
-437.000000000000,-819.000000000000,
425.000000000000,115.000000000000,
557.000000000000,1443.00000000000,
-1292.00000000000,207.000000000000,
-317.000000000000,611.000000000000,
191.000000000000,-369.000000000000,
-1057.00000000000,672.000000000000,
-154.000000000000,188.000000000000,
-5.00000000000000,-735.000000000000,
908.000000000000,536.000000000000,
-220.000000000000,-168.000000000000,
-269.000000000000,-787.000000000000,
184.000000000000,-1519.00000000000,
-291.000000000000,135.000000000000,
1228.00000000000,-387.000000000000,
-459.000000000000,196.000000000000,
190.000000000000,798.000000000000,
83.0000000000000,-967.000000000000,
-1081.00000000000,424.000000000000,
79.0000000000000,-398.000000000000,
820.000000000000,161.000000000000,
-171.000000000000,469.000000000000,
-1311.00000000000,679.000000000000,
583.000000000000,101.000000000000,
19.0000000000000,-671.000000000000,
84.0000000000000,1205.00000000000,
-445.000000000000,314.000000000000,
-1285.00000000000,231.000000000000,
-491.000000000000,-1045.00000000000,
-868.000000000000,-868.000000000000,
906.000000000000,676.000000000000,
411.000000000000,-251.000000000000,
530.000000000000,-357.000000000000,
392.000000000000,-901.000000000000,
-850.000000000000,-747.000000000000,
238.000000000000,-502.000000000000,
365.000000000000,-624.000000000000,
483.000000000000,-287.000000000000,
-231.000000000000,249.000000000000,
67.0000000000000,-257.000000000000,
-502.000000000000,-624.000000000000,
-855.000000000000,688.000000000000,
-400.000000000000,212.000000000000,
-1208.00000000000,667.000000000000,
169.000000000000,220.000000000000,
279.000000000000,-104.000000000000,
272.000000000000,1128.00000000000,
1224.00000000000,-387.000000000000,
134.000000000000,-157.000000000000,
-477.000000000000,370.000000000000,
230.000000000000,511.000000000000,
5.00000000000000,502.000000000000,
-246.000000000000,698.000000000000,
580.000000000000,529.000000000000,
-538.000000000000,-1185.00000000000,
-325.000000000000,-974.000000000000,
348.000000000000,-456.000000000000,
-110.000000000000,-770.000000000000,
349.000000000000,473.000000000000,
-69.0000000000000,726.000000000000,
649.000000000000,120.000000000000,
435.000000000000,1438.00000000000,
-195.000000000000,629.000000000000,
19.0000000000000,-649.000000000000,
-584.000000000000,469.000000000000,
-229.000000000000,-1099.00000000000,
-179.000000000000,-727.000000000000,
360.000000000000,1051.00000000000,
656.000000000000,-534.000000000000,
-583.000000000000,-84.0000000000000,
85.0000000000000,484.000000000000,
143.000000000000,1270.00000000000,
-733.000000000000,-130.000000000000,
115.000000000000,-454.000000000000,
182.000000000000,-155.000000000000,
-325.000000000000,-975.000000000000,
23.0000000000000,1108.00000000000,
-47.0000000000000,-722.000000000000,
786.000000000000,-128.000000000000,
958.000000000000,173.000000000000,
-672.000000000000,-83.0000000000000,
435.000000000000,481.000000000000,
104.000000000000,-671.000000000000,
102.000000000000,1417.00000000000,
-50.0000000000000,128.000000000000,
-755.000000000000,-947.000000000000,
651.000000000000,-467.000000000000,
-922.000000000000,310.000000000000,
-39.0000000000000,202.000000000000,
278.000000000000,148.000000000000,
-457.000000000000,822.000000000000,
927.000000000000,-909.000000000000,
271.000000000000,366.000000000000,
-590.000000000000,171.000000000000,
-470.000000000000,221.000000000000,
169.000000000000,920.000000000000,
428.000000000000,-929.000000000000,
43.0000000000000,185.000000000000,
478.000000000000,887.000000000000,
197.000000000000,31.0000000000000,
-667.000000000000,447.000000000000,
46.0000000000000,190.000000000000,
-589.000000000000,-511.000000000000,
-1024.00000000000,378.000000000000,
453.000000000000,181.000000000000,
-670.000000000000,-737.000000000000,
65.0000000000000,-112.000000000000,
929.000000000000,751.000000000000,
-873.000000000000,208.000000000000,
954.000000000000,-1382.00000000000,
41.0000000000000,-355.000000000000,
-1122.00000000000,348.000000000000,
-229.000000000000,-1083.00000000000,
-530.000000000000,463.000000000000,
-1099.00000000000,427.000000000000,
-579.000000000000,-1281.00000000000,
1269.00000000000,154.000000000000,
-255.000000000000,-12.0000000000000,
476.000000000000,-652.000000000000,
-193.000000000000,223.000000000000,
-696.000000000000,631.000000000000,
125.000000000000,406.000000000000,
-952.000000000000,-494.000000000000,
1261.00000000000,-712.000000000000,
2.00000000000000,358.000000000000,
-15.0000000000000,90.0000000000000,
1020.00000000000,-861.000000000000,
-270.000000000000,280.000000000000,
-844.000000000000,-59.0000000000000,
-1119.00000000000,-621.000000000000,
288.000000000000,-527.000000000000,
580.000000000000,95.0000000000000,
1032.00000000000,162.000000000000,
378.000000000000,-876.000000000000,
-288.000000000000,-206.000000000000,
202.000000000000,-997.000000000000,
205.000000000000,-359.000000000000,
274.000000000000,-2.00000000000000,
-457.000000000000,-1174.00000000000,
625.000000000000,277.000000000000,
148.000000000000,997.000000000000,
-1438.00000000000,751.000000000000,
-539.000000000000,225.000000000000,
885.000000000000,-155.000000000000,
493.000000000000,-364.000000000000,
-495.000000000000,-614.000000000000,
712.000000000000,-962.000000000000,
42.0000000000000,-905.000000000000,
-811.000000000000,-137.000000000000,
149.000000000000,-500.000000000000,
17.0000000000000,-392.000000000000,
199.000000000000,778.000000000000,
213.000000000000,578.000000000000,
159.000000000000,-439.000000000000,
271.000000000000,315.000000000000,
638.000000000000,1000.00000000000,
280.000000000000,-233.000000000000,
780.000000000000,-170.000000000000,
1283.00000000000,-241.000000000000,
-365.000000000000,521.000000000000,
-708.000000000000,536.000000000000,
-423.000000000000,-1451.00000000000,
607.000000000000,-655.000000000000,
1271.00000000000,-271.000000000000,
446.000000000000,-394.000000000000,
-293.000000000000,620.000000000000,
-735.000000000000,102.000000000000,
869.000000000000,-913.000000000000,
-488.000000000000,-323.000000000000,
-316.000000000000,740.000000000000,
983.000000000000,-116.000000000000,
423.000000000000,-91.0000000000000,
1159.00000000000,48.0000000000000,
356.000000000000,-102.000000000000,
512.000000000000,-843.000000000000,
614.000000000000,-463.000000000000,
228.000000000000,760.000000000000,
123.000000000000,-551.000000000000,
750.000000000000,909.000000000000,
362.000000000000,1168.00000000000,
-1060.00000000000,-456.000000000000,
726.000000000000,300.000000000000,
687.000000000000,562.000000000000,
-39.0000000000000,703.000000000000,
-473.000000000000,460.000000000000,
386.000000000000,-519.000000000000,
902.000000000000,-413.000000000000,
-1404.00000000000,792.000000000000,
-312.000000000000,-35.0000000000000,
347.000000000000,-841.000000000000,
123.000000000000,-139.000000000000,
-773.000000000000,-66.0000000000000,
-522.000000000000,872.000000000000,
579.000000000000,-101.000000000000,
-802.000000000000,565.000000000000,
-70.0000000000000,424.000000000000,
-493.000000000000,-1975.00000000000,
-23.0000000000000,-274.000000000000,
596.000000000000,644.000000000000,
-234.000000000000,-309.000000000000,
300.000000000000,-793.000000000000,
762.000000000000,158.000000000000,
-50.0000000000000,845.000000000000,
-1624.00000000000,125.000000000000,
222.000000000000,-467.000000000000,
-412.000000000000,-517.000000000000,
-349.000000000000,-319.000000000000,
1221.00000000000,-676.000000000000,
133.000000000000,774.000000000000,
394.000000000000,215.000000000000,
-770.000000000000,-181.000000000000,
235.000000000000,1253.00000000000,
551.000000000000,240.000000000000,
-77.0000000000000,750.000000000000,
391.000000000000,1137.00000000000,
-44.0000000000000,113.000000000000,
476.000000000000,222.000000000000,
503.000000000000,149.000000000000,
1176.00000000000,-588.000000000000,
325.000000000000,-606.000000000000,
-651.000000000000,72.0000000000000,
-671.000000000000,-439.000000000000,
-1372.00000000000,-27.0000000000000,
-918.000000000000,458.000000000000,
-157.000000000000,-137.000000000000,
550.000000000000,-685.000000000000,
-451.000000000000,-1122.00000000000,
738.000000000000,-266.000000000000,
493.000000000000,105.000000000000,
-765.000000000000,-29.0000000000000,
747.000000000000,238.000000000000,
-183.000000000000,210.000000000000,
740.000000000000,-120.000000000000,
729.000000000000,-253.000000000000,
-107.000000000000,580.000000000000,
-69.0000000000000,203.000000000000,
-404.000000000000,-621.000000000000,
102.000000000000,-761.000000000000,
69.0000000000000,-405.000000000000,
486.000000000000,285.000000000000,
185.000000000000,662.000000000000,
-50.0000000000000,704.000000000000,
401.000000000000,894.000000000000,
-690.000000000000,321.000000000000,
-457.000000000000,-976.000000000000,
165.000000000000,482.000000000000,
-792.000000000000,1.00000000000000,
397.000000000000,-1190.00000000000,
839.000000000000,241.000000000000,
-4.00000000000000,-684.000000000000,
429.000000000000,-102.000000000000,
-16.0000000000000,-847.000000000000,
-232.000000000000,-911.000000000000,
99.0000000000000,600.000000000000,
-805.000000000000,52.0000000000000,
-329.000000000000,-166.000000000000,
864.000000000000,-379.000000000000,
353.000000000000,433.000000000000,
78.0000000000000,407.000000000000,
71.0000000000000,-538.000000000000,
165.000000000000,-847.000000000000,
346.000000000000,-874.000000000000,
1318.00000000000,205.000000000000,
-140.000000000000,450.000000000000,
-1306.00000000000,41.0000000000000,
-297.000000000000,-44.0000000000000,
-561.000000000000,-482.000000000000,
269.000000000000,-443.000000000000,
659.000000000000,525.000000000000,
113.000000000000,3.00000000000000,
730.000000000000,-386.000000000000,
472.000000000000,732.000000000000,
-205.000000000000,-158.000000000000,
38.0000000000000,112.000000000000,
742.000000000000,266.000000000000,
260.000000000000,102.000000000000,
-360.000000000000,353.000000000000,
511.000000000000,-1136.00000000000,
901.000000000000,-383.000000000000,
-36.0000000000000,156.000000000000,
-939.000000000000,204.000000000000,
-763.000000000000,-214.000000000000,
-137.000000000000,533.000000000000,
-503.000000000000,1018.00000000000,
-437.000000000000,343.000000000000,
943.000000000000,1108.00000000000,
688.000000000000,-594.000000000000,
3.00000000000000,4.00000000000000,
252.000000000000,186.000000000000,
-1232.00000000000,-420.000000000000,
-138.000000000000,151.000000000000,
-371.000000000000,-1492.00000000000,
77.0000000000000,-441.000000000000,
1711.00000000000,-429.000000000000,
405.000000000000,-331.000000000000,
1106.00000000000,688.000000000000,
311.000000000000,176.000000000000,
-33.0000000000000,612.000000000000,
-782.000000000000,595.000000000000,
-857.000000000000,564.000000000000,
-713.000000000000,-145.000000000000,
-1120.00000000000,-169.000000000000,
-244.000000000000,-109.000000000000,
-903.000000000000,-786.000000000000,
1111.00000000000,-927.000000000000,
977.000000000000,-703.000000000000,
-375.000000000000,321.000000000000,
-1023.00000000000,379.000000000000,
-808.000000000000,-955.000000000000,
573.000000000000,23.0000000000000,
164.000000000000,57.0000000000000,
968.000000000000,-213.000000000000,
417.000000000000,381.000000000000,
-812.000000000000,132.000000000000,
-428.000000000000,568.000000000000,
35.0000000000000,-841.000000000000,
-498.000000000000,-184.000000000000,
-133.000000000000,-83.0000000000000,
1062.00000000000,-512.000000000000,
707.000000000000,486.000000000000,
284.000000000000,-400.000000000000,
463.000000000000,937.000000000000,
-195.000000000000,1199.00000000000,
-944.000000000000,433.000000000000,
-533.000000000000,-34.0000000000000,
108.000000000000,-791.000000000000,
484.000000000000,56.0000000000000,
-118.000000000000,209.000000000000,
203.000000000000,-325.000000000000,
783.000000000000,697.000000000000,
-225.000000000000,405.000000000000,
188.000000000000,-65.0000000000000,
412.000000000000,-5.00000000000000,
-694.000000000000,-491.000000000000,
482.000000000000,-263.000000000000,
64.0000000000000,-278.000000000000,
-1062.00000000000,556.000000000000,
-401.000000000000,383.000000000000,
-657.000000000000,-670.000000000000,
960.000000000000,-781.000000000000,
1200.00000000000,-100.000000000000,
-310.000000000000,978.000000000000,
-231.000000000000,610.000000000000,
367.000000000000,77.0000000000000,
1239.00000000000,-510.000000000000,
527.000000000000,500.000000000000,
-564.000000000000,1032.00000000000,
-50.0000000000000,54.0000000000000,
-395.000000000000,576.000000000000,
-402.000000000000,569.000000000000,
673.000000000000,602.000000000000,
75.0000000000000,734.000000000000,
-1254.00000000000,696.000000000000,
-746.000000000000,-881.000000000000,
371.000000000000,-1035.00000000000,
795.000000000000,-195.000000000000,
-762.000000000000,-517.000000000000,
-362.000000000000,505.000000000000,
758.000000000000,-700.000000000000,
-782.000000000000,-449.000000000000,
-482.000000000000,409.000000000000,
20.0000000000000,-417.000000000000,
743.000000000000,692.000000000000,
-66.0000000000000,875.000000000000,
-1350.00000000000,261.000000000000,
-375.000000000000,-493.000000000000,
153.000000000000,504.000000000000,
294.000000000000,-101.000000000000,
-333.000000000000,-1024.00000000000,
522.000000000000,401.000000000000,
-443.000000000000,-92.0000000000000,
-76.0000000000000,-121.000000000000,
393.000000000000,37.0000000000000,
-1454.00000000000,-302.000000000000,
184.000000000000,-1598.00000000000,
307.000000000000,59.0000000000000,
229.000000000000,948.000000000000,
434.000000000000,-432.000000000000,
-15.0000000000000,1238.00000000000,
-133.000000000000,-559.000000000000,
-295.000000000000,-854.000000000000,
-478.000000000000,51.0000000000000,
-438.000000000000,-198.000000000000,
1048.00000000000,-46.0000000000000,
-801.000000000000,-180.000000000000,
54.0000000000000,463.000000000000,
742.000000000000,-565.000000000000,
-870.000000000000,366.000000000000,
76.0000000000000,9.00000000000000,
-1203.00000000000,-250.000000000000,
654.000000000000,285.000000000000,
598.000000000000,-927.000000000000,
109.000000000000,1366.00000000000,
82.0000000000000,918.000000000000,
65.0000000000000,-538.000000000000,
1240.00000000000,451.000000000000,
-741.000000000000,1315.00000000000,
-32.0000000000000,541.000000000000,
-1214.00000000000,28.0000000000000,
-59.0000000000000,100.000000000000,
647.000000000000,-1167.00000000000,
-1190.00000000000,756.000000000000,
1045.00000000000,33.0000000000000,
582.000000000000,-309.000000000000,
-188.000000000000,-469.000000000000,
-624.000000000000,-1298.00000000000,
-359.000000000000,100.000000000000,
726.000000000000,-476.000000000000,
336.000000000000,899.000000000000,
-622.000000000000,-510.000000000000,
-96.0000000000000,-877.000000000000,
420.000000000000,544.000000000000,
-508.000000000000,-905.000000000000,
962.000000000000,351.000000000000,
-31.0000000000000,584.000000000000,
-608.000000000000,-503.000000000000,
959.000000000000,401.000000000000,
49.0000000000000,726.000000000000,
-135.000000000000,261.000000000000,
-902.000000000000,253.000000000000,
360.000000000000,-193.000000000000,
-534.000000000000,-329.000000000000,
-694.000000000000,261.000000000000,
1039.00000000000,46.0000000000000,
-648.000000000000,671.000000000000,
48.0000000000000,-70.0000000000000,
-71.0000000000000,-1217.00000000000,
465.000000000000,-310.000000000000,
1185.00000000000,-434.000000000000,
38.0000000000000,297.000000000000,
-1116.00000000000,249.000000000000,
-805.000000000000,-716.000000000000,
-119.000000000000,-6.00000000000000,
-1444.00000000000,313.000000000000,
175.000000000000,161.000000000000,
938.000000000000,376.000000000000,
-112.000000000000,79.0000000000000,
-257.000000000000,-320.000000000000,
-371.000000000000,123.000000000000,
258.000000000000,-586.000000000000,
480.000000000000,-629.000000000000,
1171.00000000000,-103.000000000000,
746.000000000000,-609.000000000000,
330.000000000000,-332.000000000000,
904.000000000000,-479.000000000000,
638.000000000000,-141.000000000000,
460.000000000000,-911.000000000000,
50.0000000000000,-322.000000000000,
406.000000000000,173.000000000000,
-598.000000000000,-972.000000000000,
73.0000000000000,1104.00000000000,
386.000000000000,578.000000000000,
-1306.00000000000,223.000000000000,
362.000000000000,-452.000000000000,
765.000000000000,-715.000000000000,
1044.00000000000,253.000000000000,
408.000000000000,229.000000000000,
-28.0000000000000,1350.00000000000,
24.0000000000000,-521.000000000000,
-1036.00000000000,-279.000000000000,
-349.000000000000,-561.000000000000,
88.0000000000000,-1271.00000000000,
1226.00000000000,-235.000000000000,
555.000000000000,-151.000000000000,
-312.000000000000,850.000000000000,
-366.000000000000,604.000000000000,
-229.000000000000,121.000000000000,
661.000000000000,-972.000000000000,
325.000000000000,258.000000000000,
633.000000000000,1697.00000000000,
-332.000000000000,822.000000000000,
-988.000000000000,460.000000000000,
72.0000000000000,-302.000000000000,
-26.0000000000000,391.000000000000,
-445.000000000000,108.000000000000,
-61.0000000000000,242.000000000000,
537.000000000000,681.000000000000,
-404.000000000000,15.0000000000000,
-427.000000000000,-167.000000000000,
33.0000000000000,-1507.00000000000,
-520.000000000000,-1200.00000000000,
431.000000000000,-261.000000000000,
366.000000000000,495.000000000000,
-114.000000000000,-148.000000000000,
577.000000000000,-118.000000000000,
98.0000000000000,-115.000000000000,
-26.0000000000000,-821.000000000000,
1226.00000000000,1451.00000000000,
-356.000000000000,985.000000000000,
-1198.00000000000,-79.0000000000000,
1188.00000000000,-408.000000000000,
-301.000000000000,-718.000000000000,
-771.000000000000,854.000000000000,
-613.000000000000,101.000000000000,
-1329.00000000000,-99.0000000000000,
285.000000000000,-206.000000000000,
804.000000000000,-483.000000000000,
743.000000000000,-60.0000000000000,
-920.000000000000,441.000000000000,
89.0000000000000,674.000000000000,
383.000000000000,301.000000000000,
-59.0000000000000,946.000000000000,
388.000000000000,-948.000000000000,
-1030.00000000000,-339.000000000000,
-102.000000000000,947.000000000000,
-163.000000000000,290.000000000000,
643.000000000000,1186.00000000000,
-748.000000000000,357.000000000000,
-1032.00000000000,-304.000000000000,
913.000000000000,-1107.00000000000,
-301.000000000000,273.000000000000,
-528.000000000000,1179.00000000000,
-767.000000000000,-391.000000000000,
938.000000000000,-135.000000000000,
459.000000000000,-141.000000000000,
-597.000000000000,-399.000000000000,
48.0000000000000,-547.000000000000,
-26.0000000000000,59.0000000000000,
438.000000000000,259.000000000000,
-853.000000000000,209.000000000000,
-608.000000000000,70.0000000000000,
176.000000000000,-222.000000000000,
822.000000000000,-132.000000000000,
332.000000000000,-870.000000000000,
-440.000000000000,-655.000000000000,
305.000000000000,-352.000000000000,
-426.000000000000,292.000000000000,
-457.000000000000,1015.00000000000,
-658.000000000000,-127.000000000000,
-750.000000000000,-576.000000000000,
246.000000000000,-232.000000000000,
-111.000000000000,181.000000000000,
-379.000000000000,-461.000000000000,
-569.000000000000,-104.000000000000,
-755.000000000000,277.000000000000,
-1231.00000000000,-331.000000000000,
-607.000000000000,-31.0000000000000,
-861.000000000000,-577.000000000000,
-152.000000000000,204.000000000000,
992.000000000000,-488.000000000000,
-604.000000000000,-491.000000000000,
480.000000000000,-155.000000000000,
849.000000000000,-1087.00000000000,
1090.00000000000,699.000000000000,
87.0000000000000,531.000000000000,
-1045.00000000000,533.000000000000,
711.000000000000,593.000000000000,
-506.000000000000,574.000000000000,
-582.000000000000,606.000000000000,
-878.000000000000,-513.000000000000,
-688.000000000000,384.000000000000,
-948.000000000000,-198.000000000000,
-538.000000000000,-873.000000000000,
879.000000000000,159.000000000000,
-384.000000000000,654.000000000000,
615.000000000000,724.000000000000,
-84.0000000000000,1068.00000000000,
-887.000000000000,625.000000000000,
787.000000000000,-837.000000000000,
182.000000000000,-525.000000000000,
-612.000000000000,455.000000000000,
553.000000000000,-532.000000000000,
473.000000000000,82.0000000000000,
14.0000000000000,1277.00000000000,
-394.000000000000,-104.000000000000,
-1370.00000000000,-367.000000000000,
-257.000000000000,-634.000000000000,
177.000000000000,-377.000000000000,
37.0000000000000,-26.0000000000000,
832.000000000000,-425.000000000000,
536.000000000000,682.000000000000,
621.000000000000,1208.00000000000,
348.000000000000,-66.0000000000000,
438.000000000000,-191.000000000000,
624.000000000000,145.000000000000,
-672.000000000000,655.000000000000,
-267.000000000000,-35.0000000000000,
505.000000000000,-943.000000000000,
1211.00000000000,222.000000000000,
487.000000000000,294.000000000000,
224.000000000000,1178.00000000000,
43.0000000000000,1180.00000000000,
-1675.00000000000,-375.000000000000,
129.000000000000,-839.000000000000,
1036.00000000000,-819.000000000000,
49.0000000000000,-354.000000000000,
-634.000000000000,-441.000000000000,
831.000000000000,-483.000000000000,
727.000000000000,-399.000000000000,
-1319.00000000000,644.000000000000,
-452.000000000000,-386.000000000000,
155.000000000000,-1043.00000000000,
1469.00000000000,17.0000000000000,
1006.00000000000,-322.000000000000,
496.000000000000,404.000000000000,
159.000000000000,-260.000000000000,
-975.000000000000,509.000000000000,
-497.000000000000,305.000000000000,
-1111.00000000000,-957.000000000000,
995.000000000000,194.000000000000,
244.000000000000,655.000000000000,
-957.000000000000,1112.00000000000,
-55.0000000000000,128.000000000000,
-1465.00000000000,111.000000000000,
407.000000000000,-313.000000000000,
1062.00000000000,-676.000000000000,
-342.000000000000,556.000000000000,
258.000000000000,667.000000000000,
-295.000000000000,901.000000000000,
-792.000000000000,488.000000000000,
-249.000000000000,-197.000000000000,
-207.000000000000,-1327.00000000000,
-458.000000000000,427.000000000000,
1.00000000000000,349.000000000000,
791.000000000000,-403.000000000000,
-60.0000000000000,531.000000000000,
-142.000000000000,-779.000000000000,
561.000000000000,1105.00000000000,
557.000000000000,643.000000000000,
96.0000000000000,119.000000000000,
-648.000000000000,-136.000000000000,
297.000000000000,-1162.00000000000,
606.000000000000,846.000000000000,
66.0000000000000,672.000000000000,
-1063.00000000000,798.000000000000,
-1065.00000000000,241.000000000000,
-193.000000000000,669.000000000000,
-178.000000000000,-435.000000000000,
-310.000000000000,-1111.00000000000,
-291.000000000000,166.000000000000,
-358.000000000000,-1629.00000000000,
-244.000000000000,269.000000000000,
-87.0000000000000,111.000000000000,
-133.000000000000,-1379.00000000000,
1232.00000000000,540.000000000000,
587.000000000000,496.000000000000,
-208.000000000000,-844.000000000000,
38.0000000000000,-1335.00000000000,
-455.000000000000,-112.000000000000,
-343.000000000000,-557.000000000000,
-850.000000000000,-105.000000000000,
-305.000000000000,984.000000000000,
445.000000000000,462.000000000000,
-337.000000000000,-160.000000000000,
-437.000000000000,0.00000000000000,
72.0000000000000,189.000000000000,
326.000000000000,-1047.00000000000,
-221.000000000000,9.00000000000000,
-684.000000000000,-347.000000000000,
773.000000000000,-1026.00000000000,
1616.00000000000,477.000000000000,
-579.000000000000,276.000000000000,
-779.000000000000,-19.0000000000000,
431.000000000000,-1153.00000000000,
325.000000000000,-432.000000000000,
1482.00000000000,-295.000000000000,
767.000000000000,331.000000000000,
363.000000000000,1770.00000000000,
523.000000000000,-131.000000000000,
-18.0000000000000,194.000000000000,
104.000000000000,584.000000000000,
-260.000000000000,366.000000000000,
218.000000000000,633.000000000000,
-263.000000000000,-463.000000000000,
697.000000000000,27.0000000000000,
778.000000000000,791.000000000000,
-549.000000000000,717.000000000000,
-1212.00000000000,-118.000000000000,
-526.000000000000,-1064.00000000000,
734.000000000000,125.000000000000,
-46.0000000000000,1505.00000000000,
197.000000000000,1098.00000000000,
-309.000000000000,159.000000000000,
-452.000000000000,-490.000000000000,
-572.000000000000,-718.000000000000,
-601.000000000000,-500.000000000000,
838.000000000000,-184.000000000000,
436.000000000000,820.000000000000,
511.000000000000,648.000000000000,
242.000000000000,37.0000000000000,
-200.000000000000,997.000000000000,
-201.000000000000,335.000000000000,
153.000000000000,-15.0000000000000,
1154.00000000000,-92.0000000000000,
493.000000000000,568.000000000000,
205.000000000000,1131.00000000000,
-1340.00000000000,-103.000000000000,
-513.000000000000,237.000000000000,
1281.00000000000,-489.000000000000,
435.000000000000,654.000000000000,
800.000000000000,481.000000000000,
-324.000000000000,-666.000000000000,
-560.000000000000,-157.000000000000,
-1067.00000000000,-998.000000000000,
520.000000000000,-302.000000000000,
1316.00000000000,-605.000000000000,
-19.0000000000000,-594.000000000000,
370.000000000000,148.000000000000,
97.0000000000000,199.000000000000,
620.000000000000,358.000000000000,
-891.000000000000,146.000000000000,
335.000000000000,219.000000000000,
897.000000000000,-791.000000000000,
-515.000000000000,-873.000000000000,
615.000000000000,580.000000000000,
-259.000000000000,719.000000000000,
-585.000000000000,-621.000000000000,
-74.0000000000000,-554.000000000000,
-201.000000000000,55.0000000000000,
-1368.00000000000,-513.000000000000,
-403.000000000000,392.000000000000,
57.0000000000000,481.000000000000,
-569.000000000000,155.000000000000,
1378.00000000000,-15.0000000000000,
-369.000000000000,-802.000000000000,
493.000000000000,637.000000000000,
743.000000000000,548.000000000000,
528.000000000000,181.000000000000,
987.000000000000,-336.000000000000,
-1206.00000000000,207.000000000000,
959.000000000000,435.000000000000,
69.0000000000000,-803.000000000000,
417.000000000000,571.000000000000,
-458.000000000000,260.000000000000,
-761.000000000000,-258.000000000000,
1234.00000000000,-723.000000000000,
-1468.00000000000,202.000000000000,
-420.000000000000,-412.000000000000,
-311.000000000000,-848.000000000000,
-92.0000000000000,584.000000000000,
732.000000000000,-926.000000000000,
889.000000000000,-190.000000000000,
1453.00000000000,-292.000000000000,
1079.00000000000,-21.0000000000000,
1050.00000000000,1137.00000000000,
-629.000000000000,994.000000000000,
-1118.00000000000,92.0000000000000,
-662.000000000000,-1471.00000000000,
256.000000000000,-251.000000000000,
677.000000000000,249.000000000000,
540.000000000000,-173.000000000000,
1172.00000000000,618.000000000000,
-35.0000000000000,1591.00000000000,
360.000000000000,751.000000000000,
194.000000000000,-272.000000000000,
-767.000000000000,521.000000000000,
-71.0000000000000,50.0000000000000,
301.000000000000,847.000000000000,
401.000000000000,308.000000000000,
-237.000000000000,90.0000000000000,
309.000000000000,1533.00000000000,
-334.000000000000,531.000000000000,
-342.000000000000,-211.000000000000,
87.0000000000000,-615.000000000000,
-75.0000000000000,892.000000000000,
468.000000000000,-38.0000000000000,
77.0000000000000,-842.000000000000,
1207.00000000000,212.000000000000,
-272.000000000000,-548.000000000000,
-83.0000000000000,539.000000000000,
1205.00000000000,276.000000000000,
-389.000000000000,-464.000000000000,
780.000000000000,-424.000000000000,
371.000000000000,738.000000000000,
-801.000000000000,1028.00000000000,
-311.000000000000,-159.000000000000,
640.000000000000,185.000000000000,
245.000000000000,-106.000000000000,
-41.0000000000000,963.000000000000,
-252.000000000000,22.0000000000000,
-658.000000000000,-1526.00000000000,
788.000000000000,228.000000000000,
-735.000000000000,350.000000000000,
339.000000000000,-498.000000000000,
1550.00000000000,-148.000000000000,
559.000000000000,729.000000000000,
396.000000000000,607.000000000000,
-913.000000000000,17.0000000000000,
333.000000000000,858.000000000000,
-69.0000000000000,729.000000000000,
-897.000000000000,115.000000000000,
-257.000000000000,253.000000000000,
-631.000000000000,-262.000000000000,
-615.000000000000,194.000000000000,
150.000000000000,481.000000000000,
-68.0000000000000,178.000000000000,
-204.000000000000,-188.000000000000,
-226.000000000000,-619.000000000000,
-1081.00000000000,122.000000000000,
-431.000000000000,-709.000000000000,
841.000000000000,-424.000000000000,
857.000000000000,-258.000000000000,
-133.000000000000,145.000000000000,
316.000000000000,341.000000000000,
-125.000000000000,-1038.00000000000,
256.000000000000,-215.000000000000,
696.000000000000,24.0000000000000,
-1350.00000000000,27.0000000000000,
-948.000000000000,124.000000000000,
127.000000000000,-737.000000000000,
-293.000000000000,-715.000000000000,
743.000000000000,-99.0000000000000,
967.000000000000,823.000000000000,
-475.000000000000,1165.00000000000,
-949.000000000000,-760.000000000000,
121.000000000000,-325.000000000000,
359.000000000000,1303.00000000000,
-965.000000000000,-306.000000000000,
684.000000000000,-988.000000000000,
685.000000000000,-432.000000000000,
-652.000000000000,411.000000000000,
501.000000000000,520.000000000000,
286.000000000000,-514.000000000000,
-48.0000000000000,-83.0000000000000,
-757.000000000000,978.000000000000,
-848.000000000000,332.000000000000,
-649.000000000000,190.000000000000,
-659.000000000000,746.000000000000,
646.000000000000,-764.000000000000,
25.0000000000000,-102.000000000000,
-88.0000000000000,-841.000000000000,
199.000000000000,-467.000000000000,
-825.000000000000,1182.00000000000,
-562.000000000000,98.0000000000000,
-392.000000000000,62.0000000000000,
565.000000000000,-991.000000000000,
982.000000000000,230.000000000000,
-599.000000000000,-638.000000000000,
80.0000000000000,-1698.00000000000,
1669.00000000000,240.000000000000,
-223.000000000000,188.000000000000,
-428.000000000000,592.000000000000,
302.000000000000,65.0000000000000,
-477.000000000000,-42.0000000000000,
864.000000000000,-363.000000000000,
425.000000000000,-625.000000000000,
671.000000000000,-196.000000000000,
993.000000000000,146.000000000000,
-1061.00000000000,844.000000000000,
-794.000000000000,382.000000000000,
90.0000000000000,882.000000000000,
-506.000000000000,821.000000000000,
-887.000000000000,176.000000000000,
-469.000000000000,-434.000000000000,
64.0000000000000,-498.000000000000,
298.000000000000,-287.000000000000,
217.000000000000,-655.000000000000,
-540.000000000000,528.000000000000,
-531.000000000000,554.000000000000,
-21.0000000000000,-446.000000000000,
-234.000000000000,-509.000000000000,
723.000000000000,-38.0000000000000,
434.000000000000,299.000000000000,
-375.000000000000,196.000000000000,
-645.000000000000,521.000000000000,
-1002.00000000000,445.000000000000,
-294.000000000000,-519.000000000000,
275.000000000000,-581.000000000000,
690.000000000000,578.000000000000,
-572.000000000000,-108.000000000000,
-496.000000000000,540.000000000000,
-605.000000000000,675.000000000000,
-404.000000000000,-1485.00000000000,
662.000000000000,286.000000000000,
-587.000000000000,501.000000000000,
181.000000000000,-298.000000000000,
-253.000000000000,442.000000000000,
-734.000000000000,-338.000000000000,
-679.000000000000,260.000000000000,
-179.000000000000,313.000000000000,
595.000000000000,291.000000000000,
-694.000000000000,-303.000000000000,
-986.000000000000,143.000000000000,
-872.000000000000,28.0000000000000,
-158.000000000000,-1671.00000000000,
1533.00000000000,14.0000000000000,
906.000000000000,-564.000000000000,
-893.000000000000,-28.0000000000000,
334.000000000000,581.000000000000,
-522.000000000000,-575.000000000000,
112.000000000000,1015.00000000000,
186.000000000000,369.000000000000,
-1079.00000000000,467.000000000000,
161.000000000000,-195.000000000000,
135.000000000000,-574.000000000000,
134.000000000000,519.000000000000,
-1046.00000000000,12.0000000000000,
692.000000000000,-1022.00000000000,
1403.00000000000,-242.000000000000,
-146.000000000000,1335.00000000000,
318.000000000000,-799.000000000000,
-433.000000000000,-59.0000000000000,
-477.000000000000,-252.000000000000,
107.000000000000,-1508.00000000000,
940.000000000000,281.000000000000,
-276.000000000000,-571.000000000000,
180.000000000000,331.000000000000,
233.000000000000,802.000000000000,
-833.000000000000,-68.0000000000000,
1425.00000000000,-441.000000000000,
944.000000000000,-51.0000000000000,
1278.00000000000,361.000000000000,
783.000000000000,-236.000000000000,
87.0000000000000,1607.00000000000,
-197.000000000000,965.000000000000,
-1166.00000000000,-1156.00000000000,
-60.0000000000000,-296.000000000000,
-795.000000000000,-208.000000000000,
-542.000000000000,-741.000000000000,
-109.000000000000,-177.000000000000,
-171.000000000000,-225.000000000000,
81.0000000000000,-814.000000000000,
754.000000000000,451.000000000000,
374.000000000000,787.000000000000,
-1190.00000000000,-132.000000000000,
14.0000000000000,-885.000000000000,
439.000000000000,-657.000000000000,
565.000000000000,-5.00000000000000,
885.000000000000,-790.000000000000,
-222.000000000000,-439.000000000000,
171.000000000000,-831.000000000000,
1038.00000000000,-375.000000000000,
622.000000000000,1113.00000000000,
-218.000000000000,1084.00000000000,
-375.000000000000,612.000000000000,
-88.0000000000000,-232.000000000000,
-168.000000000000,986.000000000000,
-597.000000000000,618.000000000000,
-1484.00000000000,-347.000000000000,
-239.000000000000,-318.000000000000,
900.000000000000,-374.000000000000,
270.000000000000,-587.000000000000,
972.000000000000,-695.000000000000,
220.000000000000,1238.00000000000,
-930.000000000000,506.000000000000,
-100.000000000000,286.000000000000,
449.000000000000,-16.0000000000000,
593.000000000000,-391.000000000000,
1012.00000000000,424.000000000000,
451.000000000000,-134.000000000000,
163.000000000000,1206.00000000000,
817.000000000000,285.000000000000,
192.000000000000,-399.000000000000,
-6.00000000000000,-192.000000000000,
-406.000000000000,-1246.00000000000,
-722.000000000000,-73.0000000000000,
-264.000000000000,110.000000000000,
1108.00000000000,-24.0000000000000,
861.000000000000,-319.000000000000,
-686.000000000000,-564.000000000000,
870.000000000000,-246.000000000000,
158.000000000000,-453.000000000000,
111.000000000000,-58.0000000000000,
-364.000000000000,343.000000000000,
-182.000000000000,411.000000000000,
294.000000000000,-1116.00000000000,
-889.000000000000,21.0000000000000,
390.000000000000,442.000000000000,
-794.000000000000,-804.000000000000,
187.000000000000,-31.0000000000000,
-56.0000000000000,-1018.00000000000,
-348.000000000000,-310.000000000000,
1943.00000000000,-246.000000000000,
532.000000000000,275.000000000000,
847.000000000000,-224.000000000000,
215.000000000000,-2.00000000000000,
-220.000000000000,578.000000000000,
599.000000000000,-1045.00000000000,
621.000000000000,800.000000000000,
191.000000000000,-32.0000000000000,
-549.000000000000,-324.000000000000,
324.000000000000,-370.000000000000,
-224.000000000000,-48.0000000000000,
158.000000000000,1126.00000000000,
24.0000000000000,176.000000000000,
-1166.00000000000,965.000000000000,
-230.000000000000,-261.000000000000,
200.000000000000,-238.000000000000,
171.000000000000,-38.0000000000000,
23.0000000000000,-67.0000000000000,
154.000000000000,-466.000000000000,
426.000000000000,-703.000000000000,
548.000000000000,839.000000000000,
646.000000000000,671.000000000000,
178.000000000000,415.000000000000,
-183.000000000000,539.000000000000,
354.000000000000,110.000000000000,
-241.000000000000,445.000000000000,
-792.000000000000,-142.000000000000,
-644.000000000000,-1093.00000000000,
-30.0000000000000,69.0000000000000,
948.000000000000,104.000000000000,
533.000000000000,848.000000000000,
-131.000000000000,1250.00000000000,
-534.000000000000,-403.000000000000,
122.000000000000,-166.000000000000,
905.000000000000,47.0000000000000,
1.00000000000000,-309.000000000000,
-91.0000000000000,166.000000000000,
496.000000000000,-244.000000000000,
-3.00000000000000,1045.00000000000,
50.0000000000000,809.000000000000,
-925.000000000000,-264.000000000000,
-503.000000000000,561.000000000000,
192.000000000000,-366.000000000000,
-647.000000000000,561.000000000000,
874.000000000000,122.000000000000,
518.000000000000,-597.000000000000,
-319.000000000000,-35.0000000000000,
-96.0000000000000,-304.000000000000,
-518.000000000000,-434.000000000000,
364.000000000000,-400.000000000000,
317.000000000000,1424.00000000000,
318.000000000000,-356.000000000000,
150.000000000000,-424.000000000000,
161.000000000000,490.000000000000,
262.000000000000,346.000000000000,
-190.000000000000,854.000000000000,
-1155.00000000000,-478.000000000000,
-125.000000000000,475.000000000000,
698.000000000000,-476.000000000000,
-658.000000000000,-524.000000000000,
156.000000000000,746.000000000000,
-678.000000000000,248.000000000000,
209.000000000000,414.000000000000,
551.000000000000,-998.000000000000,
-1193.00000000000,-961.000000000000,
666.000000000000,-603.000000000000,
1114.00000000000,-524.000000000000,
-506.000000000000,493.000000000000,
-436.000000000000,-22.0000000000000,
205.000000000000,-419.000000000000,
-189.000000000000,596.000000000000,
-478.000000000000,130.000000000000,
-997.000000000000,-101.000000000000,
-617.000000000000,-324.000000000000,
227.000000000000,-635.000000000000,
-664.000000000000,662.000000000000,
-799.000000000000,-39.0000000000000,
345.000000000000,-771.000000000000,
1098.00000000000,976.000000000000,
-14.0000000000000,133.000000000000,
-1024.00000000000,-305.000000000000,
-930.000000000000,8.00000000000000,
-728.000000000000,-1082.00000000000,
1273.00000000000,-364.000000000000,
-118.000000000000,121.000000000000,
-1376.00000000000,179.000000000000,
-172.000000000000,350.000000000000,
-217.000000000000,1278.00000000000,
278.000000000000,328.000000000000,
-1085.00000000000,-561.000000000000,
-752.000000000000,648.000000000000,
-193.000000000000,24.0000000000000,
-772.000000000000,-371.000000000000,
-770.000000000000,-138.000000000000,
-398.000000000000,22.0000000000000,
531.000000000000,93.0000000000000,
-131.000000000000,117.000000000000,
-532.000000000000,321.000000000000,
-104.000000000000,-14.0000000000000,
36.0000000000000,176.000000000000,
-395.000000000000,443.000000000000,
129.000000000000,653.000000000000,
511.000000000000,-171.000000000000,
-458.000000000000,-78.0000000000000,
219.000000000000,995.000000000000,
-826.000000000000,199.000000000000,
244.000000000000,285.000000000000,
455.000000000000,-128.000000000000,
-803.000000000000,-195.000000000000,
57.0000000000000,-547.000000000000,
-538.000000000000,-1357.00000000000,
569.000000000000,-224.000000000000,
18.0000000000000,94.0000000000000,
98.0000000000000,181.000000000000,
789.000000000000,709.000000000000,
-614.000000000000,971.000000000000,
-314.000000000000,462.000000000000,
-500.000000000000,105.000000000000,
243.000000000000,-548.000000000000,
868.000000000000,122.000000000000,
-164.000000000000,656.000000000000,
-118.000000000000,-826.000000000000,
474.000000000000,1134.00000000000,
-91.0000000000000,1170.00000000000,
-1191.00000000000,-448.000000000000,
-710.000000000000,-158.000000000000,
-293.000000000000,-152.000000000000,
-610.000000000000,-564.000000000000,
473.000000000000,-294.000000000000,
-488.000000000000,805.000000000000,
-926.000000000000,69.0000000000000,
702.000000000000,324.000000000000,
643.000000000000,-839.000000000000,
293.000000000000,-144.000000000000,
520.000000000000,1161.00000000000,
-1147.00000000000,-590.000000000000,
-628.000000000000,779.000000000000,
555.000000000000,221.000000000000,
-832.000000000000,241.000000000000,
487.000000000000,626.000000000000,
233.000000000000,-1020.00000000000,
185.000000000000,165.000000000000,
1602.00000000000,-464.000000000000,
258.000000000000,-422.000000000000,
-741.000000000000,524.000000000000,
-628.000000000000,-1027.00000000000,
78.0000000000000,-387.000000000000,
194.000000000000,1210.00000000000,
384.000000000000,-855.000000000000,
485.000000000000,-313.000000000000,
251.000000000000,1565.00000000000,
412.000000000000,-754.000000000000,
38.0000000000000,1.00000000000000,
-119.000000000000,527.000000000000,
-395.000000000000,226.000000000000,
-420.000000000000,635.000000000000,
1006.00000000000,-523.000000000000,
436.000000000000,21.0000000000000,
-551.000000000000,-586.000000000000,
-75.0000000000000,-1271.00000000000,
162.000000000000,-674.000000000000,
545.000000000000,98.0000000000000,
967.000000000000,-386.000000000000,
-521.000000000000,-4.00000000000000,
-163.000000000000,1145.00000000000,
665.000000000000,-765.000000000000,
405.000000000000,551.000000000000,
1238.00000000000,224.000000000000,
-693.000000000000,-706.000000000000,
-81.0000000000000,951.000000000000,
-224.000000000000,-959.000000000000,
-588.000000000000,330.000000000000,
18.0000000000000,797.000000000000,
-903.000000000000,-1001.00000000000,
970.000000000000,-758.000000000000,
1028.00000000000,28.0000000000000,
1123.00000000000,231.000000000000,
413.000000000000,-634.000000000000,
260.000000000000,-109.000000000000,
258.000000000000,-30.0000000000000,
-323.000000000000,192.000000000000,
-683.000000000000,426.000000000000,
-1147.00000000000,-404.000000000000,
1092.00000000000,188.000000000000,
575.000000000000,560.000000000000,
-436.000000000000,-494.000000000000,
317.000000000000,-1203.00000000000,
949.000000000000,-434.000000000000,
183.000000000000,-24.0000000000000,
235.000000000000,-398.000000000000,
1550.00000000000,134.000000000000,
-392.000000000000,-586.000000000000,
590.000000000000,-338.000000000000,
445.000000000000,-106.000000000000,
-336.000000000000,-496.000000000000,
512.000000000000,856.000000000000,
-1085.00000000000,-316.000000000000,
19.0000000000000,-1299.00000000000,
-286.000000000000,64.0000000000000,
-784.000000000000,69.0000000000000,
-15.0000000000000,-720.000000000000,
291.000000000000,1128.00000000000,
-262.000000000000,632.000000000000,
-409.000000000000,-1163.00000000000,
871.000000000000,263.000000000000,
-191.000000000000,856.000000000000,
608.000000000000,936.000000000000,
-643.000000000000,29.0000000000000,
-420.000000000000,-313.000000000000,
767.000000000000,-666.000000000000,
-349.000000000000,-1416.00000000000,
1386.00000000000,346.000000000000,
75.0000000000000,-531.000000000000,
87.0000000000000,-373.000000000000,
497.000000000000,683.000000000000,
291.000000000000,-450.000000000000,
-116.000000000000,-28.0000000000000,
-515.000000000000,-965.000000000000,
-130.000000000000,-529.000000000000,
-842.000000000000,260.000000000000,
900.000000000000,-688.000000000000,
-420.000000000000,-613.000000000000,
-343.000000000000,545.000000000000,
232.000000000000,709.000000000000,
-1462.00000000000,441.000000000000,
1000.00000000000,139.000000000000,
702.000000000000,-184.000000000000,
-142.000000000000,921.000000000000,
283.000000000000,800.000000000000,
-109.000000000000,368.000000000000,
402.000000000000,-286.000000000000,
126.000000000000,89.0000000000000,
-483.000000000000,-179.000000000000,
-632.000000000000,434.000000000000,
213.000000000000,884.000000000000,
-199.000000000000,160.000000000000,
-102.000000000000,1559.00000000000,
-96.0000000000000,-290.000000000000,
-1192.00000000000,-479.000000000000,
159.000000000000,-413.000000000000,
245.000000000000,-1266.00000000000,
290.000000000000,-170.000000000000,
264.000000000000,-1318.00000000000,
256.000000000000,-314.000000000000,
-225.000000000000,367.000000000000,
-277.000000000000,-416.000000000000,
782.000000000000,-233.000000000000,
-400.000000000000,133.000000000000,
508.000000000000,932.000000000000,
-207.000000000000,936.000000000000,
-812.000000000000,525.000000000000,
363.000000000000,-254.000000000000,
-269.000000000000,-171.000000000000,
-698.000000000000,-203.000000000000,
-574.000000000000,167.000000000000,
1158.00000000000,-307.000000000000,
638.000000000000,150.000000000000,
-455.000000000000,1427.00000000000,
9.00000000000000,-857.000000000000,
-156.000000000000,-153.000000000000,
-59.0000000000000,747.000000000000,
-213.000000000000,611.000000000000,
647.000000000000,130.000000000000,
-66.0000000000000,-794.000000000000,
-800.000000000000,685.000000000000,
133.000000000000,80.0000000000000,
-555.000000000000,-298.000000000000,
-200.000000000000,-310.000000000000,
-211.000000000000,557.000000000000,
-373.000000000000,615.000000000000,
647.000000000000,-274.000000000000,
386.000000000000,-335.000000000000,
-6.00000000000000,-998.000000000000,
38.0000000000000,-234.000000000000,
-268.000000000000,-148.000000000000,
-1234.00000000000,344.000000000000,
-762.000000000000,-469.000000000000,
1075.00000000000,-935.000000000000,
1148.00000000000,530.000000000000,
86.0000000000000,105.000000000000,
-135.000000000000,-401.000000000000,
93.0000000000000,421.000000000000,
-546.000000000000,1177.00000000000,
-475.000000000000,-365.000000000000,
471.000000000000,-37.0000000000000,
-80.0000000000000,1177.00000000000,
-908.000000000000,-587.000000000000,
142.000000000000,-371.000000000000,
1507.00000000000,222.000000000000,
701.000000000000,-293.000000000000,
179.000000000000,8.00000000000000,
-126.000000000000,-142.000000000000,
-377.000000000000,-923.000000000000,
750.000000000000,-354.000000000000,
958.000000000000,308.000000000000,
372.000000000000,-600.000000000000,
452.000000000000,-106.000000000000,
449.000000000000,-16.0000000000000,
481.000000000000,-432.000000000000,
744.000000000000,1071.00000000000,
-291.000000000000,955.000000000000,
-53.0000000000000,-38.0000000000000,
551.000000000000,187.000000000000,
355.000000000000,416.000000000000,
79.0000000000000,859.000000000000,
-841.000000000000,686.000000000000,
-225.000000000000,717.000000000000,
-162.000000000000,682.000000000000,
-139.000000000000,-346.000000000000,
-560.000000000000,-1341.00000000000,
-2.00000000000000,-662.000000000000,
530.000000000000,813.000000000000,
-1251.00000000000,-351.000000000000,
913.000000000000,-370.000000000000,
1014.00000000000,877.000000000000,
-862.000000000000,516.000000000000,
-10.0000000000000,-719.000000000000,
369.000000000000,-709.000000000000,
1386.00000000000,-175.000000000000,
615.000000000000,735.000000000000,
-587.000000000000,-21.0000000000000,
-286.000000000000,-1214.00000000000,
-263.000000000000,918.000000000000,
-307.000000000000,776.000000000000,
49.0000000000000,616.000000000000,
361.000000000000,-443.000000000000,
-888.000000000000,-268.000000000000,
-267.000000000000,907.000000000000,
-106.000000000000,231.000000000000,
265.000000000000,447.000000000000,
451.000000000000,-386.000000000000,
-727.000000000000,783.000000000000,
488.000000000000,-131.000000000000,
-497.000000000000,-598.000000000000,
-1259.00000000000,705.000000000000,
-177.000000000000,-1045.00000000000,
-515.000000000000,-1118.00000000000,
110.000000000000,380.000000000000,
-355.000000000000,837.000000000000,
-405.000000000000,-108.000000000000,
780.000000000000,-234.000000000000,
13.0000000000000,-324.000000000000,
99.0000000000000,387.000000000000,
42.0000000000000,139.000000000000,
-939.000000000000,-756.000000000000,
-707.000000000000,351.000000000000,
-673.000000000000,-1013.00000000000,
-530.000000000000,-815.000000000000,
1240.00000000000,-192.000000000000,
662.000000000000,-285.000000000000,
-418.000000000000,1011.00000000000,
-543.000000000000,-617.000000000000,
-384.000000000000,46.0000000000000,
112.000000000000,1043.00000000000,
-887.000000000000,-266.000000000000,
121.000000000000,-447.000000000000,
576.000000000000,-353.000000000000,
1006.00000000000,83.0000000000000,
-246.000000000000,-1023.00000000000,
23.0000000000000,-516.000000000000,
544.000000000000,257.000000000000,
-527.000000000000,-310.000000000000,
1678.00000000000,-375.000000000000,
-131.000000000000,-56.0000000000000,
56.0000000000000,1313.00000000000,
-298.000000000000,64.0000000000000,
-478.000000000000,148.000000000000,
971.000000000000,-190.000000000000,
-1038.00000000000,-488.000000000000,
-642.000000000000,526.000000000000,
-959.000000000000,-585.000000000000,
932.000000000000,1.00000000000000,
446.000000000000,-323.000000000000,
-1062.00000000000,-848.000000000000,
587.000000000000,-559.000000000000,
485.000000000000,-249.000000000000,
81.0000000000000,318.000000000000,
-520.000000000000,449.000000000000,
-86.0000000000000,453.000000000000,
-430.000000000000,-195.000000000000,
319.000000000000,-451.000000000000,
-13.0000000000000,-922.000000000000,
-449.000000000000,-392.000000000000,
230.000000000000,544.000000000000,
-1434.00000000000,52.0000000000000,
-1016.00000000000,-476.000000000000,
386.000000000000,-1388.00000000000,
1351.00000000000,10.0000000000000,
635.000000000000,1095.00000000000,
789.000000000000,-64.0000000000000,
805.000000000000,662.000000000000,
-1230.00000000000,142.000000000000,
718.000000000000,-554.000000000000,
569.000000000000,-666.000000000000,
564.000000000000,660.000000000000,
-47.0000000000000,1043.00000000000,
-1268.00000000000,-978.000000000000,
555.000000000000,-846.000000000000,
-144.000000000000,594.000000000000,
110.000000000000,946.000000000000,
-312.000000000000,-133.000000000000,
-417.000000000000,556.000000000000,
119.000000000000,446.000000000000,
38.0000000000000,-86.0000000000000,
-316.000000000000,115.000000000000,
-514.000000000000,-624.000000000000,
1430.00000000000,-164.000000000000,
164.000000000000,-588.000000000000,
557.000000000000,-63.0000000000000,
-207.000000000000,405.000000000000,
-1028.00000000000,237.000000000000,
1022.00000000000,90.0000000000000,
445.000000000000,-578.000000000000,
820.000000000000,1046.00000000000,
411.000000000000,1381.00000000000,
-620.000000000000,-550.000000000000,
-255.000000000000,43.0000000000000,
249.000000000000,713.000000000000,
257.000000000000,-895.000000000000,
-984.000000000000,215.000000000000,
-494.000000000000,-126.000000000000,
-191.000000000000,-1677.00000000000,
-224.000000000000,-571.000000000000,
1011.00000000000,-754.000000000000,
207.000000000000,93.0000000000000,
-335.000000000000,-571.000000000000,
852.000000000000,-502.000000000000,
1372.00000000000,388.000000000000,
192.000000000000,320.000000000000,
411.000000000000,318.000000000000,
342.000000000000,-1039.00000000000,
-839.000000000000,661.000000000000,
152.000000000000,679.000000000000,
202.000000000000,-398.000000000000,
155.000000000000,585.000000000000,
-432.000000000000,1018.00000000000,
-792.000000000000,6.00000000000000,
15.0000000000000,-1365.00000000000,
479.000000000000,-792.000000000000,
365.000000000000,-551.000000000000,
-244.000000000000,479.000000000000,
-71.0000000000000,872.000000000000,
-440.000000000000,-1.00000000000000,
-557.000000000000,-673.000000000000,
641.000000000000,-116.000000000000,
-92.0000000000000,1112.00000000000,
10.0000000000000,-154.000000000000,
801.000000000000,487.000000000000,
-547.000000000000,957.000000000000,
-1298.00000000000,-103.000000000000,
-746.000000000000,-146.000000000000,
-67.0000000000000,-15.0000000000000,
633.000000000000,518.000000000000,
462.000000000000,764.000000000000,
-284.000000000000,933.000000000000,
-124.000000000000,555.000000000000,
-61.0000000000000,-588.000000000000,
-122.000000000000,-1117.00000000000,
699.000000000000,-749.000000000000,
1372.00000000000,343.000000000000,
46.0000000000000,417.000000000000,
-717.000000000000,-692.000000000000,
243.000000000000,-465.000000000000,
846.000000000000,-144.000000000000,
562.000000000000,627.000000000000,
-415.000000000000,603.000000000000,
347.000000000000,-577.000000000000,
950.000000000000,889.000000000000,
-114.000000000000,388.000000000000,
-906.000000000000,-380.000000000000,
-249.000000000000,236.000000000000,
708.000000000000,-785.000000000000,
860.000000000000,172.000000000000,
-645.000000000000,1196.00000000000,
-731.000000000000,314.000000000000,
-354.000000000000,146.000000000000,
-601.000000000000,12.0000000000000,
-204.000000000000,444.000000000000,
-773.000000000000,64.0000000000000,
-337.000000000000,181.000000000000,
-2.00000000000000,472.000000000000,
125.000000000000,-1126.00000000000,
510.000000000000,265.000000000000,
903.000000000000,605.000000000000,
439.000000000000,-435.000000000000,
-297.000000000000,-323.000000000000,
-232.000000000000,-1216.00000000000,
103.000000000000,-609.000000000000,
-572.000000000000,-471.000000000000,
79.0000000000000,-854.000000000000,
1672.00000000000,216.000000000000,
319.000000000000,712.000000000000,
36.0000000000000,-366.000000000000,
-249.000000000000,-345.000000000000,
-615.000000000000,58.0000000000000,
102.000000000000,-549.000000000000,
-131.000000000000,1016.00000000000,
585.000000000000,261.000000000000,
492.000000000000,623.000000000000,
496.000000000000,733.000000000000,
-88.0000000000000,-380.000000000000,
184.000000000000,894.000000000000,
1049.00000000000,-185.000000000000,
-415.000000000000,117.000000000000,
489.000000000000,169.000000000000,
508.000000000000,-509.000000000000,
-404.000000000000,-282.000000000000,
323.000000000000,356.000000000000,
-622.000000000000,242.000000000000,
-912.000000000000,41.0000000000000,
-713.000000000000,700.000000000000,
-416.000000000000,-1316.00000000000,
806.000000000000,14.0000000000000,
329.000000000000,1209.00000000000,
-502.000000000000,-747.000000000000,
610.000000000000,-49.0000000000000,
386.000000000000,61.0000000000000,
-427.000000000000,-1175.00000000000,
77.0000000000000,-607.000000000000,
-151.000000000000,-814.000000000000,
589.000000000000,-945.000000000000,
464.000000000000,1205.00000000000,
-968.000000000000,277.000000000000,
166.000000000000,-703.000000000000,
446.000000000000,1027.00000000000,
486.000000000000,324.000000000000,
720.000000000000,-397.000000000000,
-224.000000000000,215.000000000000,
-395.000000000000,860.000000000000,
-808.000000000000,119.000000000000,
-444.000000000000,-1412.00000000000,
827.000000000000,-642.000000000000,
-119.000000000000,17.0000000000000,
-434.000000000000,725.000000000000,
343.000000000000,706.000000000000,
98.0000000000000,-707.000000000000,
951.000000000000,440.000000000000,
-286.000000000000,584.000000000000,
624.000000000000,-171.000000000000,
689.000000000000,140.000000000000,
-1028.00000000000,-268.000000000000,
579.000000000000,-525.000000000000,
-447.000000000000,-965.000000000000,
-729.000000000000,-119.000000000000,
-312.000000000000,-461.000000000000,
-508.000000000000,-1360.00000000000,
674.000000000000,-138.000000000000,
364.000000000000,379.000000000000,
-272.000000000000,-486.000000000000,
366.000000000000,-806.000000000000,
455.000000000000,-339.000000000000,
105.000000000000,12.0000000000000,
1158.00000000000,408.000000000000,
552.000000000000,273.000000000000,
54.0000000000000,217.000000000000,
988.000000000000,23.0000000000000,
537.000000000000,85.0000000000000,
267.000000000000,-9.00000000000000,
611.000000000000,-432.000000000000,
612.000000000000,688.000000000000,
-1003.00000000000,746.000000000000,
-1237.00000000000,192.000000000000,
-146.000000000000,-224.000000000000,
-451.000000000000,-958.000000000000,
461.000000000000,-282.000000000000,
208.000000000000,-621.000000000000,
2.00000000000000,-1021.00000000000,
493.000000000000,371.000000000000,
355.000000000000,794.000000000000,
860.000000000000,-193.000000000000,
-290.000000000000,339.000000000000,
-497.000000000000,-266.000000000000,
428.000000000000,-1209.00000000000,
609.000000000000,-313.000000000000,
598.000000000000,-395.000000000000,
-575.000000000000,345.000000000000,
-10.0000000000000,20.0000000000000,
271.000000000000,854.000000000000,
-735.000000000000,808.000000000000,
-714.000000000000,-90.0000000000000,
240.000000000000,104.000000000000,
344.000000000000,-772.000000000000,
-351.000000000000,429.000000000000,
3.00000000000000,-273.000000000000,
-1189.00000000000,-133.000000000000,
-419.000000000000,-139.000000000000,
836.000000000000,-861.000000000000,
-510.000000000000,653.000000000000,
-912.000000000000,-217.000000000000,
-501.000000000000,-536.000000000000,
-521.000000000000,152.000000000000,
-322.000000000000,7.00000000000000,
77.0000000000000,-1005.00000000000,
-147.000000000000,-1193.00000000000,
601.000000000000,22.0000000000000,
321.000000000000,483.000000000000,
-38.0000000000000,597.000000000000,
-457.000000000000,-239.000000000000,
-470.000000000000,-762.000000000000,
1033.00000000000,558.000000000000,
-666.000000000000,890.000000000000,
-771.000000000000,149.000000000000,
907.000000000000,-172.000000000000,
169.000000000000,558.000000000000,
432.000000000000,-25.0000000000000,
1079.00000000000,-388.000000000000,
-301.000000000000,288.000000000000,
-961.000000000000,-192.000000000000,
997.000000000000,-220.000000000000,
-74.0000000000000,969.000000000000,
-405.000000000000,1151.00000000000,
487.000000000000,-788.000000000000,
51.0000000000000,305.000000000000,
561.000000000000,711.000000000000,
-719.000000000000,-706.000000000000,
425.000000000000,98.0000000000000,
1181.00000000000,-54.0000000000000,
77.0000000000000,439.000000000000,
484.000000000000,249.000000000000,
352.000000000000,213.000000000000,
-19.0000000000000,-32.0000000000000,
-755.000000000000,8.00000000000000,
725.000000000000,78.0000000000000,
858.000000000000,-596.000000000000,
802.000000000000,1069.00000000000,
410.000000000000,24.0000000000000,
-617.000000000000,-19.0000000000000,
603.000000000000,374.000000000000,
-1374.00000000000,205.000000000000,
-398.000000000000,-15.0000000000000,
1068.00000000000,-514.000000000000,
-317.000000000000,1063.00000000000,
-807.000000000000,-926.000000000000,
257.000000000000,-755.000000000000,
1544.00000000000,355.000000000000,
872.000000000000,19.0000000000000,
1017.00000000000,1104.00000000000,
-981.000000000000,-150.000000000000,
-84.0000000000000,-355.000000000000,
1318.00000000000,-172.000000000000,
703.000000000000,396.000000000000,
837.000000000000,332.000000000000,
54.0000000000000,-617.000000000000,
372.000000000000,443.000000000000,
-395.000000000000,206.000000000000,
695.000000000000,-123.000000000000,
596.000000000000,789.000000000000,
-896.000000000000,640.000000000000,
345.000000000000,378.000000000000,
-377.000000000000,1137.00000000000,
-224.000000000000,681.000000000000,
935.000000000000,-301.000000000000,
-17.0000000000000,-253.000000000000,
-848.000000000000,129.000000000000,
-377.000000000000,778.000000000000,
-451.000000000000,-885.000000000000,
-23.0000000000000,14.0000000000000,
-74.0000000000000,1408.00000000000,
-1258.00000000000,-827.000000000000,
837.000000000000,182.000000000000,
345.000000000000,230.000000000000,
143.000000000000,40.0000000000000,
674.000000000000,626.000000000000,
-689.000000000000,-950.000000000000,
667.000000000000,-699.000000000000,
-521.000000000000,554.000000000000,
543.000000000000,679.000000000000,
-2.00000000000000,-290.000000000000,
-1392.00000000000,87.0000000000000,
373.000000000000,-794.000000000000,
-232.000000000000,-117.000000000000,
558.000000000000,395.000000000000,
-145.000000000000,-1024.00000000000,
173.000000000000,138.000000000000,
436.000000000000,204.000000000000,
9.00000000000000,1142.00000000000,
138.000000000000,807.000000000000,
-872.000000000000,616.000000000000,
120.000000000000,105.000000000000,
-473.000000000000,-1125.00000000000,
-686.000000000000,126.000000000000,
-142.000000000000,162.000000000000,
773.000000000000,-144.000000000000,
1164.00000000000,-268.000000000000,
17.0000000000000,599.000000000000,
-449.000000000000,457.000000000000,
-993.000000000000,-190.000000000000,
-138.000000000000,-52.0000000000000,
-861.000000000000,-933.000000000000,
265.000000000000,-73.0000000000000,
908.000000000000,-540.000000000000,
-901.000000000000,131.000000000000,
288.000000000000,1071.00000000000,
-299.000000000000,227.000000000000,
-155.000000000000,-64.0000000000000,
403.000000000000,-1458.00000000000,
103.000000000000,-400.000000000000,
-262.000000000000,426.000000000000,
-695.000000000000,-598.000000000000,
144.000000000000,-511.000000000000,
-176.000000000000,-129.000000000000,
200.000000000000,-950.000000000000,
260.000000000000,-536.000000000000,
-488.000000000000,1037.00000000000,
-170.000000000000,96.0000000000000,
-330.000000000000,-669.000000000000,
395.000000000000,-771.000000000000,
616.000000000000,-346.000000000000,
-625.000000000000,-108.000000000000,
51.0000000000000,-56.0000000000000,
336.000000000000,0.00000000000000,
-189.000000000000,-101.000000000000,
836.000000000000,602.000000000000,
149.000000000000,-370.000000000000,
-962.000000000000,-121.000000000000,
907.000000000000,456.000000000000,
557.000000000000,305.000000000000,
-417.000000000000,466.000000000000,
275.000000000000,-646.000000000000,
941.000000000000,-57.0000000000000,
1306.00000000000,-21.0000000000000,
-420.000000000000,839.000000000000,
473.000000000000,940.000000000000,
458.000000000000,-363.000000000000,
-404.000000000000,699.000000000000,
221.000000000000,-878.000000000000,
388.000000000000,-492.000000000000,
766.000000000000,-10.0000000000000,
-147.000000000000,-110.000000000000,
-222.000000000000,938.000000000000,
-873.000000000000,11.0000000000000,
469.000000000000,716.000000000000,
-115.000000000000,15.0000000000000,
-206.000000000000,-846.000000000000,
701.000000000000,-125.000000000000,
-500.000000000000,704.000000000000,
521.000000000000,245.000000000000,
-883.000000000000,-448.000000000000,
-571.000000000000,172.000000000000,
-331.000000000000,-1031.00000000000,
-215.000000000000,67.0000000000000,
1167.00000000000,724.000000000000,
50.0000000000000,-800.000000000000,
77.0000000000000,128.000000000000,
272.000000000000,353.000000000000,
-534.000000000000,-106.000000000000,
-1236.00000000000,-663.000000000000,
511.000000000000,-839.000000000000,
309.000000000000,86.0000000000000,
-1115.00000000000,282.000000000000,
579.000000000000,-153.000000000000,
510.000000000000,-197.000000000000,
-162.000000000000,-520.000000000000,
525.000000000000,-83.0000000000000,
-348.000000000000,629.000000000000,
-232.000000000000,466.000000000000,
-217.000000000000,1008.00000000000,
-963.000000000000,112.000000000000,
-596.000000000000,-68.0000000000000,
-695.000000000000,412.000000000000,
-376.000000000000,-429.000000000000,
100.000000000000,-808.000000000000,
654.000000000000,-787.000000000000,
1164.00000000000,368.000000000000,
-346.000000000000,136.000000000000,
-1024.00000000000,-252.000000000000,
-124.000000000000,708.000000000000,
-978.000000000000,10.0000000000000,
-93.0000000000000,-645.000000000000,
545.000000000000,-508.000000000000,
-1295.00000000000,58.0000000000000,
-265.000000000000,-311.000000000000,
-109.000000000000,-81.0000000000000,
-698.000000000000,579.000000000000,
-429.000000000000,-468.000000000000,
50.0000000000000,-379.000000000000,
105.000000000000,798.000000000000,
-716.000000000000,1175.00000000000,
201.000000000000,-717.000000000000,
285.000000000000,-557.000000000000,
-593.000000000000,769.000000000000,
-995.000000000000,-868.000000000000,
358.000000000000,153.000000000000,
52.0000000000000,938.000000000000,
-1420.00000000000,249.000000000000,
-546.000000000000,-644.000000000000,
164.000000000000,-877.000000000000,
765.000000000000,318.000000000000,
17.0000000000000,7.00000000000000,
793.000000000000,776.000000000000,
-262.000000000000,324.000000000000,
148.000000000000,-552.000000000000,
903.000000000000,482.000000000000,
-1193.00000000000,-768.000000000000,
-15.0000000000000,-862.000000000000,
-417.000000000000,-718.000000000000,
613.000000000000,-932.000000000000,
1138.00000000000,-343.000000000000,
-142.000000000000,1113.00000000000,
204.000000000000,1300.00000000000,
-788.000000000000,-607.000000000000,
-29.0000000000000,-571.000000000000,
250.000000000000,494.000000000000,
88.0000000000000,-170.000000000000,
913.000000000000,-575.000000000000,
-241.000000000000,496.000000000000,
-740.000000000000,-484.000000000000,
332.000000000000,-286.000000000000,
190.000000000000,403.000000000000,
-126.000000000000,-48.0000000000000,
820.000000000000,-162.000000000000,
629.000000000000,-83.0000000000000,
-840.000000000000,507.000000000000,
0.00000000000000,-509.000000000000,
1438.00000000000,-432.000000000000,
276.000000000000,874.000000000000,
135.000000000000,407.000000000000,
660.000000000000,194.000000000000,
-151.000000000000,709.000000000000,
-470.000000000000,-414.000000000000,
159.000000000000,-1075.00000000000,
1204.00000000000,68.0000000000000,
1104.00000000000,72.0000000000000,
-824.000000000000,120.000000000000,
391.000000000000,-106.000000000000,
1066.00000000000,7.00000000000000,
-441.000000000000,1614.00000000000,
330.000000000000,-105.000000000000,
-789.000000000000,53.0000000000000,
-460.000000000000,-397.000000000000,
505.000000000000,-45.0000000000000,
-126.000000000000,1357.00000000000,
-591.000000000000,-839.000000000000,
-773.000000000000,-10.0000000000000,
109.000000000000,-631.000000000000,
-786.000000000000,-701.000000000000,
511.000000000000,-276.000000000000,
467.000000000000,564.000000000000,
-880.000000000000,413.000000000000,
401.000000000000,-224.000000000000,
-831.000000000000,759.000000000000,
-921.000000000000,-331.000000000000,
376.000000000000,-350.000000000000,
763.000000000000,-607.000000000000,
1185.00000000000,-47.0000000000000,
593.000000000000,-3.00000000000000,
623.000000000000,-646.000000000000,
-91.0000000000000,95.0000000000000,
-212.000000000000,114.000000000000,
73.0000000000000,111.000000000000,
-746.000000000000,-117.000000000000,
-681.000000000000,342.000000000000,
-553.000000000000,244.000000000000,
-1227.00000000000,-537.000000000000,
-76.0000000000000,560.000000000000,
266.000000000000,932.000000000000,
-123.000000000000,-340.000000000000,
691.000000000000,-1426.00000000000,
-177.000000000000,33.0000000000000,
539.000000000000,570.000000000000,
289.000000000000,-1204.00000000000,
-686.000000000000,-228.000000000000,
-139.000000000000,436.000000000000,
-103.000000000000,732.000000000000,
349.000000000000,976.000000000000,
-302.000000000000,272.000000000000,
-163.000000000000,-529.000000000000,
827.000000000000,-432.000000000000,
518.000000000000,938.000000000000,
8.00000000000000,1143.00000000000,
-369.000000000000,533.000000000000,
-395.000000000000,750.000000000000,
-399.000000000000,1171.00000000000,
-400.000000000000,1031.00000000000,
-103.000000000000,570.000000000000,
-445.000000000000,50.0000000000000,
-710.000000000000,303.000000000000,
-137.000000000000,1023.00000000000,
-82.0000000000000,650.000000000000,
523.000000000000,22.0000000000000,
561.000000000000,563.000000000000,
-630.000000000000,1247.00000000000,
-272.000000000000,863.000000000000,
-332.000000000000,139.000000000000,
-1124.00000000000,-188.000000000000,
-376.000000000000,-489.000000000000,
201.000000000000,-198.000000000000,
-378.000000000000,-188.000000000000,
-829.000000000000,-618.000000000000,
410.000000000000,268.000000000000,
-1097.00000000000,77.0000000000000,
-872.000000000000,501.000000000000,
1437.00000000000,-87.0000000000000,
491.000000000000,-267.000000000000,
-150.000000000000,365.000000000000,
-1090.00000000000,-255.000000000000,
242.000000000000,626.000000000000,
-224.000000000000,-843.000000000000,
-202.000000000000,-480.000000000000,
1086.00000000000,327.000000000000,
-1473.00000000000,-13.0000000000000,
-429.000000000000,616.000000000000,
-272.000000000000,383.000000000000,
-978.000000000000,-522.000000000000,
330.000000000000,-95.0000000000000,
-4.00000000000000,1006.00000000000,
73.0000000000000,-501.000000000000,
-391.000000000000,-85.0000000000000,
127.000000000000,-738.000000000000,
963.000000000000,-687.000000000000,
-212.000000000000,-159.000000000000,
462.000000000000,-1096.00000000000,
662.000000000000,159.000000000000,
428.000000000000,1163.00000000000,
296.000000000000,317.000000000000,
-473.000000000000,-770.000000000000,
-441.000000000000,61.0000000000000,
-1265.00000000000,89.0000000000000,
-248.000000000000,-86.0000000000000,
1372.00000000000,103.000000000000,
1165.00000000000,368.000000000000,
-71.0000000000000,1084.00000000000,
-1353.00000000000,305.000000000000,
-221.000000000000,-567.000000000000,
948.000000000000,244.000000000000,
-904.000000000000,283.000000000000,
68.0000000000000,-127.000000000000,
434.000000000000,-512.000000000000,
-935.000000000000,450.000000000000,
727.000000000000,-499.000000000000,
-320.000000000000,-934.000000000000,
223.000000000000,-362.000000000000,
-202.000000000000,-912.000000000000,
-763.000000000000,761.000000000000,
544.000000000000,103.000000000000,
-294.000000000000,1258.00000000000,
469.000000000000,762.000000000000,
-296.000000000000,-1620.00000000000,
126.000000000000,-837.000000000000,
734.000000000000,162.000000000000,
-7.00000000000000,719.000000000000,
333.000000000000,-604.000000000000,
1067.00000000000,442.000000000000,
570.000000000000,34.0000000000000,
-1078.00000000000,-417.000000000000,
716.000000000000,921.000000000000,
679.000000000000,13.0000000000000,
138.000000000000,213.000000000000,
330.000000000000,267.000000000000,
-365.000000000000,148.000000000000,
44.0000000000000,-104.000000000000,
-554.000000000000,277.000000000000,
390.000000000000,-432.000000000000,
431.000000000000,-863.000000000000,
1169.00000000000,136.000000000000,
1557.00000000000,367.000000000000,
-914.000000000000,1112.00000000000,
259.000000000000,-537.000000000000,
176.000000000000,537.000000000000,
-993.000000000000,669.000000000000,
-195.000000000000,-1253.00000000000,
635.000000000000,71.0000000000000,
297.000000000000,730.000000000000,
-92.0000000000000,1655.00000000000,
283.000000000000,-384.000000000000,
-664.000000000000,-563.000000000000,
-415.000000000000,436.000000000000,
-839.000000000000,-190.000000000000,
93.0000000000000,-41.0000000000000,
-515.000000000000,-724.000000000000,
-484.000000000000,947.000000000000,
912.000000000000,-313.000000000000,
-299.000000000000,-778.000000000000,
1243.00000000000,991.000000000000,
104.000000000000,517.000000000000,
-1039.00000000000,272.000000000000,
-316.000000000000,-1135.00000000000,
264.000000000000,315.000000000000,
527.000000000000,599.000000000000,
78.0000000000000,-502.000000000000,
1142.00000000000,194.000000000000,
532.000000000000,471.000000000000,
282.000000000000,1537.00000000000,
-807.000000000000,546.000000000000,
202.000000000000,251.000000000000,
-5.00000000000000,240.000000000000,
-773.000000000000,63.0000000000000,
1295.00000000000,-68.0000000000000,
-79.0000000000000,-690.000000000000,
835.000000000000,58.0000000000000,
261.000000000000,515.000000000000,
-1133.00000000000,422.000000000000,
-492.000000000000,-1151.00000000000,
-943.000000000000,79.0000000000000,
14.0000000000000,1124.00000000000,
-416.000000000000,1006.00000000000,
409.000000000000,903.000000000000,
-338.000000000000,-423.000000000000,
-1749.00000000000,-172.000000000000,
982.000000000000,-965.000000000000,
561.000000000000,170.000000000000,
-465.000000000000,376.000000000000,
465.000000000000,-849.000000000000,
-484.000000000000,-192.000000000000,
-664.000000000000,65.0000000000000,
910.000000000000,-324.000000000000,
543.000000000000,-930.000000000000,
429.000000000000,-402.000000000000,
385.000000000000,91.0000000000000,
35.0000000000000,-173.000000000000,
981.000000000000,-78.0000000000000,
389.000000000000,157.000000000000,
-284.000000000000,1027.00000000000,
-366.000000000000,490.000000000000,
806.000000000000,-150.000000000000,
251.000000000000,1135.00000000000,
-1037.00000000000,294.000000000000,
636.000000000000,-690.000000000000,
-188.000000000000,-41.0000000000000,
-616.000000000000,750.000000000000,
-52.0000000000000,-234.000000000000,
-267.000000000000,-782.000000000000,
-485.000000000000,-178.000000000000,
-335.000000000000,-342.000000000000,
791.000000000000,-139.000000000000,
339.000000000000,-703.000000000000,
1153.00000000000,222.000000000000,
531.000000000000,306.000000000000,
272.000000000000,-316.000000000000,
1203.00000000000,886.000000000000,
-855.000000000000,1474.00000000000,
-545.000000000000,3.00000000000000,
-29.0000000000000,-1191.00000000000,
159.000000000000,-727.000000000000,
1016.00000000000,-708.000000000000,
253.000000000000,413.000000000000,
-406.000000000000,458.000000000000,
-811.000000000000,841.000000000000,
223.000000000000,-174.000000000000,
211.000000000000,-1161.00000000000,
750.000000000000,-231.000000000000,
809.000000000000,-50.0000000000000,
-783.000000000000,948.000000000000,
160.000000000000,386.000000000000,
-689.000000000000,549.000000000000,
-631.000000000000,-616.000000000000,
498.000000000000,147.000000000000,
137.000000000000,1470.00000000000,
163.000000000000,-1386.00000000000,
705.000000000000,538.000000000000,
-171.000000000000,724.000000000000,
-1200.00000000000,-903.000000000000,
419.000000000000,77.0000000000000,
243.000000000000,180.000000000000,
-48.0000000000000,1484.00000000000,
-322.000000000000,3.00000000000000,
400.000000000000,-595.000000000000,
-7.00000000000000,738.000000000000,
-1012.00000000000,-1136.00000000000,
356.000000000000,-1046.00000000000,
434.000000000000,72.0000000000000,
739.000000000000,-68.0000000000000,
159.000000000000,396.000000000000,
-125.000000000000,-202.000000000000,
602.000000000000,281.000000000000,
-173.000000000000,1014.00000000000,
-438.000000000000,-195.000000000000,
571.000000000000,332.000000000000,
1038.00000000000,107.000000000000,
649.000000000000,642.000000000000,
-832.000000000000,1139.00000000000,
-531.000000000000,-592.000000000000,
-871.000000000000,299.000000000000,
-462.000000000000,-519.000000000000,
831.000000000000,-3.00000000000000,
122.000000000000,324.000000000000,
-495.000000000000,-1073.00000000000,
-560.000000000000,920.000000000000,
292.000000000000,629.000000000000,
260.000000000000,-19.0000000000000,
-381.000000000000,47.0000000000000,
-570.000000000000,92.0000000000000,
735.000000000000,599.000000000000,
501.000000000000,-344.000000000000,
198.000000000000,372.000000000000,
-326.000000000000,586.000000000000,
-1444.00000000000,-769.000000000000,
257.000000000000,-936.000000000000,
553.000000000000,-268.000000000000,
225.000000000000,-259.000000000000,
454.000000000000,515.000000000000,
408.000000000000,1223.00000000000,
110.000000000000,-16.0000000000000,
208.000000000000,97.0000000000000,
1021.00000000000,83.0000000000000,
941.000000000000,-315.000000000000,
-317.000000000000,53.0000000000000,
-577.000000000000,-1035.00000000000,
261.000000000000,-739.000000000000,
-1010.00000000000,209.000000000000,
-760.000000000000,-292.000000000000,
506.000000000000,557.000000000000,
340.000000000000,492.000000000000,
796.000000000000,-44.0000000000000,
1008.00000000000,93.0000000000000,
-336.000000000000,-126.000000000000,
-58.0000000000000,-21.0000000000000,
583.000000000000,-697.000000000000,
-211.000000000000,114.000000000000,
460.000000000000,490.000000000000,
286.000000000000,716.000000000000,
-344.000000000000,626.000000000000,
-125.000000000000,-1059.00000000000,
-13.0000000000000,-85.0000000000000,
-237.000000000000,373.000000000000,
-333.000000000000,-1497.00000000000,
665.000000000000,-1039.00000000000,
595.000000000000,592.000000000000,
-490.000000000000,1052.00000000000,
310.000000000000,282.000000000000,
1201.00000000000,-219.000000000000,
867.000000000000,99.0000000000000,
828.000000000000,-514.000000000000,
114.000000000000,-231.000000000000,
397.000000000000,-453.000000000000,
541.000000000000,-785.000000000000,
283.000000000000,391.000000000000,
-335.000000000000,336.000000000000,
-927.000000000000,592.000000000000,
-393.000000000000,0.00000000000000,
-543.000000000000,181.000000000000,
-103.000000000000,430.000000000000,
-309.000000000000,-312.000000000000,
-2.00000000000000,57.0000000000000,
148.000000000000,-697.000000000000,
-485.000000000000,-396.000000000000,
-169.000000000000,-317.000000000000,
-440.000000000000,-872.000000000000,
299.000000000000,-769.000000000000,
195.000000000000,264.000000000000,
-170.000000000000,276.000000000000,
562.000000000000,208.000000000000,
348.000000000000,1037.00000000000,
964.000000000000,-38.0000000000000,
804.000000000000,-533.000000000000,
-837.000000000000,237.000000000000,
9.00000000000000,-61.0000000000000,
70.0000000000000,-885.000000000000,
-1382.00000000000,-420.000000000000,
-284.000000000000,595.000000000000,
186.000000000000,103.000000000000,
98.0000000000000,-608.000000000000,
775.000000000000,-558.000000000000,
221.000000000000,-823.000000000000,
519.000000000000,-266.000000000000,
1004.00000000000,153.000000000000,
270.000000000000,18.0000000000000,
-161.000000000000,424.000000000000,
138.000000000000,-356.000000000000,
739.000000000000,-1010.00000000000,
475.000000000000,317.000000000000,
520.000000000000,505.000000000000,
753.000000000000,-358.000000000000,
802.000000000000,977.000000000000,
36.0000000000000,825.000000000000,
7.00000000000000,407.000000000000,
532.000000000000,239.000000000000,
364.000000000000,73.0000000000000,
648.000000000000,313.000000000000,
-1058.00000000000,191.000000000000,
-299.000000000000,691.000000000000,
52.0000000000000,-647.000000000000,
-1537.00000000000,-162.000000000000,
-772.000000000000,11.0000000000000,
304.000000000000,-951.000000000000,
1332.00000000000,696.000000000000,
-470.000000000000,143.000000000000,
38.0000000000000,356.000000000000,
800.000000000000,383.000000000000,
-291.000000000000,41.0000000000000,
-290.000000000000,96.0000000000000,
-960.000000000000,136.000000000000,
-708.000000000000,426.000000000000,
-721.000000000000,-1077.00000000000,
-8.00000000000000,-801.000000000000,
-23.0000000000000,-518.000000000000,
750.000000000000,-396.000000000000,
211.000000000000,592.000000000000,
-981.000000000000,-218.000000000000,
353.000000000000,-751.000000000000,
-73.0000000000000,-437.000000000000,
694.000000000000,80.0000000000000,
340.000000000000,-1113.00000000000,
704.000000000000,-107.000000000000,
267.000000000000,824.000000000000,
-1580.00000000000,-212.000000000000,
-236.000000000000,-402.000000000000,
-17.0000000000000,-1665.00000000000,
823.000000000000,89.0000000000000,
184.000000000000,538.000000000000,
464.000000000000,-171.000000000000,
487.000000000000,-270.000000000000,
-849.000000000000,-422.000000000000,
442.000000000000,187.000000000000,
-524.000000000000,-565.000000000000,
-270.000000000000,122.000000000000,
-626.000000000000,131.000000000000,
-766.000000000000,58.0000000000000,
187.000000000000,561.000000000000,
51.0000000000000,608.000000000000,
190.000000000000,-293.000000000000,
-432.000000000000,-457.000000000000,
248.000000000000,-83.0000000000000,
-98.0000000000000,-1633.00000000000,
547.000000000000,101.000000000000,
639.000000000000,-42.0000000000000,
325.000000000000,-809.000000000000,
929.000000000000,1357.00000000000,
-414.000000000000,146.000000000000,
-27.0000000000000,-134.000000000000,
160.000000000000,107.000000000000,
896.000000000000,-23.0000000000000,
-411.000000000000,498.000000000000,
-1067.00000000000,-107.000000000000,
929.000000000000,-387.000000000000,
133.000000000000,160.000000000000,
652.000000000000,599.000000000000,
693.000000000000,-982.000000000000,
807.000000000000,376.000000000000,
-56.0000000000000,887.000000000000,
-765.000000000000,-45.0000000000000,
27.0000000000000,530.000000000000,
177.000000000000,-159.000000000000,
518.000000000000,446.000000000000,
-288.000000000000,28.0000000000000,
580.000000000000,-413.000000000000,
-78.0000000000000,582.000000000000,
-675.000000000000,179.000000000000,
458.000000000000,-25.0000000000000,
-342.000000000000,737.000000000000,
639.000000000000,611.000000000000,
806.000000000000,541.000000000000,
-652.000000000000,413.000000000000,
637.000000000000,-351.000000000000,
919.000000000000,-46.0000000000000,
84.0000000000000,4.00000000000000,
-7.00000000000000,1029.00000000000,
-417.000000000000,1179.00000000000,
230.000000000000,241.000000000000,
338.000000000000,897.000000000000,
-952.000000000000,-35.0000000000000,
-532.000000000000,-452.000000000000,
-211.000000000000,108.000000000000,
36.0000000000000,-1081.00000000000,
305.000000000000,303.000000000000,
169.000000000000,746.000000000000,
525.000000000000,359.000000000000,
-372.000000000000,837.000000000000,
-178.000000000000,-1121.00000000000,
267.000000000000,432.000000000000,
-341.000000000000,849.000000000000,
33.0000000000000,-1358.00000000000,
673.000000000000,-130.000000000000,
-519.000000000000,129.000000000000,
-888.000000000000,-263.000000000000,
320.000000000000,-73.0000000000000,
164.000000000000,-1082.00000000000,
-131.000000000000,-685.000000000000,
-422.000000000000,195.000000000000,
-703.000000000000,-179.000000000000,
845.000000000000,-478.000000000000,
62.0000000000000,-237.000000000000,
-804.000000000000,611.000000000000,
296.000000000000,-688.000000000000,
-283.000000000000,158.000000000000,
842.000000000000,815.000000000000,
284.000000000000,-1380.00000000000,
-168.000000000000,-737.000000000000,
1130.00000000000,-286.000000000000,
138.000000000000,-337.000000000000,
-226.000000000000,21.0000000000000,
137.000000000000,805.000000000000,
823.000000000000,514.000000000000,
816.000000000000,-368.000000000000,
-143.000000000000,269.000000000000,
-79.0000000000000,244.000000000000,
1034.00000000000,724.000000000000,
-112.000000000000,698.000000000000,
-460.000000000000,-503.000000000000,
213.000000000000,165.000000000000,
-219.000000000000,65.0000000000000,
-192.000000000000,-338.000000000000,
-949.000000000000,-136.000000000000,
-498.000000000000,-451.000000000000,
-613.000000000000,-1072.00000000000,
328.000000000000,-925.000000000000,
919.000000000000,959.000000000000,
-70.0000000000000,35.0000000000000,
-78.0000000000000,41.0000000000000,
-545.000000000000,-212.000000000000,
-86.0000000000000,-1324.00000000000,
525.000000000000,166.000000000000,
1198.00000000000,131.000000000000,
108.000000000000,712.000000000000,
-336.000000000000,101.000000000000,
570.000000000000,-106.000000000000,
-1065.00000000000,352.000000000000,
-435.000000000000,-186.000000000000,
-585.000000000000,-634.000000000000,
-1173.00000000000,33.0000000000000,
-57.0000000000000,-243.000000000000,
-234.000000000000,-1405.00000000000,
705.000000000000,-601.000000000000,
-120.000000000000,-783.000000000000,
-302.000000000000,-58.0000000000000,
150.000000000000,-763.000000000000,
-4.00000000000000,-987.000000000000,
730.000000000000,540.000000000000,
103.000000000000,439.000000000000,
40.0000000000000,246.000000000000,
-212.000000000000,-287.000000000000,
616.000000000000,421.000000000000,
643.000000000000,-391.000000000000,
842.000000000000,422.000000000000,
161.000000000000,823.000000000000,
-1288.00000000000,-513.000000000000,
772.000000000000,622.000000000000,
-1186.00000000000,-116.000000000000,
-1090.00000000000,-377.000000000000,
389.000000000000,369.000000000000,
-690.000000000000,1089.00000000000,
402.000000000000,-67.0000000000000,
-107.000000000000,457.000000000000,
93.0000000000000,973.000000000000,
-501.000000000000,17.0000000000000,
-155.000000000000,714.000000000000,
560.000000000000,-72.0000000000000,
-724.000000000000,782.000000000000,
618.000000000000,117.000000000000,
383.000000000000,418.000000000000,
-127.000000000000,1119.00000000000,
-87.0000000000000,424.000000000000,
596.000000000000,720.000000000000,
719.000000000000,-398.000000000000,
-259.000000000000,-165.000000000000,
114.000000000000,-753.000000000000,
354.000000000000,249.000000000000,
913.000000000000,536.000000000000,
-433.000000000000,-901.000000000000,
82.0000000000000,-694.000000000000,
352.000000000000,-376.000000000000,
-99.0000000000000,1054.00000000000,
1281.00000000000,155.000000000000,
-333.000000000000,1059.00000000000,
-87.0000000000000,1570.00000000000,
-159.000000000000,320.000000000000,
-973.000000000000,706.000000000000,
6.00000000000000,39.0000000000000,
-168.000000000000,-315.000000000000,
-124.000000000000,-45.0000000000000,
-877.000000000000,-44.0000000000000,
-420.000000000000,-929.000000000000,
-119.000000000000,536.000000000000,
-1195.00000000000,62.0000000000000,
243.000000000000,-458.000000000000,
957.000000000000,608.000000000000,
-130.000000000000,-498.000000000000,
-646.000000000000,164.000000000000,
-168.000000000000,-790.000000000000,
-134.000000000000,-577.000000000000,
-162.000000000000,1078.00000000000,
-820.000000000000,38.0000000000000,
-166.000000000000,623.000000000000,
764.000000000000,-137.000000000000,
221.000000000000,-396.000000000000,
123.000000000000,370.000000000000,
-1337.00000000000,-616.000000000000,
-539.000000000000,-144.000000000000,
-547.000000000000,-78.0000000000000,
-389.000000000000,-105.000000000000,
63.0000000000000,-347.000000000000,
-1114.00000000000,260.000000000000,
-450.000000000000,-315.000000000000,
-1086.00000000000,-217.000000000000,
253.000000000000,569.000000000000,
753.000000000000,116.000000000000,
-178.000000000000,1230.00000000000,
643.000000000000,718.000000000000,
-337.000000000000,387.000000000000,
-115.000000000000,-188.000000000000,
917.000000000000,-592.000000000000,
-175.000000000000,285.000000000000,
-261.000000000000,-414.000000000000,
334.000000000000,-686.000000000000,
-762.000000000000,446.000000000000,
68.0000000000000,14.0000000000000,
1239.00000000000,-808.000000000000,
-478.000000000000,683.000000000000,
-466.000000000000,-252.000000000000,
-375.000000000000,-461.000000000000,
-520.000000000000,853.000000000000,
236.000000000000,-790.000000000000,
-501.000000000000,-341.000000000000,
730.000000000000,-350.000000000000,
843.000000000000,-657.000000000000,
539.000000000000,-479.000000000000,
1040.00000000000,-509.000000000000,
843.000000000000,831.000000000000,
-472.000000000000,300.000000000000,
-685.000000000000,1151.00000000000,
-725.000000000000,362.000000000000,
-1227.00000000000,424.000000000000,
327.000000000000,981.000000000000,
-943.000000000000,-940.000000000000,
-58.0000000000000,389.000000000000,
-81.0000000000000,-292.000000000000,
-605.000000000000,-521.000000000000,
349.000000000000,136.000000000000,
-1712.00000000000,-559.000000000000,
-615.000000000000,-450.000000000000,
-471.000000000000,-524.000000000000,
-340.000000000000,-218.000000000000,
1014.00000000000,-326.000000000000,
1141.00000000000,314.000000000000,
1008.00000000000,18.0000000000000,
840.000000000000,450.000000000000,
922.000000000000,472.000000000000,
45.0000000000000,-685.000000000000,
-196.000000000000,-229.000000000000,
-1287.00000000000,-373.000000000000,
-614.000000000000,806.000000000000,
-143.000000000000,-105.000000000000,
-892.000000000000,-590.000000000000,
605.000000000000,553.000000000000,
-356.000000000000,-621.000000000000,
-477.000000000000,-525.000000000000,
-530.000000000000,-301.000000000000,
-339.000000000000,139.000000000000,
607.000000000000,553.000000000000,
-661.000000000000,39.0000000000000,
-469.000000000000,-396.000000000000,
631.000000000000,-643.000000000000,
661.000000000000,-406.000000000000,
245.000000000000,-310.000000000000,
-72.0000000000000,-302.000000000000,
121.000000000000,-491.000000000000,
389.000000000000,92.0000000000000,
-1066.00000000000,144.000000000000,
-296.000000000000,-75.0000000000000,
1285.00000000000,486.000000000000,
-1301.00000000000,325.000000000000,
-627.000000000000,-181.000000000000,
1190.00000000000,-593.000000000000,
-16.0000000000000,899.000000000000,
-375.000000000000,1059.00000000000,
-697.000000000000,-1312.00000000000,
792.000000000000,-714.000000000000,
625.000000000000,723.000000000000,
-368.000000000000,65.0000000000000,
1093.00000000000,-277.000000000000,
-334.000000000000,960.000000000000,
-1116.00000000000,588.000000000000,
-194.000000000000,286.000000000000,
-938.000000000000,301.000000000000,
-87.0000000000000,-553.000000000000,
625.000000000000,-246.000000000000,
-263.000000000000,-88.0000000000000,
28.0000000000000,-719.000000000000,
393.000000000000,-761.000000000000,
566.000000000000,-263.000000000000,
357.000000000000,-326.000000000000,
-723.000000000000,122.000000000000,
106.000000000000,799.000000000000,
191.000000000000,224.000000000000,
-238.000000000000,717.000000000000,
-527.000000000000,1198.00000000000,
170.000000000000,-216.000000000000,
999.000000000000,655.000000000000,
159.000000000000,34.0000000000000,
364.000000000000,344.000000000000,
-361.000000000000,977.000000000000,
232.000000000000,-115.000000000000,
422.000000000000,608.000000000000,
208.000000000000,458.000000000000,
319.000000000000,438.000000000000,
-1024.00000000000,-796.000000000000,
628.000000000000,211.000000000000,
-671.000000000000,610.000000000000,
-686.000000000000,-482.000000000000,
346.000000000000,728.000000000000,
-816.000000000000,764.000000000000,
-225.000000000000,700.000000000000,
-680.000000000000,-103.000000000000,
395.000000000000,-468.000000000000,
43.0000000000000,-251.000000000000,
-333.000000000000,637.000000000000,
828.000000000000,-337.000000000000,
78.0000000000000,-1059.00000000000,
79.0000000000000,-60.0000000000000,
254.000000000000,-910.000000000000,
140.000000000000,220.000000000000,
-334.000000000000,363.000000000000,
-267.000000000000,-1337.00000000000,
329.000000000000,-281.000000000000,
-200.000000000000,633.000000000000,
-613.000000000000,554.000000000000,
383.000000000000,351.000000000000,
-59.0000000000000,417.000000000000,
-455.000000000000,724.000000000000,
797.000000000000,590.000000000000,
-443.000000000000,398.000000000000,
-885.000000000000,351.000000000000,
-557.000000000000,-433.000000000000,
-635.000000000000,-1043.00000000000,
1223.00000000000,-990.000000000000,
-92.0000000000000,-786.000000000000,
-782.000000000000,486.000000000000,
613.000000000000,144.000000000000,
-657.000000000000,836.000000000000,
2.00000000000000,936.000000000000,
-1101.00000000000,-436.000000000000,
-814.000000000000,-616.000000000000,
637.000000000000,-761.000000000000,
-477.000000000000,315.000000000000,
-499.000000000000,-1146.00000000000,
33.0000000000000,339.000000000000,
335.000000000000,690.000000000000,
-977.000000000000,-783.000000000000,
47.0000000000000,747.000000000000,
-65.0000000000000,-378.000000000000,
-348.000000000000,146.000000000000,
-379.000000000000,-128.000000000000,
-895.000000000000,-303.000000000000,
1101.00000000000,609.000000000000,
-422.000000000000,1008.00000000000,
-72.0000000000000,481.000000000000,
209.000000000000,102.000000000000,
-82.0000000000000,1289.00000000000,
136.000000000000,175.000000000000,
-1525.00000000000,23.0000000000000,
-638.000000000000,-744.000000000000,
-217.000000000000,-186.000000000000,
515.000000000000,178.000000000000,
135.000000000000,-563.000000000000,
-685.000000000000,608.000000000000,
-67.0000000000000,-973.000000000000,
-837.000000000000,-111.000000000000,
-645.000000000000,-282.000000000000,
371.000000000000,-1458.00000000000,
495.000000000000,501.000000000000,
-434.000000000000,-176.000000000000,
776.000000000000,-38.0000000000000,
574.000000000000,683.000000000000,
535.000000000000,94.0000000000000,
373.000000000000,-91.0000000000000,
-956.000000000000,-587.000000000000,
1139.00000000000,-798.000000000000,
208.000000000000,913.000000000000,
-226.000000000000,950.000000000000,
691.000000000000,-450.000000000000,
-420.000000000000,1042.00000000000,
632.000000000000,-216.000000000000,
389.000000000000,-843.000000000000,
-487.000000000000,23.0000000000000,
-1027.00000000000,-490.000000000000,
-404.000000000000,-918.000000000000,
227.000000000000,-1313.00000000000,
-704.000000000000,593.000000000000,
684.000000000000,-212.000000000000,
498.000000000000,-367.000000000000,
-219.000000000000,304.000000000000,
-133.000000000000,-764.000000000000,
214.000000000000,-144.000000000000,
16.0000000000000,399.000000000000,
301.000000000000,635.000000000000,
715.000000000000,-360.000000000000,
-168.000000000000,478.000000000000,
876.000000000000,181.000000000000,
437.000000000000,-422.000000000000,
315.000000000000,837.000000000000,
157.000000000000,-943.000000000000,
-335.000000000000,-517.000000000000,
60.0000000000000,106.000000000000,
674.000000000000,-138.000000000000,
559.000000000000,1024.00000000000,
-1243.00000000000,705.000000000000,
-349.000000000000,710.000000000000,
-242.000000000000,-180.000000000000,
-147.000000000000,-317.000000000000,
-390.000000000000,-276.000000000000,
-932.000000000000,-11.0000000000000,
334.000000000000,771.000000000000,
-1077.00000000000,-64.0000000000000,
-621.000000000000,62.0000000000000,
-47.0000000000000,990.000000000000,
-1137.00000000000,221.000000000000,
822.000000000000,-955.000000000000,
725.000000000000,124.000000000000,
-865.000000000000,-506.000000000000,
241.000000000000,-1310.00000000000,
1029.00000000000,405.000000000000,
487.000000000000,79.0000000000000,
295.000000000000,188.000000000000,
-358.000000000000,958.000000000000,
528.000000000000,591.000000000000,
-402.000000000000,183.000000000000,
-1417.00000000000,-70.0000000000000,
755.000000000000,-561.000000000000,
-223.000000000000,-621.000000000000,
266.000000000000,1017.00000000000,
370.000000000000,-280.000000000000,
-688.000000000000,-641.000000000000,
671.000000000000,1352.00000000000,
-516.000000000000,571.000000000000,
447.000000000000,236.000000000000,
1382.00000000000,44.0000000000000,
32.0000000000000,-17.0000000000000,
-279.000000000000,-840.000000000000,
-271.000000000000,-964.000000000000,
73.0000000000000,-349.000000000000,
-103.000000000000,370.000000000000,
862.000000000000,-376.000000000000,
-2.00000000000000,-391.000000000000,
-888.000000000000,616.000000000000,
-342.000000000000,-991.000000000000,
-506.000000000000,-233.000000000000,
530.000000000000,-771.000000000000,
276.000000000000,-233.000000000000,
161.000000000000,1464.00000000000,
297.000000000000,408.000000000000,
404.000000000000,1006.00000000000,
-99.0000000000000,1020.00000000000,
-503.000000000000,61.0000000000000,
319.000000000000,-864.000000000000,
-58.0000000000000,-321.000000000000,
-498.000000000000,81.0000000000000,
-1653.00000000000,-549.000000000000,
36.0000000000000,489.000000000000,
782.000000000000,-9.00000000000000,
36.0000000000000,972.000000000000,
-201.000000000000,944.000000000000,
-1275.00000000000,332.000000000000,
-38.0000000000000,805.000000000000,
-639.000000000000,-717.000000000000,
173.000000000000,149.000000000000,
571.000000000000,520.000000000000,
12.0000000000000,860.000000000000,
392.000000000000,-166.000000000000,
-402.000000000000,178.000000000000,
91.0000000000000,1166.00000000000,
-1346.00000000000,-738.000000000000,
-365.000000000000,-153.000000000000,
50.0000000000000,-1035.00000000000,
-495.000000000000,-900.000000000000,
-215.000000000000,85.0000000000000,
-1119.00000000000,551.000000000000,
761.000000000000,41.0000000000000,
554.000000000000,387.000000000000,
261.000000000000,1585.00000000000,
-61.0000000000000,24.0000000000000,
-524.000000000000,583.000000000000,
612.000000000000,-173.000000000000,
128.000000000000,-1003.00000000000,
379.000000000000,147.000000000000,
169.000000000000,418.000000000000,
177.000000000000,-931.000000000000,
299.000000000000,-671.000000000000,
-381.000000000000,897.000000000000,
59.0000000000000,553.000000000000,
-735.000000000000,894.000000000000,
-1410.00000000000,-361.000000000000,
-369.000000000000,-1283.00000000000,
929.000000000000,-29.0000000000000,
943.000000000000,-268.000000000000,
636.000000000000,-236.000000000000,
278.000000000000,505.000000000000,
-525.000000000000,1416.00000000000,
-322.000000000000,134.000000000000,
-196.000000000000,-392.000000000000,
569.000000000000,642.000000000000,
-212.000000000000,-916.000000000000,
375.000000000000,-747.000000000000,
1346.00000000000,564.000000000000,
87.0000000000000,616.000000000000,
1232.00000000000,200.000000000000,
0.00000000000000,1033.00000000000,
-806.000000000000,-160.000000000000,
753.000000000000,-667.000000000000,
325.000000000000,557.000000000000,
149.000000000000,-1092.00000000000,
103.000000000000,-454.000000000000,
281.000000000000,511.000000000000,
-348.000000000000,994.000000000000,
586.000000000000,379.000000000000,
561.000000000000,270.000000000000,
-1200.00000000000,756.000000000000,
-320.000000000000,-362.000000000000,
23.0000000000000,953.000000000000,
362.000000000000,44.0000000000000,
195.000000000000,68.0000000000000,
1263.00000000000,609.000000000000,
407.000000000000,-55.0000000000000,
-1217.00000000000,604.000000000000,
-288.000000000000,-1153.00000000000,
-203.000000000000,-648.000000000000,
191.000000000000,-9.00000000000000,
-179.000000000000,-778.000000000000,
387.000000000000,-679.000000000000,
-191.000000000000,311.000000000000,
-91.0000000000000,808.000000000000,
1041.00000000000,-295.000000000000,
198.000000000000,157.000000000000,
778.000000000000,-225.000000000000,
-182.000000000000,528.000000000000,
-668.000000000000,1294.00000000000,
354.000000000000,363.000000000000,
-339.000000000000,128.000000000000,
-338.000000000000,696.000000000000,
259.000000000000,-360.000000000000,
886.000000000000,-697.000000000000,
190.000000000000,1190.00000000000,
290.000000000000,-481.000000000000,
-290.000000000000,239.000000000000,
-860.000000000000,-156.000000000000,
682.000000000000,-1244.00000000000,
-145.000000000000,1326.00000000000,
474.000000000000,195.000000000000,
-353.000000000000,408.000000000000,
-1057.00000000000,-224.000000000000,
-782.000000000000,-992.000000000000,
-755.000000000000,278.000000000000,
185.000000000000,-794.000000000000,
-185.000000000000,309.000000000000,
-468.000000000000,361.000000000000,
-510.000000000000,397.000000000000,
691.000000000000,760.000000000000,
394.000000000000,-291.000000000000,
-40.0000000000000,-215.000000000000,
-327.000000000000,-521.000000000000,
116.000000000000,323.000000000000,
-148.000000000000,-52.0000000000000,
-222.000000000000,-325.000000000000,
520.000000000000,1104.00000000000,
-717.000000000000,1098.00000000000,
105.000000000000,1094.00000000000,
-826.000000000000,-132.000000000000,
-1123.00000000000,-75.0000000000000,
235.000000000000,-165.000000000000,
-111.000000000000,-501.000000000000,
143.000000000000,-317.000000000000,
-351.000000000000,-768.000000000000,
809.000000000000,-655.000000000000,
453.000000000000,-678.000000000000,
270.000000000000,204.000000000000,
901.000000000000,-443.000000000000,
-616.000000000000,16.0000000000000,
-369.000000000000,-484.000000000000,
780.000000000000,-1192.00000000000,
681.000000000000,880.000000000000,
-637.000000000000,-119.000000000000,
-495.000000000000,-584.000000000000,
-405.000000000000,382.000000000000,
-650.000000000000,459.000000000000,
-486.000000000000,329.000000000000,
-648.000000000000,-913.000000000000,
862.000000000000,-578.000000000000,
1142.00000000000,588.000000000000,
227.000000000000,-742.000000000000,
695.000000000000,-430.000000000000,
48.0000000000000,467.000000000000,
-630.000000000000,-808.000000000000,
-218.000000000000,60.0000000000000,
68.0000000000000,-609.000000000000,
-187.000000000000,-915.000000000000,
3.00000000000000,880.000000000000,
-5.00000000000000,-290.000000000000,
-473.000000000000,-104.000000000000,
675.000000000000,-725.000000000000,
-423.000000000000,-536.000000000000,
-389.000000000000,-63.0000000000000,
-76.0000000000000,-272.000000000000,
68.0000000000000,1190.00000000000,
-292.000000000000,-188.000000000000,
-804.000000000000,435.000000000000,
956.000000000000,-360.000000000000,
-173.000000000000,-594.000000000000,
657.000000000000,511.000000000000,
-257.000000000000,-509.000000000000,
-985.000000000000,223.000000000000,
451.000000000000,-684.000000000000,
-550.000000000000,-548.000000000000,
-9.00000000000000,403.000000000000,
128.000000000000,622.000000000000,
305.000000000000,28.0000000000000,
-345.000000000000,767.000000000000,
-414.000000000000,521.000000000000,
258.000000000000,-1690.00000000000,
395.000000000000,595.000000000000,
98.0000000000000,298.000000000000,
-761.000000000000,-33.0000000000000,
317.000000000000,810.000000000000,
-339.000000000000,-685.000000000000,
566.000000000000,-302.000000000000,
163.000000000000,-565.000000000000,
-250.000000000000,696.000000000000,
1177.00000000000,342.000000000000,
195.000000000000,-2.00000000000000,
739.000000000000,751.000000000000,
-377.000000000000,-510.000000000000,
280.000000000000,-1060.00000000000,
1204.00000000000,-167.000000000000,
-139.000000000000,702.000000000000,
727.000000000000,-574.000000000000,
386.000000000000,606.000000000000,
768.000000000000,744.000000000000,
-236.000000000000,568.000000000000,
-1278.00000000000,966.000000000000,
-403.000000000000,213.000000000000,
-684.000000000000,679.000000000000,
-676.000000000000,-994.000000000000,
-448.000000000000,-652.000000000000,
628.000000000000,355.000000000000,
619.000000000000,96.0000000000000,
788.000000000000,-78.0000000000000,
547.000000000000,-927.000000000000,
696.000000000000,211.000000000000,
288.000000000000,905.000000000000,
-1067.00000000000,1106.00000000000,
-101.000000000000,298.000000000000,
-653.000000000000,66.0000000000000,
-360.000000000000,-497.000000000000,
422.000000000000,-1643.00000000000,
-362.000000000000,24.0000000000000,
-732.000000000000,-443.000000000000,
-22.0000000000000,-830.000000000000,
726.000000000000,616.000000000000,
-619.000000000000,-103.000000000000,
-562.000000000000,-296.000000000000,
479.000000000000,492.000000000000,
-147.000000000000,173.000000000000,
-418.000000000000,436.000000000000,
-22.0000000000000,669.000000000000,
-208.000000000000,-519.000000000000,
-61.0000000000000,124.000000000000,
-352.000000000000,751.000000000000,
-642.000000000000,-35.0000000000000,
487.000000000000,568.000000000000,
-14.0000000000000,-350.000000000000,
-746.000000000000,-990.000000000000,
-559.000000000000,-670.000000000000,
-581.000000000000,-1092.00000000000,
933.000000000000,-526.000000000000,
398.000000000000,-34.0000000000000,
-122.000000000000,316.000000000000,
331.000000000000,-111.000000000000,
205.000000000000,-32.0000000000000,
19.0000000000000,254.000000000000,
-468.000000000000,610.000000000000,
45.0000000000000,476.000000000000,
250.000000000000,-1073.00000000000,
418.000000000000,276.000000000000,
209.000000000000,512.000000000000,
-71.0000000000000,-143.000000000000,
-382.000000000000,676.000000000000,
528.000000000000,364.000000000000,
-69.0000000000000,455.000000000000,
-1212.00000000000,-456.000000000000,
1629.00000000000,-300.000000000000,
691.000000000000,-298.000000000000,
-159.000000000000,-911.000000000000,
695.000000000000,-1062.00000000000,
-482.000000000000,-319.000000000000,
-573.000000000000,697.000000000000,
-555.000000000000,-1174.00000000000,
197.000000000000,-498.000000000000,
357.000000000000,80.0000000000000,
1003.00000000000,115.000000000000,
195.000000000000,346.000000000000,
-630.000000000000,-249.000000000000,
-45.0000000000000,-188.000000000000,
-751.000000000000,-282.000000000000,
-316.000000000000,886.000000000000,
-398.000000000000,347.000000000000,
335.000000000000,-192.000000000000,
1210.00000000000,747.000000000000,
180.000000000000,478.000000000000,
625.000000000000,-82.0000000000000,
-450.000000000000,239.000000000000,
-621.000000000000,-399.000000000000,
409.000000000000,-270.000000000000,
377.000000000000,1413.00000000000,
399.000000000000,-805.000000000000,
-732.000000000000,-279.000000000000,
18.0000000000000,-127.000000000000,
-338.000000000000,-913.000000000000,
85.0000000000000,952.000000000000,
221.000000000000,479.000000000000,
-668.000000000000,658.000000000000,
-133.000000000000,-527.000000000000,
-535.000000000000,249.000000000000,
13.0000000000000,1344.00000000000,
-432.000000000000,541.000000000000,
-420.000000000000,1167.00000000000,
-600.000000000000,134.000000000000,
-45.0000000000000,480.000000000000,
-709.000000000000,-381.000000000000,
-418.000000000000,-816.000000000000,
1636.00000000000,387.000000000000,
549.000000000000,113.000000000000,
611.000000000000,662.000000000000,
-849.000000000000,385.000000000000,
-1215.00000000000,90.0000000000000,
746.000000000000,-403.000000000000,
-33.0000000000000,17.0000000000000,
-575.000000000000,325.000000000000,
-295.000000000000,421.000000000000,
486.000000000000,760.000000000000,
11.0000000000000,-197.000000000000,
10.0000000000000,-637.000000000000,
476.000000000000,-1261.00000000000,
19.0000000000000,-229.000000000000,
-181.000000000000,-187.000000000000,
-1028.00000000000,-740.000000000000,
283.000000000000,-624.000000000000,
743.000000000000,106.000000000000,
241.000000000000,1802.00000000000,
-295.000000000000,-485.000000000000,
-28.0000000000000,-592.000000000000,
808.000000000000,453.000000000000,
-1223.00000000000,-170.000000000000,
-190.000000000000,-49.0000000000000,
642.000000000000,87.0000000000000,
96.0000000000000,819.000000000000,
159.000000000000,576.000000000000,
-454.000000000000,943.000000000000,
-320.000000000000,774.000000000000,
181.000000000000,12.0000000000000,
756.000000000000,348.000000000000,
911.000000000000,106.000000000000,
437.000000000000,523.000000000000,
-685.000000000000,772.000000000000,
-1096.00000000000,-89.0000000000000,
133.000000000000,-591.000000000000,
772.000000000000,-583.000000000000,
65.0000000000000,-5.00000000000000,
-5.00000000000000,874.000000000000,
-75.0000000000000,-176.000000000000,
-89.0000000000000,-853.000000000000,
1138.00000000000,215.000000000000,
87.0000000000000,-139.000000000000,
-1157.00000000000,140.000000000000,
-305.000000000000,170.000000000000,
-588.000000000000,-727.000000000000,
1092.00000000000,102.000000000000,
158.000000000000,-569.000000000000,
-889.000000000000,140.000000000000,
1181.00000000000,-27.0000000000000,
163.000000000000,719.000000000000,
-830.000000000000,468.000000000000,
-700.000000000000,-1199.00000000000,
98.0000000000000,1233.00000000000,
-1033.00000000000,-499.000000000000,
-98.0000000000000,-107.000000000000,
37.0000000000000,811.000000000000,
-1208.00000000000,-391.000000000000,
665.000000000000,618.000000000000,
-834.000000000000,-1183.00000000000,
-337.000000000000,-953.000000000000,
423.000000000000,510.000000000000,
-913.000000000000,475.000000000000,
-674.000000000000,-672.000000000000,
-120.000000000000,-1417.00000000000,
525.000000000000,-786.000000000000,
182.000000000000,1006.00000000000,
667.000000000000,456.000000000000,
-62.0000000000000,-541.000000000000,
-109.000000000000,264.000000000000,
701.000000000000,-1015.00000000000,
-715.000000000000,550.000000000000,
-240.000000000000,948.000000000000,
-1134.00000000000,-490.000000000000,
-422.000000000000,-714.000000000000,
1106.00000000000,15.0000000000000,
-338.000000000000,201.000000000000,
171.000000000000,-1050.00000000000,
25.0000000000000,704.000000000000,
-349.000000000000,557.000000000000,
754.000000000000,-388.000000000000,
340.000000000000,669.000000000000,
-306.000000000000,-580.000000000000,
656.000000000000,-213.000000000000,
182.000000000000,1072.00000000000,
197.000000000000,490.000000000000,
873.000000000000,-634.000000000000,
-237.000000000000,167.000000000000,
39.0000000000000,919.000000000000,
-1285.00000000000,-387.000000000000,
-333.000000000000,342.000000000000,
873.000000000000,178.000000000000,
-629.000000000000,-148.000000000000,
973.000000000000,-223.000000000000,
-33.0000000000000,138.000000000000,
-1164.00000000000,-101.000000000000,
-782.000000000000,-264.000000000000,
53.0000000000000,271.000000000000,
490.000000000000,-1121.00000000000,
-603.000000000000,748.000000000000,
-406.000000000000,732.000000000000,
-857.000000000000,-173.000000000000,
-19.0000000000000,-692.000000000000,
-33.0000000000000,-1174.00000000000,
544.000000000000,616.000000000000,
602.000000000000,-683.000000000000,
-655.000000000000,768.000000000000,
-136.000000000000,1290.00000000000,
-1194.00000000000,-756.000000000000,
-263.000000000000,-21.0000000000000,
-522.000000000000,538.000000000000,
-867.000000000000,-269.000000000000,
818.000000000000,-936.000000000000,
634.000000000000,-256.000000000000,
-11.0000000000000,66.0000000000000,
230.000000000000,656.000000000000,
1198.00000000000,170.000000000000,
190.000000000000,234.000000000000,
-464.000000000000,989.000000000000,
109.000000000000,-106.000000000000,
-89.0000000000000,6.00000000000000,
-193.000000000000,-278.000000000000,
916.000000000000,473.000000000000,
411.000000000000,684.000000000000,
-705.000000000000,-527.000000000000,
625.000000000000,944.000000000000,
-1176.00000000000,156.000000000000,
-560.000000000000,-14.0000000000000,
926.000000000000,-640.000000000000,
-55.0000000000000,-1043.00000000000,
380.000000000000,1276.00000000000,
-609.000000000000,-137.000000000000,
233.000000000000,-284.000000000000,
-11.0000000000000,285.000000000000,
-471.000000000000,629.000000000000,
277.000000000000,692.000000000000,
58.0000000000000,569.000000000000,
920.000000000000,535.000000000000,
-95.0000000000000,-73.0000000000000,
-137.000000000000,-730.000000000000,
-16.0000000000000,-748.000000000000,
-917.000000000000,-161.000000000000,
-399.000000000000,-507.000000000000,
-30.0000000000000,1159.00000000000,
359.000000000000,523.000000000000,
-350.000000000000,479.000000000000,
138.000000000000,640.000000000000,
-276.000000000000,-1233.00000000000,
-177.000000000000,392.000000000000,
1048.00000000000,121.000000000000,
-716.000000000000,447.000000000000,
-284.000000000000,813.000000000000,
-4.00000000000000,-859.000000000000,
-799.000000000000,-172.000000000000,
-174.000000000000,-256.000000000000,
809.000000000000,-764.000000000000,
609.000000000000,309.000000000000,
320.000000000000,881.000000000000,
593.000000000000,-174.000000000000,
-1056.00000000000,358.000000000000,
-159.000000000000,-476.000000000000,
-410.000000000000,-1141.00000000000,
-616.000000000000,608.000000000000,
1138.00000000000,289.000000000000,
-615.000000000000,700.000000000000,
-165.000000000000,-688.000000000000,
-291.000000000000,-639.000000000000,
16.0000000000000,325.000000000000,
639.000000000000,149.000000000000,
-874.000000000000,307.000000000000,
-591.000000000000,106.000000000000,
-253.000000000000,1409.00000000000,
443.000000000000,169.000000000000,
2.00000000000000,524.000000000000,
564.000000000000,306.000000000000,
75.0000000000000,-301.000000000000,
135.000000000000,1041.00000000000,
377.000000000000,-203.000000000000,
-1397.00000000000,-35.0000000000000,
656.000000000000,-582.000000000000,
402.000000000000,-96.0000000000000,
-177.000000000000,757.000000000000,
-74.0000000000000,127.000000000000,
386.000000000000,575.000000000000,
625.000000000000,59.0000000000000,
-205.000000000000,390.000000000000,
394.000000000000,-1046.00000000000,
-444.000000000000,-264.000000000000,
33.0000000000000,241.000000000000,
-496.000000000000,-857.000000000000,
-467.000000000000,1306.00000000000,
-757.000000000000,-496.000000000000,
-459.000000000000,-456.000000000000,
200.000000000000,871.000000000000,
-1433.00000000000,264.000000000000,
-114.000000000000,-719.000000000000,
-449.000000000000,-1132.00000000000,
676.000000000000,521.000000000000,
983.000000000000,258.000000000000,
-760.000000000000,897.000000000000,
485.000000000000,294.000000000000,
861.000000000000,-132.000000000000,
-140.000000000000,969.000000000000,
-326.000000000000,367.000000000000,
626.000000000000,87.0000000000000,
3.00000000000000,-475.000000000000,
-20.0000000000000,-122.000000000000,
-231.000000000000,-61.0000000000000,
-778.000000000000,492.000000000000,
-449.000000000000,1489.00000000000,
-182.000000000000,17.0000000000000,
-212.000000000000,-305.000000000000,
-1202.00000000000,-635.000000000000,
523.000000000000,-300.000000000000,
1032.00000000000,590.000000000000,
0.00000000000000,769.000000000000,
670.000000000000,438.000000000000,
-202.000000000000,667.000000000000,
400.000000000000,1020.00000000000,
-807.000000000000,-369.000000000000,
-484.000000000000,20.0000000000000,
1411.00000000000,370.000000000000,
-647.000000000000,201.000000000000,
183.000000000000,-958.000000000000,
-235.000000000000,46.0000000000000,
-697.000000000000,209.000000000000,
37.0000000000000,-1142.00000000000,
-124.000000000000,1062.00000000000,
-431.000000000000,165.000000000000,
-1877.00000000000,-403.000000000000,
596.000000000000,-1161.00000000000,
-134.000000000000,-308.000000000000,
-553.000000000000,-247.000000000000,
374.000000000000,-1358.00000000000,
-426.000000000000,1596.00000000000,
-303.000000000000,461.000000000000,
-330.000000000000,-668.000000000000,
1294.00000000000,-752.000000000000,
-256.000000000000,416.000000000000,
722.000000000000,632.000000000000,
344.000000000000,-582.000000000000,
-1108.00000000000,156.000000000000,
480.000000000000,-458.000000000000,
-622.000000000000,1502.00000000000,
-410.000000000000,-290.000000000000,
-710.000000000000,-831.000000000000,
-27.0000000000000,1503.00000000000,
-478.000000000000,456.000000000000,
-205.000000000000,242.000000000000,
1072.00000000000,-306.000000000000,
415.000000000000,-105.000000000000,
1398.00000000000,-174.000000000000,
-629.000000000000,702.000000000000,
-224.000000000000,-375.000000000000,
654.000000000000,-491.000000000000,
-542.000000000000,522.000000000000,
-656.000000000000,-1360.00000000000,
-140.000000000000,353.000000000000,
362.000000000000,838.000000000000,
-1691.00000000000,326.000000000000,
288.000000000000,-265.000000000000,
810.000000000000,-340.000000000000,
-294.000000000000,221.000000000000,
174.000000000000,-1395.00000000000,
-805.000000000000,31.0000000000000,
287.000000000000,139.000000000000,
256.000000000000,-216.000000000000,
-407.000000000000,-461.000000000000,
-551.000000000000,-1076.00000000000,
938.000000000000,-422.000000000000,
686.000000000000,-857.000000000000,
243.000000000000,126.000000000000,
1019.00000000000,-273.000000000000,
227.000000000000,-772.000000000000,
436.000000000000,-207.000000000000,
-398.000000000000,-279.000000000000,
-349.000000000000,89.0000000000000,
360.000000000000,-433.000000000000,
-202.000000000000,84.0000000000000,
-323.000000000000,715.000000000000,
632.000000000000,332.000000000000,
725.000000000000,445.000000000000,
-283.000000000000,-213.000000000000,
818.000000000000,-1296.00000000000,
913.000000000000,66.0000000000000,
-468.000000000000,1640.00000000000,
-1194.00000000000,-106.000000000000,
-1353.00000000000,-680.000000000000,
105.000000000000,-210.000000000000,
493.000000000000,173.000000000000,
-498.000000000000,746.000000000000,
87.0000000000000,-316.000000000000,
454.000000000000,-641.000000000000,
229.000000000000,795.000000000000,
204.000000000000,-280.000000000000,
-266.000000000000,-363.000000000000,
559.000000000000,418.000000000000,
392.000000000000,-343.000000000000,
-595.000000000000,1280.00000000000,
-894.000000000000,57.0000000000000,
-512.000000000000,-1063.00000000000,
342.000000000000,227.000000000000,
751.000000000000,-1129.00000000000,
-258.000000000000,40.0000000000000,
-231.000000000000,384.000000000000,
45.0000000000000,-951.000000000000,
-802.000000000000,355.000000000000,
-235.000000000000,15.0000000000000,
89.0000000000000,446.000000000000,
520.000000000000,456.000000000000,
35.0000000000000,-588.000000000000,
-60.0000000000000,221.000000000000,
62.0000000000000,-793.000000000000,
424.000000000000,-404.000000000000,
310.000000000000,409.000000000000,
-57.0000000000000,979.000000000000,
-252.000000000000,95.0000000000000,
-474.000000000000,-748.000000000000,
992.000000000000,56.0000000000000,
28.0000000000000,-1021.00000000000,
242.000000000000,418.000000000000,
665.000000000000,163.000000000000,
-259.000000000000,-351.000000000000,
-258.000000000000,1137.00000000000,
-220.000000000000,-280.000000000000,
661.000000000000,-867.000000000000,
361.000000000000,-601.000000000000,
762.000000000000,-1223.00000000000,
1102.00000000000,-149.000000000000,
400.000000000000,1211.00000000000,
344.000000000000,1.00000000000000,
-706.000000000000,271.000000000000,
-529.000000000000,707.000000000000,
-442.000000000000,33.0000000000000,
-288.000000000000,209.000000000000,
1556.00000000000,44.0000000000000,
133.000000000000,-79.0000000000000,
-510.000000000000,-149.000000000000,
1050.00000000000,486.000000000000,
-216.000000000000,529.000000000000,
-1450.00000000000,-476.000000000000,
143.000000000000,-571.000000000000,
93.0000000000000,-201.000000000000,
-542.000000000000,1162.00000000000,
-961.000000000000,121.000000000000,
-669.000000000000,-566.000000000000,
247.000000000000,238.000000000000,
14.0000000000000,-962.000000000000,
898.000000000000,521.000000000000,
-375.000000000000,889.000000000000,
-470.000000000000,15.0000000000000,
859.000000000000,2.00000000000000,
-157.000000000000,-15.0000000000000,
567.000000000000,392.000000000000,
-193.000000000000,671.000000000000,
-626.000000000000,396.000000000000,
196.000000000000,-429.000000000000,
446.000000000000,-54.0000000000000,
652.000000000000,-972.000000000000,
-1112.00000000000,-308.000000000000,
-603.000000000000,-430.000000000000,
-559.000000000000,-859.000000000000,
-935.000000000000,-27.0000000000000,
-256.000000000000,-432.000000000000,
284.000000000000,1200.00000000000,
-481.000000000000,172.000000000000,
-955.000000000000,25.0000000000000,
1261.00000000000,636.000000000000,
151.000000000000,135.000000000000,
-915.000000000000,207.000000000000,
-1016.00000000000,-918.000000000000,
-623.000000000000,433.000000000000,
117.000000000000,-25.0000000000000,
41.0000000000000,-1160.00000000000,
513.000000000000,409.000000000000,
-564.000000000000,299.000000000000,
-41.0000000000000,-932.000000000000,
177.000000000000,-559.000000000000,
555.000000000000,775.000000000000,
430.000000000000,-627.000000000000,
-666.000000000000,-322.000000000000,
1083.00000000000,320.000000000000,
685.000000000000,268.000000000000,
-621.000000000000,242.000000000000,
269.000000000000,-1517.00000000000,
716.000000000000,24.0000000000000,
-460.000000000000,576.000000000000,
13.0000000000000,-932.000000000000,
856.000000000000,210.000000000000,
-467.000000000000,1237.00000000000,
-721.000000000000,599.000000000000,
162.000000000000,-290.000000000000,
148.000000000000,-394.000000000000,
-393.000000000000,-660.000000000000,
944.000000000000,-286.000000000000,
826.000000000000,886.000000000000,
635.000000000000,540.000000000000,
615.000000000000,867.000000000000,
-1198.00000000000,686.000000000000,
-930.000000000000,-738.000000000000,
982.000000000000,-216.000000000000,
62.0000000000000,-200.000000000000,
-443.000000000000,-193.000000000000,
601.000000000000,720.000000000000,
1001.00000000000,62.0000000000000,
415.000000000000,758.000000000000,
-697.000000000000,1210.00000000000,
-1363.00000000000,-687.000000000000,
-526.000000000000,-151.000000000000,
425.000000000000,-780.000000000000,
-76.0000000000000,-815.000000000000,
286.000000000000,-56.0000000000000,
-984.000000000000,-321.000000000000,
202.000000000000,887.000000000000,
1083.00000000000,-113.000000000000,
-679.000000000000,1053.00000000000,
-198.000000000000,1245.00000000000,
-1344.00000000000,-125.000000000000,
-50.0000000000000,-321.000000000000,
972.000000000000,-346.000000000000,
713.000000000000,867.000000000000,
636.000000000000,69.0000000000000,
92.0000000000000,-865.000000000000,
1139.00000000000,-791.000000000000,
-743.000000000000,494.000000000000,
-1052.00000000000,247.000000000000,
-478.000000000000,114.000000000000,
-250.000000000000,412.000000000000,
877.000000000000,150.000000000000,
-27.0000000000000,281.000000000000,
320.000000000000,-613.000000000000,
393.000000000000,859.000000000000,
-500.000000000000,1235.00000000000,
-399.000000000000,-30.0000000000000,
396.000000000000,-293.000000000000,
-184.000000000000,371.000000000000,
-437.000000000000,388.000000000000,
8.00000000000000,-1164.00000000000,
-191.000000000000,613.000000000000,
-99.0000000000000,850.000000000000,
-340.000000000000,-1502.00000000000,
97.0000000000000,-84.0000000000000,
-706.000000000000,98.0000000000000,
-1283.00000000000,-638.000000000000,
-280.000000000000,-51.0000000000000,
319.000000000000,270.000000000000,
625.000000000000,381.000000000000,
-1142.00000000000,2.00000000000000,
-420.000000000000,-341.000000000000,
1157.00000000000,136.000000000000,
451.000000000000,-321.000000000000,
831.000000000000,-832.000000000000,
21.0000000000000,187.000000000000,
-473.000000000000,-894.000000000000,
-171.000000000000,-922.000000000000,
-403.000000000000,80.0000000000000,
194.000000000000,-355.000000000000,
654.000000000000,-346.000000000000,
319.000000000000,-1224.00000000000,
995.000000000000,-522.000000000000,
263.000000000000,387.000000000000,
43.0000000000000,-172.000000000000,
-220.000000000000,1034.00000000000,
-707.000000000000,-791.000000000000,
353.000000000000,-989.000000000000,
-433.000000000000,505.000000000000,
439.000000000000,-900.000000000000,
-319.000000000000,-539.000000000000,
-120.000000000000,-831.000000000000,
1075.00000000000,335.000000000000,
-620.000000000000,-241.000000000000,
933.000000000000,-583.000000000000,
765.000000000000,1231.00000000000,
-835.000000000000,-5.00000000000000,
78.0000000000000,-397.000000000000,
-97.0000000000000,647.000000000000,
124.000000000000,-8.00000000000000,
275.000000000000,94.0000000000000,
-312.000000000000,-184.000000000000,
350.000000000000,-1544.00000000000,
216.000000000000,615.000000000000,
-504.000000000000,897.000000000000,
-109.000000000000,-209.000000000000,
1098.00000000000,394.000000000000,
655.000000000000,421.000000000000,
687.000000000000,565.000000000000,
1053.00000000000,583.000000000000,
-739.000000000000,660.000000000000,
-947.000000000000,-348.000000000000,
217.000000000000,-679.000000000000,
540.000000000000,461.000000000000,
552.000000000000,253.000000000000,
172.000000000000,-415.000000000000,
-664.000000000000,309.000000000000,
-645.000000000000,-320.000000000000,
376.000000000000,-1483.00000000000,
236.000000000000,-1052.00000000000,
767.000000000000,-247.000000000000,
811.000000000000,762.000000000000,
-143.000000000000,-257.000000000000,
431.000000000000,-64.0000000000000,
29.0000000000000,829.000000000000,
386.000000000000,338.000000000000,
126.000000000000,310.000000000000,
-75.0000000000000,-180.000000000000,
757.000000000000,351.000000000000,
-69.0000000000000,175.000000000000,
-56.0000000000000,448.000000000000,
53.0000000000000,116.000000000000,
560.000000000000,-637.000000000000,
998.000000000000,477.000000000000,
632.000000000000,-432.000000000000,
-106.000000000000,44.0000000000000,
-223.000000000000,1404.00000000000,
-702.000000000000,-539.000000000000,
-235.000000000000,-388.000000000000,
983.000000000000,191.000000000000,
528.000000000000,496.000000000000,
1194.00000000000,701.000000000000,
-473.000000000000,-242.000000000000,
-1025.00000000000,-168.000000000000,
696.000000000000,-917.000000000000,
163.000000000000,-609.000000000000,
-253.000000000000,-367.000000000000,
901.000000000000,225.000000000000,
259.000000000000,850.000000000000,
-915.000000000000,-244.000000000000,
480.000000000000,-231.000000000000,
141.000000000000,-218.000000000000,
-102.000000000000,-264.000000000000,
515.000000000000,-169.000000000000,
590.000000000000,550.000000000000,
631.000000000000,584.000000000000,
-923.000000000000,108.000000000000,
-107.000000000000,-526.000000000000,
-397.000000000000,-869.000000000000,
-191.000000000000,814.000000000000,
1111.00000000000,173.000000000000,
-920.000000000000,653.000000000000,
-505.000000000000,1145.00000000000,
-496.000000000000,389.000000000000,
-887.000000000000,-340.000000000000,
-363.000000000000,-795.000000000000,
-223.000000000000,561.000000000000,
272.000000000000,64.0000000000000,
786.000000000000,427.000000000000,
501.000000000000,475.000000000000,
-139.000000000000,271.000000000000,
476.000000000000,912.000000000000,
-423.000000000000,-185.000000000000,
-409.000000000000,-551.000000000000,
434.000000000000,-780.000000000000,
22.0000000000000,-184.000000000000,
-724.000000000000,-34.0000000000000,
-1241.00000000000,-696.000000000000,
-492.000000000000,-632.000000000000,
-657.000000000000,-875.000000000000,
982.000000000000,-412.000000000000,
630.000000000000,-870.000000000000,
-973.000000000000,209.000000000000,
817.000000000000,-193.000000000000,
1016.00000000000,215.000000000000,
907.000000000000,1005.00000000000,
-189.000000000000,-1050.00000000000,
10.0000000000000,-101.000000000000,
-334.000000000000,-777.000000000000,
-59.0000000000000,-74.0000000000000,
1196.00000000000,789.000000000000,
-615.000000000000,596.000000000000,
840.000000000000,318.000000000000,
-153.000000000000,-303.000000000000,
-1153.00000000000,371.000000000000,
576.000000000000,-597.000000000000,
-266.000000000000,773.000000000000,
-611.000000000000,934.000000000000,
483.000000000000,-141.000000000000,
182.000000000000,1188.00000000000,
-651.000000000000,701.000000000000,
-541.000000000000,-371.000000000000,
-651.000000000000,-533.000000000000,
837.000000000000,-260.000000000000,
378.000000000000,-593.000000000000,
-691.000000000000,-690.000000000000,
-135.000000000000,261.000000000000,
-466.000000000000,832.000000000000,
-616.000000000000,1198.00000000000,
65.0000000000000,-1.00000000000000,
770.000000000000,211.000000000000,
-441.000000000000,1026.00000000000,
-505.000000000000,390.000000000000,
89.0000000000000,480.000000000000,
-152.000000000000,361.000000000000,
916.000000000000,-96.0000000000000,
-390.000000000000,-381.000000000000,
-610.000000000000,792.000000000000,
288.000000000000,613.000000000000,
-825.000000000000,-141.000000000000,
-144.000000000000,-394.000000000000,
400.000000000000,-137.000000000000,
45.0000000000000,273.000000000000,
175.000000000000,-514.000000000000,
-269.000000000000,205.000000000000,
-663.000000000000,-273.000000000000,
203.000000000000,-1333.00000000000,
-157.000000000000,-329.000000000000,
-656.000000000000,646.000000000000,
41.0000000000000,796.000000000000,
-411.000000000000,-397.000000000000,
-230.000000000000,-3.00000000000000,
-91.0000000000000,-732.000000000000,
770.000000000000,-391.000000000000,
763.000000000000,749.000000000000,
-373.000000000000,-1072.00000000000,
98.0000000000000,254.000000000000,
48.0000000000000,732.000000000000,
113.000000000000,61.0000000000000,
-667.000000000000,756.000000000000,
-488.000000000000,906.000000000000,
-262.000000000000,-182.000000000000,
-1419.00000000000,-461.000000000000,
278.000000000000,335.000000000000,
677.000000000000,-138.000000000000,
-279.000000000000,-191.000000000000,
-139.000000000000,-1022.00000000000,
411.000000000000,-828.000000000000,
541.000000000000,-899.000000000000,
-696.000000000000,86.0000000000000,
88.0000000000000,1051.00000000000,
-188.000000000000,-357.000000000000,
10.0000000000000,469.000000000000,
988.000000000000,823.000000000000,
-1161.00000000000,318.000000000000,
-642.000000000000,241.000000000000,
209.000000000000,179.000000000000,
171.000000000000,-1035.00000000000,
435.000000000000,-352.000000000000,
1133.00000000000,953.000000000000,
180.000000000000,-856.000000000000,
-1004.00000000000,241.000000000000,
194.000000000000,-158.000000000000,
313.000000000000,-58.0000000000000,
-110.000000000000,1328.00000000000,
-873.000000000000,69.0000000000000,
-171.000000000000,963.000000000000,
-1157.00000000000,-27.0000000000000,
-1277.00000000000,-599.000000000000,
246.000000000000,-499.000000000000,
-567.000000000000,-394.000000000000,
294.000000000000,615.000000000000,
-513.000000000000,-244.000000000000,
-415.000000000000,-742.000000000000,
1009.00000000000,-11.0000000000000,
510.000000000000,284.000000000000,
33.0000000000000,-850.000000000000,
470.000000000000,325.000000000000,
1317.00000000000,243.000000000000,
-630.000000000000,-637.000000000000,
-113.000000000000,233.000000000000,
850.000000000000,-730.000000000000,
8.00000000000000,823.000000000000,
195.000000000000,300.000000000000,
259.000000000000,-25.0000000000000,
1071.00000000000,-361.000000000000,
-787.000000000000,-576.000000000000,
258.000000000000,633.000000000000,
-54.0000000000000,-1427.00000000000,
66.0000000000000,520.000000000000,
1118.00000000000,-400.000000000000,
-1109.00000000000,-277.000000000000,
36.0000000000000,1006.00000000000,
36.0000000000000,-1398.00000000000,
1136.00000000000,834.000000000000,
817.000000000000,1168.00000000000,
-1089.00000000000,171.000000000000,
-459.000000000000,388.000000000000,
-440.000000000000,-258.000000000000,
-312.000000000000,-616.000000000000,
91.0000000000000,104.000000000000,
295.000000000000,-281.000000000000,
-592.000000000000,67.0000000000000,
-80.0000000000000,1067.00000000000,
979.000000000000,-7.00000000000000,
130.000000000000,998.000000000000,
-395.000000000000,475.000000000000,
-69.0000000000000,-211.000000000000,
1014.00000000000,334.000000000000,
233.000000000000,-40.0000000000000,
618.000000000000,542.000000000000,
594.000000000000,-633.000000000000,
3.00000000000000,-274.000000000000,
1010.00000000000,-83.0000000000000,
-1006.00000000000,-722.000000000000,
-172.000000000000,-149.000000000000,
1449.00000000000,-126.000000000000,
154.000000000000,1491.00000000000,
-647.000000000000,1096.00000000000,
-924.000000000000,687.000000000000,
-360.000000000000,466.000000000000,
210.000000000000,-777.000000000000,
69.0000000000000,-679.000000000000,
-321.000000000000,-177.000000000000,
825.000000000000,211.000000000000,
-78.0000000000000,-462.000000000000,
-952.000000000000,419.000000000000,
-519.000000000000,-184.000000000000,
-412.000000000000,-1385.00000000000,
466.000000000000,230.000000000000,
-558.000000000000,687.000000000000,
23.0000000000000,980.000000000000,
376.000000000000,-475.000000000000,
-672.000000000000,-34.0000000000000,
-99.0000000000000,998.000000000000,
134.000000000000,-383.000000000000,
306.000000000000,216.000000000000,
490.000000000000,441.000000000000,
69.0000000000000,115.000000000000,
-1124.00000000000,279.000000000000,
-1132.00000000000,-227.000000000000,
-767.000000000000,-1097.00000000000,
-18.0000000000000,-276.000000000000,
1089.00000000000,-444.000000000000,
-291.000000000000,-825.000000000000,
22.0000000000000,-433.000000000000,
661.000000000000,-1018.00000000000,
368.000000000000,369.000000000000,
471.000000000000,100.000000000000,
-324.000000000000,-132.000000000000,
567.000000000000,406.000000000000,
-998.000000000000,-363.000000000000,
-726.000000000000,-290.000000000000,
1346.00000000000,-844.000000000000,
233.000000000000,294.000000000000,
807.000000000000,262.000000000000,
770.000000000000,309.000000000000,
311.000000000000,1103.00000000000,
-478.000000000000,958.000000000000,
345.000000000000,39.0000000000000,
619.000000000000,93.0000000000000,
-669.000000000000,1687.00000000000,
-622.000000000000,453.000000000000,
-819.000000000000,-240.000000000000,
-30.0000000000000,-416.000000000000,
-688.000000000000,-848.000000000000,
-642.000000000000,-396.000000000000,
220.000000000000,146.000000000000,
-507.000000000000,234.000000000000,
-442.000000000000,-957.000000000000,
-161.000000000000,-86.0000000000000,
798.000000000000,697.000000000000,
790.000000000000,45.0000000000000,
391.000000000000,-127.000000000000,
391.000000000000,166.000000000000,
-230.000000000000,-9.00000000000000,
-784.000000000000,-623.000000000000,
-900.000000000000,-110.000000000000,
625.000000000000,276.000000000000,
561.000000000000,617.000000000000,
904.000000000000,303.000000000000,
311.000000000000,748.000000000000,
-467.000000000000,1027.00000000000,
622.000000000000,-822.000000000000,
-301.000000000000,-505.000000000000,
73.0000000000000,-324.000000000000,
-224.000000000000,633.000000000000,
-677.000000000000,505.000000000000,
-556.000000000000,-839.000000000000,
-357.000000000000,817.000000000000,
326.000000000000,-781.000000000000,
434.000000000000,-372.000000000000,
272.000000000000,1649.00000000000,
-334.000000000000,328.000000000000,
494.000000000000,-461.000000000000,
-131.000000000000,57.0000000000000,
704.000000000000,645.000000000000,
1039.00000000000,336.000000000000,
-364.000000000000,1157.00000000000,
484.000000000000,338.000000000000,
-94.0000000000000,-172.000000000000,
404.000000000000,-143.000000000000,
436.000000000000,-1529.00000000000,
377.000000000000,364.000000000000,
575.000000000000,1242.00000000000,
-1114.00000000000,263.000000000000,
-788.000000000000,-606.000000000000,
-24.0000000000000,-570.000000000000,
358.000000000000,68.0000000000000,
721.000000000000,456.000000000000,
791.000000000000,1053.00000000000,
-454.000000000000,327.000000000000,
-398.000000000000,-340.000000000000,
-53.0000000000000,-1306.00000000000,
-1066.00000000000,-196.000000000000,
814.000000000000,-275.000000000000,
-12.0000000000000,-931.000000000000,
-797.000000000000,1284.00000000000,
228.000000000000,79.0000000000000,
385.000000000000,-212.000000000000,
-220.000000000000,-497.000000000000,
-891.000000000000,141.000000000000,
702.000000000000,553.000000000000,
-633.000000000000,-969.000000000000,
-316.000000000000,1024.00000000000,
-77.0000000000000,-830.000000000000,
-618.000000000000,-1046.00000000000,
798.000000000000,44.0000000000000,
271.000000000000,881.000000000000,
-226.000000000000,1148.00000000000,
-1108.00000000000,-744.000000000000,
185.000000000000,109.000000000000,
-494.000000000000,-867.000000000000,
-486.000000000000,-267.000000000000,
996.000000000000,-54.0000000000000,
-92.0000000000000,409.000000000000,
65.0000000000000,522.000000000000,
-1332.00000000000,-517.000000000000,
331.000000000000,362.000000000000,
624.000000000000,-33.0000000000000,
90.0000000000000,621.000000000000,
1168.00000000000,-251.000000000000,
-605.000000000000,517.000000000000,
867.000000000000,100.000000000000,
-503.000000000000,-584.000000000000,
-935.000000000000,-104.000000000000,
1189.00000000000,-1678.00000000000,
495.000000000000,93.0000000000000,
803.000000000000,774.000000000000,
122.000000000000,-129.000000000000,
-797.000000000000,-233.000000000000,
-233.000000000000,469.000000000000,
865.000000000000,362.000000000000,
448.000000000000,-807.000000000000,
411.000000000000,-141.000000000000,
462.000000000000,-810.000000000000,
167.000000000000,-906.000000000000,
-141.000000000000,26.0000000000000,
-125.000000000000,-535.000000000000,
-122.000000000000,-658.000000000000,
-647.000000000000,-367.000000000000,
783.000000000000,-211.000000000000,
606.000000000000,-34.0000000000000,
-180.000000000000,-132.000000000000,
-176.000000000000,-774.000000000000,
-774.000000000000,-325.000000000000,
229.000000000000,207.000000000000,
710.000000000000,-166.000000000000,
230.000000000000,899.000000000000,
-373.000000000000,63.0000000000000,
-213.000000000000,78.0000000000000,
589.000000000000,239.000000000000,
-28.0000000000000,-132.000000000000,
54.0000000000000,334.000000000000,
-180.000000000000,-1186.00000000000,
550.000000000000,-161.000000000000,
180.000000000000,668.000000000000,
-1254.00000000000,265.000000000000,
-500.000000000000,-289.000000000000,
240.000000000000,-923.000000000000,
599.000000000000,-236.000000000000,
576.000000000000,-240.000000000000,
634.000000000000,-139.000000000000,
140.000000000000,822.000000000000,
195.000000000000,1047.00000000000,
509.000000000000,240.000000000000,
-678.000000000000,846.000000000000,
-890.000000000000,762.000000000000,
-17.0000000000000,-28.0000000000000,
586.000000000000,342.000000000000,
490.000000000000,-681.000000000000,
572.000000000000,-593.000000000000,
509.000000000000,153.000000000000,
1.00000000000000,-52.0000000000000,
402.000000000000,270.000000000000,
342.000000000000,674.000000000000,
906.000000000000,483.000000000000,
30.0000000000000,80.0000000000000,
-734.000000000000,1270.00000000000,
32.0000000000000,136.000000000000,
-1329.00000000000,-883.000000000000,
239.000000000000,-248.000000000000,
607.000000000000,349.000000000000,
-701.000000000000,1108.00000000000,
252.000000000000,-182.000000000000,
250.000000000000,492.000000000000,
-247.000000000000,1008.00000000000,
-467.000000000000,-209.000000000000,
373.000000000000,-446.000000000000,
619.000000000000,452.000000000000,
933.000000000000,-130.000000000000,
91.0000000000000,-699.000000000000,
-449.000000000000,31.0000000000000,
924.000000000000,-995.000000000000,
121.000000000000,-988.000000000000,
715.000000000000,310.000000000000,
532.000000000000,634.000000000000,
-523.000000000000,-308.000000000000,
438.000000000000,385.000000000000,
345.000000000000,344.000000000000,
148.000000000000,-1286.00000000000,
1019.00000000000,529.000000000000,
789.000000000000,574.000000000000,
-1106.00000000000,395.000000000000,
-252.000000000000,1265.00000000000,
-471.000000000000,-727.000000000000,
-178.000000000000,-238.000000000000,
1132.00000000000,14.0000000000000,
-586.000000000000,22.0000000000000,
383.000000000000,-56.0000000000000,
-214.000000000000,-288.000000000000,
-1153.00000000000,42.0000000000000,
-273.000000000000,-1505.00000000000,
702.000000000000,-864.000000000000,
262.000000000000,-223.000000000000,
-664.000000000000,871.000000000000,
-2.00000000000000,799.000000000000,
-123.000000000000,50.0000000000000,
623.000000000000,442.000000000000,
285.000000000000,-165.000000000000,
-59.0000000000000,-26.0000000000000,
684.000000000000,-476.000000000000,
927.000000000000,421.000000000000,
323.000000000000,628.000000000000,
-306.000000000000,-768.000000000000,
676.000000000000,-181.000000000000,
281.000000000000,-144.000000000000,
-338.000000000000,-87.0000000000000,
-365.000000000000,238.000000000000,
-725.000000000000,-230.000000000000,
480.000000000000,-474.000000000000,
1183.00000000000,644.000000000000,
564.000000000000,700.000000000000,
96.0000000000000,-840.000000000000,
659.000000000000,-547.000000000000,
357.000000000000,594.000000000000,
85.0000000000000,396.000000000000,
603.000000000000,-1016.00000000000,
229.000000000000,9.00000000000000,
320.000000000000,411.000000000000,
292.000000000000,-205.000000000000,
-24.0000000000000,1137.00000000000,
-910.000000000000,-336.000000000000,
52.0000000000000,-506.000000000000,
638.000000000000,929.000000000000,
-1390.00000000000,170.000000000000,
280.000000000000,-377.000000000000,
912.000000000000,473.000000000000,
-904.000000000000,1068.00000000000,
-319.000000000000,-751.000000000000,
440.000000000000,-711.000000000000,
581.000000000000,311.000000000000,
526.000000000000,492.000000000000,
-873.000000000000,325.000000000000,
-251.000000000000,-701.000000000000,
641.000000000000,577.000000000000,
-1079.00000000000,197.000000000000,
16.0000000000000,-783.000000000000,
555.000000000000,-920.000000000000,
-102.000000000000,-44.0000000000000,
448.000000000000,1338.00000000000,
-214.000000000000,655.000000000000,
812.000000000000,257.000000000000,
-112.000000000000,-420.000000000000,
-513.000000000000,-801.000000000000,
558.000000000000,-367.000000000000,
-908.000000000000,236.000000000000,
715.000000000000,-607.000000000000,
-141.000000000000,220.000000000000,
-547.000000000000,665.000000000000,
1068.00000000000,-401.000000000000,
667.000000000000,1302.00000000000,
714.000000000000,-521.000000000000,
-626.000000000000,-302.000000000000,
-160.000000000000,346.000000000000,
-859.000000000000,-1278.00000000000,
-867.000000000000,-223.000000000000,
1027.00000000000,-435.000000000000,
536.000000000000,574.000000000000,
38.0000000000000,1216.00000000000,
307.000000000000,370.000000000000,
-755.000000000000,332.000000000000,
-415.000000000000,-1095.00000000000,
659.000000000000,-636.000000000000,
-486.000000000000,1004.00000000000,
-56.0000000000000,26.0000000000000,
-162.000000000000,109.000000000000,
-990.000000000000,102.000000000000,
-5.00000000000000,-937.000000000000,
521.000000000000,752.000000000000,
55.0000000000000,743.000000000000,
167.000000000000,-459.000000000000,
33.0000000000000,401.000000000000,
-835.000000000000,208.000000000000,
-151.000000000000,204.000000000000,
860.000000000000,-12.0000000000000,
91.0000000000000,-184.000000000000,
1054.00000000000,521.000000000000,
407.000000000000,406.000000000000,
-1474.00000000000,331.000000000000,
-624.000000000000,-1002.00000000000,
-224.000000000000,-668.000000000000,
138.000000000000,1081.00000000000,
-718.000000000000,447.000000000000,
-204.000000000000,-790.000000000000,
800.000000000000,244.000000000000,
273.000000000000,84.0000000000000,
261.000000000000,-466.000000000000,
381.000000000000,-43.0000000000000,
1100.00000000000,31.0000000000000,
-724.000000000000,518.000000000000,
-290.000000000000,-397.000000000000,
1333.00000000000,154.000000000000,
-655.000000000000,567.000000000000,
-249.000000000000,62.0000000000000,
624.000000000000,1138.00000000000,
-581.000000000000,249.000000000000,
-66.0000000000000,-321.000000000000,
-118.000000000000,891.000000000000,
-637.000000000000,424.000000000000,
1252.00000000000,-41.0000000000000,
246.000000000000,48.0000000000000,
-1042.00000000000,491.000000000000,
-211.000000000000,492.000000000000,
-1246.00000000000,771.000000000000,
27.0000000000000,-84.0000000000000,
-486.000000000000,-819.000000000000,
-695.000000000000,361.000000000000,
14.0000000000000,67.0000000000000,
-974.000000000000,772.000000000000,
1053.00000000000,628.000000000000,
353.000000000000,-255.000000000000,
-561.000000000000,365.000000000000,
-10.0000000000000,596.000000000000,
75.0000000000000,-628.000000000000,
946.000000000000,-584.000000000000,
582.000000000000,-286.000000000000,
629.000000000000,-801.000000000000,
351.000000000000,899.000000000000,
563.000000000000,810.000000000000,
-140.000000000000,304.000000000000,
105.000000000000,-67.0000000000000,
432.000000000000,228.000000000000,
351.000000000000,1067.00000000000,
832.000000000000,-86.0000000000000,
-1072.00000000000,140.000000000000,
-124.000000000000,-619.000000000000,
-478.000000000000,-370.000000000000,
276.000000000000,727.000000000000,
693.000000000000,-414.000000000000,
-1403.00000000000,790.000000000000,
-435.000000000000,-242.000000000000,
52.0000000000000,-183.000000000000,
544.000000000000,149.000000000000,
371.000000000000,-563.000000000000,
925.000000000000,990.000000000000,
843.000000000000,220.000000000000,
596.000000000000,673.000000000000,
662.000000000000,600.000000000000,
-47.0000000000000,-155.000000000000,
357.000000000000,380.000000000000,
140.000000000000,489.000000000000,
-393.000000000000,1262.00000000000,
-832.000000000000,417.000000000000,
-658.000000000000,-689.000000000000,
-507.000000000000,-8.00000000000000,
3.00000000000000,618.000000000000,
-171.000000000000,-404.000000000000,
102.000000000000,-807.000000000000,
207.000000000000,-604.000000000000,
-824.000000000000,-903.000000000000,
249.000000000000,357.000000000000,
601.000000000000,-76.0000000000000,
-151.000000000000,-263.000000000000,
-437.000000000000,-165.000000000000,
-311.000000000000,-581.000000000000,
182.000000000000,1094.00000000000,
-596.000000000000,-268.000000000000,
571.000000000000,-952.000000000000,
1239.00000000000,281.000000000000,
-113.000000000000,291.000000000000,
174.000000000000,-1077.00000000000,
170.000000000000,-870.000000000000,
1039.00000000000,-29.0000000000000,
354.000000000000,535.000000000000,
467.000000000000,974.000000000000,
240.000000000000,-577.000000000000,
-1119.00000000000,42.0000000000000,
998.000000000000,-381.000000000000,
-188.000000000000,-608.000000000000,
-61.0000000000000,-559.000000000000,
210.000000000000,-1199.00000000000,
-372.000000000000,-34.0000000000000,
578.000000000000,482.000000000000,
-731.000000000000,981.000000000000,
-862.000000000000,-100.000000000000,
-351.000000000000,302.000000000000,
66.0000000000000,992.000000000000,
-301.000000000000,560.000000000000,
-916.000000000000,1343.00000000000,
-362.000000000000,309.000000000000,
394.000000000000,521.000000000000,
-408.000000000000,263.000000000000,
-152.000000000000,-254.000000000000,
1481.00000000000,437.000000000000,
8.00000000000000,-610.000000000000,
555.000000000000,-558.000000000000,
464.000000000000,-685.000000000000,
-200.000000000000,312.000000000000,
630.000000000000,-410.000000000000,
-30.0000000000000,-154.000000000000,
897.000000000000,143.000000000000,
500.000000000000,-759.000000000000,
739.000000000000,1251.00000000000,
-369.000000000000,479.000000000000,
-1324.00000000000,-136.000000000000,
322.000000000000,-443.000000000000,
-952.000000000000,220.000000000000,
-537.000000000000,919.000000000000,
-819.000000000000,532.000000000000,
-631.000000000000,922.000000000000,
244.000000000000,427.000000000000,
-763.000000000000,136.000000000000,
-482.000000000000,-1341.00000000000,
-87.0000000000000,-1204.00000000000,
-99.0000000000000,-771.000000000000,
-755.000000000000,-595.000000000000,
-263.000000000000,259.000000000000,
-324.000000000000,-511.000000000000,
387.000000000000,663.000000000000,
1049.00000000000,-250.000000000000,
684.000000000000,-337.000000000000,
602.000000000000,961.000000000000,
-544.000000000000,522.000000000000,
-142.000000000000,670.000000000000,
-971.000000000000,-221.000000000000,
-20.0000000000000,-17.0000000000000,
824.000000000000,-671.000000000000,
-1149.00000000000,-264.000000000000,
-275.000000000000,908.000000000000,
-318.000000000000,188.000000000000,
-715.000000000000,248.000000000000,
-283.000000000000,412.000000000000,
-684.000000000000,-45.0000000000000,
274.000000000000,-373.000000000000,
1052.00000000000,1347.00000000000,
-289.000000000000,372.000000000000,
-128.000000000000,-1069.00000000000,
1088.00000000000,257.000000000000,
-947.000000000000,475.000000000000,
-178.000000000000,798.000000000000,
246.000000000000,211.000000000000,
-1316.00000000000,148.000000000000,
669.000000000000,-840.000000000000,
-4.00000000000000,208.000000000000,
-613.000000000000,1176.00000000000,
-490.000000000000,-1351.00000000000,
-333.000000000000,480.000000000000,
-410.000000000000,332.000000000000,
581.000000000000,-101.000000000000,
1641.00000000000,531.000000000000,
-1136.00000000000,-47.0000000000000,
-170.000000000000,-763.000000000000,
604.000000000000,-1062.00000000000,
281.000000000000,151.000000000000,
-197.000000000000,-589.000000000000,
-1184.00000000000,26.0000000000000,
603.000000000000,456.000000000000,
-235.000000000000,410.000000000000,
428.000000000000,-497.000000000000,
222.000000000000,-614.000000000000,
310.000000000000,-69.0000000000000,
669.000000000000,-1076.00000000000,
-923.000000000000,701.000000000000,
579.000000000000,60.0000000000000,
-13.0000000000000,140.000000000000,
467.000000000000,-202.000000000000,
-83.0000000000000,-1109.00000000000,
262.000000000000,364.000000000000,
573.000000000000,-968.000000000000,
-1036.00000000000,106.000000000000,
295.000000000000,563.000000000000,
125.000000000000,-514.000000000000,
1256.00000000000,-49.0000000000000,
235.000000000000,1026.00000000000,
-1188.00000000000,490.000000000000,
68.0000000000000,-532.000000000000,
198.000000000000,42.0000000000000,
-57.0000000000000,95.0000000000000,
-642.000000000000,715.000000000000,
-488.000000000000,219.000000000000,
-682.000000000000,-475.000000000000,
5.00000000000000,-498.000000000000,
65.0000000000000,-155.000000000000,
-247.000000000000,838.000000000000,
-185.000000000000,679.000000000000,
-1314.00000000000,81.0000000000000,
387.000000000000,-564.000000000000,
1055.00000000000,-216.000000000000,
116.000000000000,48.0000000000000,
1143.00000000000,-142.000000000000,
383.000000000000,-71.0000000000000,
-814.000000000000,352.000000000000,
-192.000000000000,167.000000000000,
-783.000000000000,-350.000000000000,
-915.000000000000,-579.000000000000,
416.000000000000,-598.000000000000,
783.000000000000,415.000000000000,
607.000000000000,478.000000000000,
573.000000000000,438.000000000000,
134.000000000000,83.0000000000000,
-694.000000000000,-173.000000000000,
329.000000000000,452.000000000000,
751.000000000000,192.000000000000,
123.000000000000,441.000000000000,
-400.000000000000,559.000000000000,
-896.000000000000,-328.000000000000,
229.000000000000,-1433.00000000000,
1301.00000000000,-762.000000000000,
-259.000000000000,705.000000000000,
-470.000000000000,367.000000000000,
-1024.00000000000,99.0000000000000,
-873.000000000000,-732.000000000000,
1164.00000000000,-268.000000000000,
-118.000000000000,929.000000000000,
507.000000000000,338.000000000000,
-424.000000000000,1008.00000000000,
-148.000000000000,-23.0000000000000,
-14.0000000000000,49.0000000000000,
-993.000000000000,484.000000000000,
1320.00000000000,-482.000000000000,
91.0000000000000,-42.0000000000000,
35.0000000000000,-598.000000000000,
707.000000000000,317.000000000000,
474.000000000000,-119.000000000000,
454.000000000000,-1209.00000000000,
411.000000000000,22.0000000000000,
457.000000000000,-1284.00000000000,
-310.000000000000,627.000000000000,
-535.000000000000,1409.00000000000,
216.000000000000,157.000000000000,
97.0000000000000,969.000000000000,
-341.000000000000,-1084.00000000000,
1335.00000000000,602.000000000000,
28.0000000000000,-22.0000000000000,
436.000000000000,-896.000000000000,
992.000000000000,1234.00000000000,
-1383.00000000000,607.000000000000,
-891.000000000000,-89.0000000000000,
-952.000000000000,-477.000000000000,
345.000000000000,-270.000000000000,
601.000000000000,-100.000000000000,
-682.000000000000,1417.00000000000,
-668.000000000000,227.000000000000,
-1053.00000000000,-313.000000000000,
870.000000000000,710.000000000000,
105.000000000000,261.000000000000,
-34.0000000000000,429.000000000000,
1304.00000000000,-125.000000000000,
-771.000000000000,742.000000000000,
-789.000000000000,410.000000000000,
-116.000000000000,356.000000000000,
-269.000000000000,347.000000000000,
-638.000000000000,229.000000000000,
568.000000000000,846.000000000000,
544.000000000000,-523.000000000000,
330.000000000000,146.000000000000,
614.000000000000,787.000000000000,
-1170.00000000000,219.000000000000,
-571.000000000000,41.0000000000000,
379.000000000000,-198.000000000000,
748.000000000000,2.00000000000000,
384.000000000000,331.000000000000,
-743.000000000000,-163.000000000000,
-349.000000000000,-1010.00000000000,
-231.000000000000,-711.000000000000,
-804.000000000000,-554.000000000000,
287.000000000000,-249.000000000000,
1084.00000000000,662.000000000000,
885.000000000000,997.000000000000,
107.000000000000,301.000000000000,
-283.000000000000,-339.000000000000,
768.000000000000,760.000000000000,
-639.000000000000,545.000000000000,
-783.000000000000,-1252.00000000000,
378.000000000000,-375.000000000000,
-979.000000000000,180.000000000000,
-889.000000000000,-75.0000000000000};
