shortreal out[256] = '{0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
2.66509092572420e-10,
4.61373126370290e-08,
8.88102675844493e-08,
2.40444421706343e-07,
3.75227330096095e-07,
7.02720228673570e-07,
9.68885160546051e-07,
1.28994133774540e-06,
1.44176726735168e-06,
1.16348769552133e-06,
5.54416374143329e-07,
-1.50671303345007e-06,
-4.11884411732899e-06,
-9.95987466012593e-06,
-1.65829023899278e-05,
-2.92648292088415e-05,
-4.32401866419241e-05,
-6.28012639936060e-05,
-8.24869930511341e-05,
-0.000109443266410381,
-0.000135262962430716,
-0.000169655118952505,
-0.000196373308426701,
-0.000232294376473874,
-0.000268995063379407,
-0.000319092359859496,
-0.000365189247531816,
-0.000412089983001351,
-0.000462468044133857,
-0.000483716867165640,
-0.000517295440658927,
-0.000480718270409852,
-0.000459422910353169,
-0.000377413205569610,
-0.000303582055494189,
-0.000138340023113415,
3.89154592994601e-05,
0.000345375941833481,
0.000707449391484261,
0.00133225915487856,
0.00203267880715430,
0.000826355768367648,
-0.000163685297593474,
0.000442691496573389,
0.00152463337872177,
0.00253183161839843,
0.00245912885293365,
0.00145507056731731,
-0.00277410028502345,
-0.00927543826401234,
-0.0150782559067011,
-0.0211231745779514,
-0.0273839086294174,
-0.0330593287944794,
-0.0381380058825016,
-0.0401630885899067,
-0.0425003059208393,
-0.0487441942095757,
-0.0525458492338657,
-0.0556293204426765,
-0.0593254901468754,
-0.0634186938405037,
-0.0680719092488289,
-0.0721101686358452,
-0.0783602744340897,
-0.0832021981477737,
-0.0897725224494934,
-0.0973846688866615,
-0.102064333856106,
-0.106065139174461,
-0.109658837318420,
-0.112591877579689,
-0.112577855587006,
-0.115370012819767,
-0.120329752564430,
-0.123550817370415,
-0.129484817385674,
-0.137580111622810,
-0.144542515277863,
-0.148416638374329,
-0.152123183012009,
-0.154995545744896,
-0.157224565744400,
-0.161946207284927,
-0.164249628782272,
-0.164953604340553,
-0.166232600808144,
-0.165594831109047,
-0.164933457970619,
-0.165674477815628,
-0.165187105536461,
-0.164969965815544,
-0.168054789304733,
-0.172671675682068,
-0.180064320564270,
-0.190728619694710,
-0.205018892884254,
-0.221605673432350,
-0.236788377165794,
-0.251209467649460,
-0.266243666410446,
-0.282457083463669,
-0.299866735935211,
-0.321500808000565,
-0.342596441507340,
-0.364256680011749,
-0.389486312866211,
-0.411321371793747,
-0.434028476476669,
-0.458701789379120,
-0.485420435667038,
-0.513122558593750,
-0.539874434471130,
-0.569842636585236,
-0.599001765251160,
-0.625391304492950,
-0.651307046413422,
-0.677643716335297,
-0.707461118698120,
-0.737938582897186,
-0.765931665897369,
-0.796017229557037,
-0.827176332473755,
-0.856641054153442,
-0.886234462261200,
-0.918056726455689,
-0.951689720153809,
-0.984218776226044,
-1.01964545249939,
-1.05308079719543,
-1.08798730373383,
-1.12210524082184,
-1.16020810604095,
-1.19282150268555,
-1.23325490951538,
-1.26595175266266,
-1.29865431785584,
-1.33520233631134,
-1.35154008865356,
-1.40526676177979,
-1.40052199363709,
-1.48026192188263,
-1.43507218360901,
-1.55214452743530,
-1.52207088470459,
-1.65377736091614,
-1.58081030845642,
-1.76459228992462,
-1.65098106861115,
-1.96331787109375,
-1.73259103298187,
-1.91794991493225,
-1.76102685928345,
-2.09321665763855,
-2.06416344642639,
-2.07215213775635,
-2.65714764595032,
-2.03192353248596,
-3.43564867973328,
-2.08765602111816,
-3.38544273376465,
-2.30686426162720,
-3.98799681663513,
-2.74154710769653,
-4.71619939804077,
-3.56363129615784,
-7.01465988159180,
-4.00696945190430,
28.4115219116211,
-6.42915916442871,
-29.0981693267822,
-10.7974786758423,
-1.84854602813721,
14.5533351898193,
12.0550689697266,
49.5718917846680,
33.9042358398438,
-14.8161058425903,
0.544351816177368,
0.0613934993743897,
-13.1170434951782,
-13.3595561981201,
-53.6686935424805,
1.41266775131226,
60.2425003051758,
-43.8310089111328,
-15.6436042785645,
6.10202884674072,
2.51057767868042,
5.12387990951538,
-14.1841926574707,
32.0684967041016,
-27.2989768981934,
24.0272960662842,
12.7188243865967,
-52.4527549743652,
-15.5973968505859,
-11.2145204544067,
-15.4370269775391,
-52.9664192199707,
41.2193031311035,
30.6836585998535,
-33.3864326477051,
39.4732780456543,
30.3626613616943,
-23.6771831512451,
-55.7813415527344,
-8.00340270996094,
-19.0007972717285,
-15.9499473571777,
35.3487434387207,
-45.1872024536133,
-31.8529720306397,
3.68921899795532,
-37.2195434570313,
-6.29013347625732,
16.9848823547363,
-26.2062358856201,
-1.74663782119751,
47.8320159912109,
18.7461204528809,
39.0357360839844,
47.0817260742188,
52.8130531311035,
30.9606361389160,
-29.7364768981934,
-19.2794361114502,
3.17606210708618,
12.3802356719971,
12.5912513732910,
62.1434669494629,
-15.9460315704346,
2.06738853454590,
51.2389335632324,
-62.9108047485352};
