shortreal out[65536] = '{0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
0.00000000000000,0.00000000000000,
-4.38911592937075e-06,4.38911592937075e-06,
0.000857615086715668,-0.000857615086715668,
-0.000130425411043689,1.70185739989392e-05,
-0.00294469785876572,0.00207644514739513,
0.000517314590979368,1.76012399606407e-05,
0.00888451281934977,-0.00483433110639453,
-0.00118979322724044,0.000103017773653846,
-0.0161311868578196,0.00776506913825870,
0.00295175332576036,2.91678588837385e-05,
0.0268595926463604,-0.0121033936738968,
-0.00542815960943699,-0.000286702532321215,
-0.0429344065487385,0.0182635802775621,
0.00903866346925497,0.00127281760796905,
0.0665498822927475,-0.0269927643239498,
-0.0118200145661831,-0.00539663946256042,
-0.102336540818214,0.0404747426509857,
-0.00669883098453283,0.0324266813695431,
0.102436713874340,-0.00545950885862112,
-0.0174739174544811,0.00462837843224406,
-0.116872042417526,0.0232486426830292,
0.0690425336360931,-0.0238357298076153,
0.144421368837357,-0.0498520135879517,
-0.297323763370514,0.0632123351097107,
-0.164491370320320,0.00982888787984848,
0.0569290779531002,0.0451888702809811,
0.410083800554276,-0.188530549407005,
-0.263645827770233,-0.163308382034302,
-0.392919868230820,0.294498562812805,
0.248755723237991,0.527588486671448,
0.539202868938446,-0.752772688865662,
-0.0791890770196915,-1.00755190849304,
-1.08938050270081,1.32884073257446,
-0.215780973434448,1.43418073654175,
1.63814187049866,-0.830794334411621,
0.647801756858826,-2.17863845825195,
-2.32431459426880,0.731393396854401,
-1.56910765171051,3.40720629692078,
3.05108094215393,-0.447411268949509,
3.71394872665405,-5.43856191635132,
-5.30884361267090,0.408017694950104,
-18.5073852539063,13.5823020935059,
-26.0687789916992,17.8305664062500,
-28.1438484191895,5.64882326126099,
-27.3125762939453,-3.57323980331421,
-20.3192501068115,9.07210254669190,
-3.06076955795288,28.3982944488525,
16.2501296997070,21.1651439666748,
21.8685855865479,-17.6394557952881,
8.75393104553223,-54.3817596435547,
-8.53807926177979,-55.1090316772461,
-11.0397119522095,-24.6573352813721,
1.02949464321136,4.37941741943359,
13.3652048110962,13.7510213851929,
13.9070215225220,3.96203231811523,
4.06555795669556,-19.4358692169189,
-4.13289737701416,-50.0434646606445,
2.87850165367126,-70.5329132080078,
27.5136985778809,-61.6138153076172,
47.3335075378418,-26.0172405242920,
40.0484199523926,2.96577715873718,
10.2771854400635,2.14516091346741,
-9.71932601928711,-15.2516822814941,
1.37613129615784,-14.6399679183960,
21.4920043945313,10.9131145477295,
15.6205263137817,32.8808593750000,
-15.7349863052368,21.8783817291260,
-35.0897102355957,-19.6480388641357,
-24.3956718444824,-51.8982734680176,
-6.97463178634644,-48.0531120300293,
-8.70646953582764,-18.2234382629395,
-12.2946414947510,3.50951695442200,
12.9963006973267,-2.89965510368347,
57.2841720581055,-22.2843322753906,
77.2303085327148,-24.6693058013916,
50.2490196228027,0.0566104650497437,
2.92156696319580,33.6583976745606,
-23.9154262542725,47.3199920654297,
-20.0616226196289,46.7733306884766,
-5.97481489181519,49.2110786437988,
2.03339838981628,50.7554435729981,
2.69306135177612,30.5889549255371,
-0.108316153287888,-13.7981605529785,
1.29324328899384,-46.2840957641602,
18.7352943420410,-36.4782638549805,
47.7942390441895,-4.14428710937500,
53.8056297302246,7.31033372879028,
15.2749395370483,-2.31932544708252,
-36.8956527709961,4.34524011611939,
-47.5175819396973,29.9348716735840,
-12.7465744018555,27.3365516662598,
12.6147241592407,-25.0556068420410,
-8.91567230224609,-74.2345199584961,
-42.5316429138184,-51.9048118591309,
-26.5903263092041,19.5662117004395,
27.5510616302490,51.9542617797852,
53.4687347412109,9.22649192810059,
28.7906131744385,-52.0507659912109,
-3.69163370132446,-62.5675773620606,
-4.66626405715942,-34.5553359985352,
4.20142698287964,-20.3649253845215,
-6.33035755157471,-27.3562221527100,
-20.2456588745117,-11.4876937866211,
-8.33281803131104,35.9198532104492,
9.35693740844727,68.7326660156250,
-5.61313056945801,45.9990768432617,
-44.1722297668457,-12.0187349319458,
-48.9561843872070,-54.1802940368652,
-2.50499916076660,-59.5849685668945,
37.1852455139160,-42.8602180480957,
18.5480480194092,-26.3473911285400,
-27.9413852691650,-18.9945125579834,
-37.1573448181152,-18.3413562774658,
3.89629125595093,-21.1473903656006,
48.9551849365234,-19.7709445953369,
61.2755432128906,-5.79500436782837,
47.0730171203613,5.51590156555176,
27.8348236083984,-8.94002342224121,
10.5473279953003,-39.5007019042969,
-0.0273989457637072,-58.4990653991699,
7.40352487564087,-50.6911430358887,
32.2767868041992,-28.8785610198975,
48.4044609069824,-8.44538593292236,
34.6210441589356,8.60961151123047,
13.4867267608643,24.7781238555908,
16.8414020538330,31.9543399810791,
36.2639312744141,24.0462989807129,
35.3924751281738,15.9877138137817,
1.10429441928864,18.1870975494385,
-35.2256278991699,16.3131008148193,
-37.8775978088379,-12.1578168869019,
-7.13160467147827,-47.6587066650391,
22.7822074890137,-45.7200775146484,
26.9132480621338,2.92930936813355,
9.40071964263916,51.0101623535156,
-14.7207746505737,54.7210426330566,
-27.1417884826660,22.8161201477051,
-11.9297904968262,-4.77601051330566,
30.1665706634522,-15.3083324432373,
68.0091018676758,-20.0640735626221,
68.0992126464844,-19.4645061492920,
30.9273719787598,-1.86707949638367,
-12.3457040786743,22.0311546325684,
-31.5797119140625,18.0947341918945,
-31.8735599517822,-19.3171215057373,
-29.6625957489014,-43.1945037841797,
-26.9857959747314,-18.6163043975830,
-16.3895149230957,27.7248992919922,
-2.98618698120117,40.7750892639160,
-3.13201212882996,14.7924823760986,
-7.88606548309326,-9.57822418212891,
5.95898056030273,-2.50069618225098,
33.5983734130859,23.8106460571289,
37.3028793334961,41.4497756958008,
-4.82509994506836,42.6442375183106,
-55.0846748352051,33.4928550720215,
-57.6059913635254,9.79997539520264,
-6.49112510681152,-19.7549571990967,
46.0440597534180,-29.1352500915527,
52.9615516662598,-6.98758172988892,
23.3557434082031,18.7935123443604,
-11.7792081832886,21.0396003723145,
-40.8622283935547,13.4913539886475,
-66.6282501220703,21.1762237548828,
-77.6283721923828,26.2149868011475,
-55.9571075439453,-4.23179435729981,
-13.6485261917114,-55.9317855834961,
14.1716871261597,-69.4300155639648,
8.73586559295654,-19.5681648254395,
-9.53743839263916,34.8970184326172,
-18.7843208312988,29.2749195098877,
-25.4863910675049,-17.6775512695313,
-42.6562919616699,-38.4082832336426,
-59.3494606018066,-17.2154083251953,
-45.7973480224609,1.21346795558929,
-0.205030083656311,-8.48309516906738,
42.1709403991699,-21.9156017303467,
53.9113655090332,-17.3996562957764,
40.7770347595215,-11.5123949050903,
24.4410972595215,-23.9305152893066,
11.4643392562866,-33.9880142211914,
-4.19113779067993,-16.4085559844971,
-20.5017833709717,9.69088554382324,
-21.9217262268066,7.05931949615479,
1.00590634346008,-19.0483608245850,
28.7771987915039,-23.9460945129395,
34.2491950988770,3.18482971191406,
10.9558706283569,20.7789306640625,
-20.4599800109863,8.69445323944092,
-29.1962852478027,-1.99883651733398,
-3.00394177436829,20.2738456726074,
31.1015586853027,49.9884757995606,
29.4189205169678,43.1768264770508,
-11.4587583541870,-2.16996383666992,
-44.1469268798828,-44.0053939819336,
-20.7753486633301,-50.5594062805176,
47.2187042236328,-36.5870666503906,
92.9870529174805,-20.8913040161133,
77.8048019409180,-5.04611730575562,
32.6939392089844,6.95841598510742,
10.6222858428955,-5.17940568923950,
16.9489459991455,-39.2432556152344,
14.1535377502441,-55.1126899719238,
-9.41647148132324,-25.0282154083252,
-19.7329063415527,25.4618053436279,
1.11973285675049,53.9027900695801,
26.7054653167725,54.3557052612305,
18.1411037445068,50.8901786804199,
-16.9510936737061,48.1896972656250,
-40.4639053344727,18.3057422637939,
-33.2517242431641,-38.3367843627930,
-11.2994003295898,-72.5606460571289,
7.15167856216431,-51.7928733825684,
14.3057546615601,-11.0955476760864,
9.80239582061768,3.57282781600952,
-5.23140096664429,-6.88323545455933,
-18.4049930572510,-2.53695821762085,
-2.56518840789795,18.3603630065918,
35.8605155944824,23.0923633575439,
56.0335922241211,4.26714420318604,
29.0087852478027,-2.46972060203552,
-21.4559669494629,20.5976715087891,
-51.8498992919922,33.8353347778320,
-52.1152725219727,-0.810570240020752,
-40.7262382507324,-52.2777328491211,
-35.9006271362305,-56.4195404052734,
-36.9305152893066,-10.6171598434448,
-36.1817779541016,25.1636028289795,
-36.2265625000000,5.99644088745117,
-33.9795341491699,-39.4470024108887,
-18.8519153594971,-65.1496810913086,
7.48417711257935,-63.7376976013184,
23.6309871673584,-58.9323081970215,
18.0784645080566,-51.2300910949707,
1.44241058826447,-22.4642581939697,
-19.4191455841064,17.6930294036865,
-45.5572357177734,26.2119960784912,
-62.3404884338379,-13.3392810821533,
-35.5853805541992,-55.4147796630859,
31.0128822326660,-45.9538421630859,
79.2675781250000,4.62320423126221,
55.8786659240723,34.1914100646973,
-12.1378250122070,11.2575073242188,
-40.6799545288086,-32.6628417968750,
-4.35183382034302,-47.1170845031738,
29.0308322906494,-24.3400554656982,
3.00010824203491,-1.00057470798492,
-46.5107116699219,-5.33539628982544,
-43.9417381286621,-22.6494960784912,
14.5774707794189,-27.9222831726074,
57.0981254577637,-13.6681327819824,
45.2847442626953,-0.564868032932282,
15.0569162368774,-4.82756233215332,
13.4653196334839,-25.4282684326172,
30.9633502960205,-43.0845642089844,
26.8818950653076,-39.4383430480957,
2.12143707275391,-21.8590183258057,
-10.1298036575317,-11.3917675018311,
1.17571198940277,-16.4385452270508,
7.50333023071289,-27.7668170928955,
-12.1914529800415,-30.2099323272705,
-35.7882575988770,-26.3712539672852,
-33.7778816223145,-26.6884822845459,
-4.17641735076904,-29.9942550659180,
30.2465991973877,-23.2654914855957,
51.2579879760742,-8.61830902099609,
52.1892547607422,-7.23266315460205,
36.4940261840820,-19.9264907836914,
9.43214797973633,-20.0912170410156,
-16.8643836975098,9.47378349304199,
-29.7300739288330,42.6430435180664,
-33.8567657470703,38.4569435119629,
-39.7887229919434,-2.94017982482910,
-44.5572853088379,-34.2966995239258,
-27.9390144348145,-25.0168209075928,
9.87220954895020,9.61887645721436,
37.8430976867676,34.2591018676758,
21.6681308746338,40.4452819824219,
-25.9141616821289,39.7287826538086,
-61.0189704895020,31.0130443572998,
-53.5990867614746,3.83141183853149,
-22.7159519195557,-31.5245914459229,
-9.36859321594238,-45.0982322692871,
-25.3189525604248,-23.8271121978760,
-42.3138542175293,10.6881971359253,
-30.8088417053223,24.0554733276367,
-0.636928319931030,9.94328975677490,
23.2393016815186,-13.3863048553467,
27.5704765319824,-26.0020885467529,
25.5264854431152,-19.1103057861328,
33.1331443786621,3.15988945960999,
38.2472305297852,31.0171813964844,
15.1840343475342,44.2909126281738,
-41.1996459960938,24.5319957733154,
-89.3054122924805,-15.6574621200562,
-83.8349990844727,-38.5932083129883,
-33.2427787780762,-22.8453159332275,
5.39091539382935,12.8726463317871,
-7.63584518432617,24.4505500793457,
-44.0378646850586,-1.54310333728790,
-37.8247299194336,-36.2280769348145,
23.1665477752686,-43.4158363342285,
78.1962585449219,-20.5252914428711,
77.0092163085938,5.49344396591187,
37.1911239624023,17.4205551147461,
3.62185716629028,18.4340152740479,
-11.6778182983398,18.1659259796143,
-26.3371524810791,19.8872394561768,
-35.4469184875488,25.5581760406494,
-16.8134174346924,32.4775238037109,
21.7851085662842,34.5393333435059,
31.9171619415283,18.4581336975098,
-2.75431537628174,-10.5986862182617,
-27.8525905609131,-31.7279548645020,
-3.10062313079834,-27.9604606628418,
39.3936691284180,-3.79732632637024,
34.6541595458984,21.6534175872803,
-11.7183456420898,35.5174713134766,
-28.3652000427246,36.7869567871094,
13.8303871154785,23.7964706420898,
56.5894660949707,5.73681879043579,
42.4757499694824,3.21064257621765,
-5.82997941970825,29.6584033966064,
-22.6990470886230,63.9391403198242,
-0.951124429702759,67.1399917602539,
7.66995191574097,29.7003536224365,
-16.2471733093262,-21.7739944458008,
-29.4828796386719,-49.3305130004883,
7.44158172607422,-42.0151138305664,
59.1254577636719,-17.9988403320313,
65.2838973999023,2.24506354331970,
26.6255302429199,4.27449274063110,
-5.10177612304688,-16.5269317626953,
0.598963499069214,-42.1703643798828,
21.0046024322510,-41.3320159912109,
17.5110416412354,-13.3227539062500,
-9.49456501007080,5.60841274261475,
-28.0136966705322,-15.4739151000977,
-18.8887557983398,-44.2179832458496,
0.315580487251282,-25.0999946594238,
4.86654615402222,40.1184349060059,
-16.1218948364258,74.2822570800781,
-47.3208770751953,29.8175659179688,
-58.1527862548828,-44.9139595031738,
-34.4165344238281,-58.9867553710938,
0.847067832946777,1.66537845134735,
6.95672416687012,56.3077850341797,
-18.4853324890137,40.6406822204590,
-36.5845680236816,-16.8451614379883,
-12.6403636932373,-38.5915260314941,
37.9157867431641,-2.52029752731323,
64.4161987304688,43.2497253417969,
48.0230751037598,50.8277702331543,
21.3283214569092,31.1080741882324,
17.3854045867920,26.8817405700684,
28.3550968170166,51.5184745788574,
27.7301578521729,68.9201889038086,
12.2689170837402,44.1647262573242,
-0.724178314208984,-9.49781703948975,
-3.67469549179077,-45.1082572937012,
-4.79153394699097,-39.4769172668457,
-6.82104253768921,-10.7644376754761,
8.17210483551025,4.21495819091797,
41.7761917114258,-8.05541038513184,
68.3775711059570,-15.8395385742188,
60.4067764282227,4.68593883514404,
24.4227409362793,34.8541183471680,
-5.44692516326904,41.8500175476074,
-11.0399675369263,21.3592758178711,
-4.57498502731323,7.47426939010620,
-0.718230307102203,21.6823577880859,
4.94607162475586,42.9799957275391,
19.8542156219482,41.1124496459961,
31.3375492095947,19.6625366210938,
20.1040763854980,13.2069549560547,
-12.2101106643677,22.6603183746338,
-38.3305282592773,12.2212247848511,
-39.5497245788574,-35.1758804321289,
-21.2517242431641,-80.8213958740234,
-2.56421756744385,-72.6467590332031,
6.18266820907593,-16.8599720001221,
6.95671224594116,28.8317871093750,
-3.10253095626831,23.0210800170898,
-24.3964843750000,-16.7582225799561,
-37.8212814331055,-50.0165252685547,
-27.6593036651611,-56.2389564514160,
6.23097753524780,-37.3311424255371,
37.1863250732422,-1.14141082763672,
37.4840888977051,40.4815788269043,
8.23232841491699,60.3647384643555,
-16.1430625915527,37.1983032226563,
-4.33002758026123,-7.52104568481445,
34.7118225097656,-27.9728870391846,
59.6390342712402,-6.04049062728882,
34.6977767944336,23.8713092803955,
-21.8243446350098,18.7417697906494,
-48.0555000305176,-19.1150341033936,
-13.0191450119019,-46.4575614929199,
39.4841308593750,-33.4633712768555,
39.6144180297852,1.55412948131561,
-17.7243175506592,24.4130783081055,
-65.2475280761719,24.0965709686279,
-51.2727012634277,12.0861196517944,
-8.75729084014893,-1.18226838111877,
-0.128374218940735,-9.43252658843994,
-32.4193954467773,-10.7910451889038,
-49.2191085815430,0.301748573780060,
-13.6667699813843,10.1586036682129,
39.1824264526367,5.65817832946777,
57.2506713867188,-9.99324893951416,
37.4747276306152,-11.1390018463135,
13.8926410675049,21.1802253723145,
4.82217073440552,60.8323974609375,
-2.05029296875000,63.5091552734375,
-12.7806568145752,17.7920379638672,
-19.2917842864990,-40.2260322570801,
-14.6931095123291,-66.8443832397461,
-5.82478713989258,-49.6007041931152,
5.91636753082275,-12.9296302795410,
23.4635314941406,13.4896125793457,
37.3348999023438,25.0179824829102,
28.4116821289063,36.6392250061035,
-5.02455139160156,57.1361656188965,
-28.3467407226563,70.9660110473633,
-13.2224779129028,52.8207283020020,
12.2013130187988,3.02936744689941,
5.54605627059937,-44.3632583618164,
-24.9425048828125,-56.7881431579590,
-25.9288845062256,-37.6904296875000,
31.4715290069580,-20.4838867187500,
93.4933319091797,-17.3477611541748,
90.8036651611328,-5.14823150634766,
21.3230934143066,21.0861053466797,
-45.7055358886719,36.7620201110840,
-56.9300918579102,21.1693572998047,
-26.4266662597656,-7.72145700454712,
1.06473898887634,-13.2195167541504,
7.84912443161011,5.18935918807983,
4.38917160034180,15.1807994842529,
-6.95699977874756,6.35090160369873,
-30.7264442443848,-0.865526914596558,
-54.8461265563965,2.96133303642273,
-51.0626411437988,-5.09713983535767,
-9.22829246520996,-36.8587760925293,
45.3533363342285,-55.1532287597656,
75.7751693725586,-23.5985984802246,
71.2973709106445,33.4152793884277,
54.2877502441406,58.3327140808106,
43.5073928833008,32.0933723449707,
35.9550514221191,-3.98493719100952,
26.7187194824219,-17.8959255218506,
8.53926467895508,-25.5022525787354,
-10.2172117233276,-49.8315277099609,
-11.3046140670776,-75.5158004760742,
12.0950727462769,-67.7344970703125,
44.7675209045410,-30.5279521942139,
59.6201858520508,-5.87583875656128,
44.9774856567383,-9.43039417266846,
21.5802268981934,-10.7510166168213,
15.5474796295166,13.6960191726685,
17.9665412902832,46.1947746276856,
-0.0878022387623787,49.8167114257813,
-37.6159667968750,16.6090011596680,
-52.3206062316895,-25.4631309509277,
-16.4084663391113,-45.0532608032227,
43.7641143798828,-35.2421379089356,
71.8169555664063,-12.3368225097656,
55.3202133178711,0.314659655094147,
28.0526084899902,-10.6774358749390,
20.0197277069092,-36.8866806030273,
17.8053684234619,-45.3546905517578,
-2.59304976463318,-17.2169208526611,
-32.1393089294434,26.8023910522461,
-36.6536865234375,35.1138610839844,
-5.76242876052856,-2.82280611991882,
33.2730369567871,-46.0771598815918,
40.0139884948731,-44.1786308288574,
12.1019134521484,0.713084697723389,
-22.1552200317383,39.7915420532227,
-34.3067588806152,34.4568595886231,
-17.2237205505371,-1.64802157878876,
9.92430686950684,-34.5344352722168,
20.3383865356445,-48.3815078735352,
11.4288768768311,-46.4577903747559,
1.17621839046478,-34.6535186767578,
-2.14067959785461,-11.9638795852661,
-1.85554242134094,14.3753252029419,
-9.09121990203857,31.5180530548096,
-17.1117725372314,35.6948051452637,
-15.0772037506104,39.9337615966797,
-9.28640747070313,48.3230628967285,
-22.4465637207031,45.8564796447754,
-51.5091552734375,23.3216667175293,
-55.2515754699707,-7.21745061874390,
-10.8298349380493,-15.1723022460938,
43.4935569763184,7.03552150726318,
49.7091331481934,28.0139274597168,
2.35833859443665,24.6748371124268,
-34.4905967712402,3.52762269973755,
-14.5415534973145,-11.1831521987915,
34.0331306457520,-10.2086706161499,
54.5741691589356,-9.91999149322510,
34.8940773010254,-16.7060871124268,
14.4889898300171,-18.2909202575684,
18.8832836151123,-0.0956823825836182,
23.2461471557617,25.6200771331787,
2.51489686965942,28.1710910797119,
-25.8667278289795,-3.86313748359680,
-26.6852512359619,-51.1551513671875,
-1.14610016345978,-74.2970504760742,
19.5289268493652,-51.5282859802246,
10.6526393890381,3.55994915962219,
-18.8446159362793,46.7855873107910,
-42.9492454528809,46.3240394592285,
-39.1508102416992,11.4834556579590,
-6.85609292984009,-19.7605457305908,
32.4875488281250,-21.9916095733643,
42.5794982910156,-10.6821470260620,
6.94010925292969,-12.0435009002686,
-41.7206039428711,-20.8321571350098,
-51.2158393859863,-7.11249542236328,
-14.7567415237427,32.8707351684570,
20.0025844573975,59.7141952514648,
19.4737606048584,45.0470466613770,
9.60366058349609,9.36259937286377,
24.6890773773193,-6.15336275100708,
48.5187568664551,5.71567058563232,
37.1658782958984,10.4509115219116,
-13.5897922515869,-10.8868265151978,
-50.3379478454590,-31.9608039855957,
-32.5783462524414,-24.4381656646729,
13.6331081390381,1.80119442939758,
37.6210975646973,16.8663349151611,
26.6825962066650,14.9989690780640,
-2.49468088150024,17.1180191040039,
-36.2974395751953,23.7122879028320,
-63.1878738403320,11.2988262176514,
-60.7946968078613,-23.7600135803223,
-18.5510139465332,-48.5128059387207,
25.6872043609619,-30.2677669525147,
25.1806888580322,16.5278663635254,
-10.9030199050903,45.1120491027832,
-22.5452232360840,28.5422515869141,
15.1252765655518,-12.6123600006104,
49.3066825866699,-42.2697830200195,
27.1856327056885,-42.7372589111328,
-25.2039146423340,-22.1135730743408,
-31.4729328155518,0.617059469223023,
19.1332244873047,6.74316978454590,
53.8703804016113,-9.66009330749512,
24.8577785491943,-24.8997745513916,
-33.6073036193848,-11.2852106094360,
-55.8306083679199,28.7469749450684,
-27.7176589965820,57.3733367919922,
5.93653964996338,44.2265129089356,
7.94404935836792,1.72164702415466,
-15.0881576538086,-27.7161407470703,
-32.5739784240723,-18.8614959716797,
-29.4551315307617,10.2247819900513,
-11.4953289031982,25.7093524932861,
2.16378641128540,15.7333297729492,
-7.82320499420166,-9.75148391723633,
-38.8384132385254,-27.7725620269775,
-51.9986648559570,-19.4505138397217,
-15.7948160171509,10.4499940872192,
38.0188560485840,34.9922180175781,
44.6334381103516,29.8631515502930,
-7.36408901214600,2.63073301315308,
-50.6690101623535,-13.4416666030884,
-26.3108596801758,-2.02796506881714,
36.5074768066406,14.7849102020264,
55.4450988769531,10.9341802597046,
11.8326730728149,-1.45292687416077,
-34.7305259704590,9.06094837188721,
-38.8524169921875,37.3431587219238,
-28.1945152282715,41.1981887817383,
-40.4917068481445,2.79991555213928,
-59.6004486083984,-37.5813026428223,
-41.7796516418457,-34.0683784484863,
2.78153228759766,0.528551101684570,
23.6602725982666,13.0562734603882,
0.678470134735107,-15.4773960113525,
-27.2880096435547,-40.1452102661133,
-24.0229492187500,-21.7400398254395,
-5.40056467056274,20.5393142700195,
-3.99309372901917,33.4671134948731,
-18.8314933776855,-2.86160469055176,
-23.5450553894043,-48.3966903686523,
-13.4071683883667,-55.0652198791504,
-9.60302829742432,-19.1083793640137,
-18.0270977020264,23.5884513854980,
-28.1188411712647,33.8299217224121,
-32.0325508117676,3.84585165977478,
-29.7207984924316,-43.5942268371582,
-17.2887554168701,-69.8140716552734,
14.5482845306396,-58.4330291748047,
48.7041549682617,-20.1350116729736,
50.5904502868652,22.4689788818359,
6.18664264678955,49.9307708740234,
-45.3101959228516,52.0163650512695,
-50.4160156250000,30.0947761535645,
-10.3080720901489,-3.87466955184937,
27.3944435119629,-28.6123847961426,
32.6929702758789,-21.9012393951416,
21.8820934295654,4.56467485427856,
18.5658111572266,19.8472957611084,
23.1397418975830,17.7763042449951,
22.1777362823486,19.9963016510010,
11.2829608917236,41.4840927124023,
-3.11468100547791,59.3691139221191,
-17.3447341918945,45.0217895507813,
-31.0420131683350,10.1984214782715,
-33.0554275512695,-5.48938322067261,
-18.4424781799316,3.75257730484009,
-5.57493305206299,3.27500748634338,
-15.4769792556763,-26.6677532196045,
-37.2008666992188,-50.3235702514648,
-37.9149551391602,-22.4990959167480,
-16.0560913085938,34.5991020202637,
-7.83947610855103,58.4433364868164,
-22.7097549438477,25.6694030761719,
-28.3769798278809,-16.7100925445557,
3.06738042831421,-21.4140090942383,
41.7672233581543,-3.66485691070557,
39.7481117248535,-5.45623922348023,
2.36249828338623,-31.4972438812256,
-17.2333793640137,-39.6483497619629,
1.32460093498230,-12.3614416122437,
15.7690124511719,18.1609897613525,
-5.60425996780396,13.7686815261841,
-36.0994415283203,-17.2428493499756,
-33.1069946289063,-40.6886482238770,
-3.92829751968384,-43.4720916748047,
16.0515804290772,-38.1265945434570,
19.7465934753418,-33.9446830749512,
28.6594791412354,-23.5236606597900,
45.2473945617676,-7.78796148300171,
43.6877136230469,2.29411745071411,
18.0179805755615,7.21397113800049,
-3.08532547950745,19.6875591278076,
-3.10310053825378,42.9116096496582,
-4.24569749832153,54.5619773864746,
-26.2954139709473,31.9444923400879,
-47.1972389221191,-9.70279693603516,
-35.9508361816406,-29.9044437408447,
-8.26738452911377,-14.2188844680786,
-4.43582630157471,13.8984584808350,
-28.7151718139648,24.3982639312744,
-39.0069160461426,17.3163528442383,
-13.9967479705811,15.6374740600586,
13.1646575927734,27.4689273834229,
-2.99349164962769,34.4472084045410,
-47.4961318969727,15.5745286941528,
-63.2604866027832,-21.7195777893066,
-26.4472370147705,-39.9442062377930,
22.9775924682617,-19.5751495361328,
28.1754093170166,20.2058963775635,
-8.06362342834473,42.8687973022461,
-41.0385665893555,33.4137573242188,
-40.8132362365723,9.63838577270508,
-26.0566902160645,-6.89800548553467,
-25.5662422180176,-13.8632688522339,
-37.1620559692383,-18.4821605682373,
-38.9956283569336,-12.0994024276733,
-29.0560951232910,8.84037399291992,
-23.8641681671143,18.4857368469238,
-22.7582492828369,-12.4126033782959,
-3.80297827720642,-62.4091453552246,
34.6120300292969,-71.0212326049805,
54.3553848266602,-16.5637931823730,
26.1797351837158,46.2214050292969,
-28.0652999877930,49.8834457397461,
-60.5979614257813,0.851349830627441,
-53.0197525024414,-35.5223999023438,
-33.1884269714356,-33.5669898986816,
-20.2866134643555,-30.3128318786621,
-5.83794879913330,-52.5906219482422,
18.4152412414551,-66.4069824218750,
36.6884002685547,-36.4750137329102,
29.5936203002930,6.62232875823975,
12.7623701095581,8.53896331787109,
10.2147893905640,-24.3686103820801,
22.8576908111572,-30.8395843505859,
23.9454383850098,12.2721843719482,
-0.855430364608765,51.2745437622070,
-33.5049438476563,37.7151184082031,
-44.8121986389160,0.588465690612793,
-29.3954925537109,-3.43382549285889,
-5.32181167602539,28.2505302429199,
13.3827838897705,40.4822463989258,
25.5121841430664,6.91979503631592,
35.6918411254883,-29.6581897735596,
44.0388488769531,-30.3138771057129,
34.0125617980957,-9.86004447937012,
-3.67859649658203,-3.42338466644287,
-49.8111000061035,-11.9898796081543,
-62.5250892639160,-7.71102476119995,
-28.0248622894287,17.1008358001709,
20.5744094848633,35.2131652832031,
32.3687705993652,24.9108371734619,
2.54011726379395,-0.469221591949463,
-30.7582550048828,-16.0505447387695,
-36.0804443359375,-14.7475137710571,
-21.8893089294434,-6.64293003082275,
-13.0571393966675,5.45279502868652,
-7.47619724273682,9.24309444427490,
7.06236600875855,-5.64834403991699,
25.0684223175049,-33.9081535339356,
27.9752864837647,-44.1189613342285,
17.1323051452637,-15.8075828552246,
12.8846435546875,33.6081314086914,
21.5777606964111,56.6804618835449,
30.8100643157959,38.5253105163574,
33.9018516540527,7.79669189453125,
40.2116050720215,-0.623613178730011,
47.8217582702637,13.2779130935669,
32.0630683898926,29.8353939056397,
-17.6307792663574,40.0335197448731,
-68.7693557739258,41.1882209777832,
-75.5570602416992,23.6190509796143,
-37.2833213806152,-21.2346897125244,
0.330258965492249,-71.0152511596680,
6.32871246337891,-84.0707015991211,
-3.92595028877258,-50.8393211364746,
-1.65581631660461,-11.2482576370239,
8.38261985778809,-11.0200138092041,
-1.51747107505798,-47.4856719970703,
-27.1437873840332,-74.6070175170898,
-35.4289741516113,-62.2653503417969,
-3.45933771133423,-29.3199062347412,
46.2225990295410,-10.7309255599976,
64.2983779907227,-17.3820285797119,
35.1552047729492,-23.5747203826904,
-6.58615541458130,-4.37498188018799,
-17.3268489837647,30.1399269104004,
4.00029706954956,47.2488632202148,
23.9831848144531,29.6531085968018,
19.4503231048584,-7.02432155609131,
1.77624595165253,-28.4010696411133,
0.394834786653519,-17.7010059356689,
13.2681121826172,7.40170478820801,
4.44045639038086,18.7761783599854,
-39.7613983154297,-1.76846683025360,
-78.0943298339844,-34.9551353454590,
-62.4979171752930,-46.6079940795898,
-2.19208717346191,-23.1090145111084,
37.8353385925293,12.7275753021240,
16.0493240356445,26.7376251220703,
-32.0909919738770,7.04057073593140,
-37.6356658935547,-24.9289398193359,
1.18101429939270,-39.3296623229981,
29.1874523162842,-31.0727329254150,
18.5062713623047,-16.0179080963135,
5.83263063430786,-6.73748445510864,
27.7297344207764,-5.97135305404663,
55.0130996704102,-4.40539264678955,
35.9230079650879,6.45900058746338,
-16.9693679809570,23.4834194183350,
-32.9625511169434,32.8661079406738,
11.2170295715332,19.8743438720703,
55.7486381530762,-6.40053653717041,
41.5184402465820,-14.3378419876099,
-1.42744064331055,8.23735427856445,
-4.14077377319336,33.9920845031738,
40.1349525451660,26.5239162445068,
66.1348648071289,-8.81558418273926,
35.1551742553711,-26.0430431365967,
-11.7531585693359,-1.69335293769836,
-22.9558944702148,31.3074073791504,
-6.69520187377930,32.6191406250000,
-3.97650742530823,2.70526862144470,
-29.5685672760010,-24.2103691101074,
-53.3510322570801,-30.6512088775635,
-46.8685684204102,-23.0860824584961,
-14.9950199127197,-10.5876770019531,
18.8020744323730,1.56959128379822,
40.4706497192383,5.14032888412476,
41.2018928527832,-13.5389118194580,
17.2002048492432,-40.4114761352539,
-13.8796854019165,-42.6516036987305,
-28.6059265136719,-13.4842138290405,
-28.2612991333008,12.3617897033691,
-24.9918422698975,2.99394893646240,
-13.3099174499512,-19.8390617370605,
19.0241127014160,-20.9327850341797,
56.9529228210449,-5.46205902099609,
58.8578224182129,-7.07733106613159,
11.3935852050781,-27.8185195922852,
-38.3283576965332,-28.9469738006592,
-35.7468948364258,7.87103176116943,
3.04919528961182,41.4633407592773,
16.7252082824707,23.1991729736328,
-3.54317188262939,-27.8638725280762,
-8.88204002380371,-52.7052116394043,
23.1353778839111,-29.3886966705322,
49.9141502380371,4.19014167785645,
25.8216609954834,12.5606298446655,
-20.6698246002197,14.3116502761841,
-32.6410865783691,37.6806068420410,
-11.3720855712891,64.5014495849609,
-4.61876821517944,59.0728187561035,
-22.4503536224365,15.3725385665894,
-19.1294879913330,-26.3484649658203,
26.5720157623291,-28.8949489593506,
65.8942337036133,-2.32617282867432,
45.7607612609863,11.7620859146118,
-4.91670846939087,-7.88216829299927,
-21.6479301452637,-38.6822853088379,
-0.313454151153564,-42.0633735656738,
6.63476657867432,-6.02944946289063,
-27.0219135284424,38.4921264648438,
-63.6328887939453,37.4625892639160,
-56.7266159057617,-21.4043350219727,
-15.3293676376343,-73.5657424926758,
20.1217594146729,-52.9314727783203,
29.9167118072510,28.0470104217529,
24.7223796844482,83.2334747314453,
8.77962303161621,62.3957023620606,
-15.9152832031250,9.61745643615723,
-26.0440425872803,-4.00394201278687,
-0.832300901412964,21.2148399353027,
38.3124160766602,27.7947502136230,
40.3224754333496,2.05416679382324,
2.95565414428711,-7.85556411743164,
-27.1001281738281,22.3335361480713,
-10.9797992706299,45.6392021179199,
27.7475128173828,21.1496810913086,
37.1675987243652,-21.2822170257568,
9.77084350585938,-18.5989875793457,
-15.0482902526855,30.4124393463135,
-15.3695926666260,65.4414978027344,
-12.0531454086304,56.9191932678223,
-20.5563755035400,33.7246589660645,
-27.3712234497070,26.4581642150879,
-16.5312175750732,23.8774356842041,
6.53903388977051,4.97411298751831,
32.6505317687988,-14.4878158569336,
58.2646255493164,-10.2655410766602,
77.8703918457031,5.88192224502564,
71.7455596923828,-1.13994479179382,
32.4040946960449,-28.7527885437012,
-9.41330623626709,-49.2092018127441,
-16.7344875335693,-50.9242744445801,
2.88730287551880,-51.2583084106445,
7.58145236968994,-57.0038604736328,
-14.7108154296875,-55.7440071105957,
-28.8459892272949,-40.1461677551270,
-15.4655342102051,-30.1504688262939,
-0.256216317415237,-39.7817420959473,
-8.53956317901611,-51.1520729064941,
-15.0176191329956,-33.7838020324707,
17.6175270080566,-0.124116897583008,
71.5307464599609,20.2221927642822,
89.7524566650391,24.7180900573730,
43.7599868774414,39.6409339904785,
-21.6851081848145,65.7816009521484,
-50.3263702392578,73.0266799926758,
-33.6477546691895,46.7665061950684,
-6.20357704162598,14.2245855331421,
9.09994983673096,10.9147405624390,
13.8100700378418,34.4378280639648,
11.9135894775391,49.8994789123535,
5.44932651519775,44.4320716857910,
-0.693093657493591,28.4114170074463,
-9.74921798706055,8.89800071716309,
-26.8358230590820,-21.4421653747559,
-45.0808753967285,-51.6881942749023,
-36.6975479125977,-53.6309089660645,
11.2233953475952,-25.3490619659424,
64.6989669799805,-2.67944097518921,
70.4014358520508,-10.1748809814453,
22.0067443847656,-25.2376594543457,
-21.0449047088623,-11.2350282669067,
-20.6396446228027,23.9169139862061,
-8.02218914031982,39.5896568298340,
-17.4658660888672,15.6499719619751,
-30.6448287963867,-14.6737270355225,
-6.95357561111450,-15.8519754409790,
38.0108146667481,6.42600297927856,
38.4258842468262,23.2157211303711,
-23.0514068603516,27.1843719482422,
-80.2653808593750,18.6518859863281,
-75.0821685791016,-3.56200957298279,
-34.2261962890625,-36.1551513671875,
-21.4121360778809,-55.1199417114258,
-30.8366222381592,-43.8097457885742,
-9.03116703033447,-19.5467548370361,
47.4974975585938,-7.17691802978516,
67.3772125244141,-7.23103857040405,
9.71710491180420,3.04651117324829,
-63.3335533142090,21.7313117980957,
-67.9162979125977,17.4868450164795,
-6.92122650146484,-12.6038217544556,
40.4061660766602,-21.5229206085205,
28.3359355926514,14.0513057708740,
-12.3211135864258,53.4621009826660,
-34.6233406066895,50.1084213256836,
-38.2606201171875,19.2115097045898,
-43.3454895019531,3.89115643501282,
-40.3939933776856,5.13010358810425,
-10.3069400787354,-12.2264289855957,
26.1515254974365,-43.4562072753906,
35.7130126953125,-36.7393074035645,
16.9478034973145,17.3343238830566,
3.27573752403259,55.6974716186523,
13.7336091995239,24.5751209259033,
30.8220844268799,-31.0348739624023,
30.5694923400879,-31.9374866485596,
12.1491422653198,16.7801322937012,
-6.42603683471680,44.9985771179199,
-19.2082233428955,22.6963806152344,
-24.3360481262207,-2.26930546760559,
-14.8564815521240,7.22478103637695,
1.12505578994751,26.9919185638428,
-2.01401162147522,18.8728103637695,
-30.2118225097656,-6.05358028411865,
-56.1622848510742,-8.28410339355469,
-48.5414657592773,9.57880401611328,
-21.5908279418945,14.5529041290283,
-8.68595027923584,5.93496513366699,
-16.6624870300293,13.4472789764404,
-18.0986328125000,33.4972648620606,
-0.0371239781379700,23.0846157073975,
12.9402360916138,-30.2383365631104,
1.76948428153992,-73.8888244628906,
-9.48955249786377,-68.0441436767578,
2.37730550765991,-39.5771331787109,
18.0218887329102,-36.6462326049805,
7.06239366531372,-58.2741203308106,
-21.5439929962158,-55.7510261535645,
-33.6889839172363,-13.6398353576660,
-26.6822738647461,21.0626640319824,
-25.6776084899902,12.3117895126343,
-30.4237136840820,-16.3478183746338,
-12.7854728698730,-25.9193000793457,
31.5287303924561,-19.0171241760254,
59.4966506958008,-22.9430141448975,
38.6786651611328,-37.6146774291992,
4.13957595825195,-43.1042022705078,
5.98659706115723,-33.4419937133789,
34.3751564025879,-20.2918071746826,
36.5904273986816,-4.63805150985718,
1.56263625621796,20.8274688720703,
-21.8939456939697,44.5315437316895,
-8.97496414184570,34.5815010070801,
10.7900638580322,-11.9335079193115,
4.15128707885742,-54.9388961791992,
-3.39201164245605,-56.6422500610352,
26.2481613159180,-30.2530555725098,
78.2922363281250,-4.48362731933594,
88.9596252441406,16.1406269073486,
39.5426521301270,38.3363647460938,
-17.7231864929199,46.1391258239746,
-26.8780746459961,23.8978309631348,
3.87738013267517,-10.4460725784302,
23.5502986907959,-18.3622112274170,
14.1006708145142,4.44574594497681,
-9.98641872406006,20.1881275177002,
-31.2808399200439,2.96965885162354,
-47.3535881042481,-19.4501266479492,
-60.2302932739258,-15.5551834106445,
-66.5097122192383,1.32806515693665,
-63.8830184936523,-1.57292830944061,
-59.5366973876953,-15.3449287414551,
-55.8621177673340,-15.1511716842651,
-46.1835212707520,-9.04748344421387,
-27.5509185791016,-22.3705215454102,
-10.3484039306641,-48.4584999084473,
5.24572849273682,-42.4026374816895,
32.8488349914551,4.97203111648560,
58.2587051391602,44.4876632690430,
50.0077438354492,36.6451797485352,
2.93808794021606,6.22987365722656,
-37.6129722595215,4.05478096008301,
-22.0970458984375,23.1613655090332,
29.7164955139160,17.6107006072998,
50.8130493164063,-13.5842552185059,
17.5515556335449,-16.5011863708496,
-18.2775459289551,27.8971309661865,
-15.4625110626221,69.4623947143555,
-2.49217438697815,58.3660202026367,
-28.5692062377930,8.34524726867676,
-75.8704605102539,-30.3651695251465,
-74.7966842651367,-43.0184478759766,
-10.0445880889893,-47.4579391479492,
58.1327438354492,-44.4509925842285,
70.5090942382813,-16.9533882141113,
44.6370811462402,28.3317127227783,
36.7636604309082,47.6255722045898,
57.4748802185059,22.5371570587158,
69.9865951538086,-10.0415229797363,
47.9630584716797,-18.3346138000488,
15.5414199829102,-14.3347215652466,
8.69315052032471,-22.8804168701172,
27.6956844329834,-35.2699966430664,
51.4656372070313,-24.9462966918945,
63.1036224365234,7.69302415847778,
53.1178016662598,36.4166526794434,
22.3306045532227,42.7434806823731,
-13.6035108566284,36.8399429321289,
-31.7200889587402,26.0279312133789,
-27.9692401885986,-1.50211429595947,
-15.8317461013794,-34.3270492553711,
-12.9319801330566,-40.2237167358398,
-21.3048171997070,-12.3416938781738,
-27.7731781005859,9.07066631317139,
-34.1788253784180,-7.04557418823242,
-41.1112899780273,-33.4478034973145,
-36.3969726562500,-25.6568222045898,
-2.79694867134094,10.6469507217407,
36.7893066406250,24.3008365631104,
46.2267074584961,0.725301504135132,
25.4483337402344,-15.9363403320313,
9.53204536437988,3.99938249588013,
15.5273132324219,23.0627956390381,
17.7673225402832,-9.44641113281250,
-3.46361660957336,-63.6365203857422,
-23.3048381805420,-67.7525253295898,
-4.71342992782593,-7.55021667480469,
34.5732536315918,45.2573318481445,
44.0809402465820,32.8110389709473,
22.3866310119629,-15.4626789093018,
16.7978801727295,-33.1781349182129,
42.6898765563965,-4.34230470657349,
52.3203506469727,24.2937450408936,
12.6591377258301,15.0446071624756,
-33.5229034423828,-18.2861137390137,
-20.5878524780273,-39.0940475463867,
35.3746337890625,-34.9191207885742,
59.9688072204590,-14.4791774749756,
26.2643394470215,12.7868862152100,
-7.53245353698731,35.1344490051270,
16.3658924102783,39.3956871032715,
67.3746871948242,30.9240608215332,
73.6817550659180,23.2289543151855,
22.7823867797852,18.7291946411133,
-24.6967258453369,9.66091918945313,
-20.3092327117920,-5.04632949829102,
17.2253570556641,-15.3736305236816,
42.4754219055176,-6.73361873626709,
39.2606964111328,10.6851692199707,
27.3053054809570,18.9937648773193,
25.7367115020752,20.6545028686523,
35.0799293518066,24.7775783538818,
43.2358016967773,21.4274635314941,
44.3774566650391,-1.50650000572205,
32.8325195312500,-21.9507141113281,
7.78198480606079,-7.74055290222168,
-20.0414752960205,36.3981132507324,
-31.1574974060059,59.7502059936523,
-20.4425029754639,34.5251350402832,
-5.08939170837402,1.83918845653534,
1.34702670574188,16.2145748138428,
-0.560872077941895,66.5222091674805,
-5.45971775054932,88.2457656860352,
-12.0475521087646,51.6596755981445,
-21.1696434020996,-0.675368010997772,
-22.9244022369385,-15.5462808609009,
-3.90871548652649,2.56861257553101,
26.1354789733887,15.8011646270752,
38.2662124633789,13.1318788528442,
12.7571277618408,17.6535263061523,
-29.2990875244141,38.6073036193848,
-49.0530853271484,49.0040626525879,
-25.6113414764404,29.6411705017090,
21.7393627166748,-3.62519836425781,
49.0307044982910,-19.3156719207764,
29.4920234680176,-9.78602027893066,
-21.4981517791748,0.998028635978699,
-58.0093765258789,-4.44162654876709,
-50.2073898315430,-16.0505752563477,
-11.9267101287842,-16.2761878967285,
13.2155809402466,-8.35906028747559,
5.08508396148682,-4.92691802978516,
-10.1106433868408,-19.0013256072998,
-4.71182680130005,-40.2992439270020,
14.9092006683350,-47.9440269470215,
15.5266456604004,-37.9147262573242,
-9.53879928588867,-25.8424358367920,
-22.7592773437500,-29.0226669311523,
3.65803194046021,-42.2811622619629,
48.1535797119141,-41.4632034301758,
63.7279815673828,-10.9225759506226,
35.7987403869629,30.7310867309570,
0.557502150535584,44.4768142700195,
-0.718612551689148,18.5355453491211,
29.6279850006104,-14.8285284042358,
51.3158569335938,-14.0048122406006,
29.8018932342529,23.6197853088379,
-23.5241489410400,52.4659576416016,
-66.4198455810547,37.6907691955566,
-63.2090148925781,-8.87759876251221,
-18.4738006591797,-43.6082229614258,
24.1407623291016,-43.7539100646973,
22.9238491058350,-27.0504837036133,
-14.8391819000244,-13.8564004898071,
-45.2540206909180,-0.825403928756714,
-42.0329055786133,24.4376106262207,
-23.3121051788330,50.3664855957031,
-17.9863834381104,50.7002487182617,
-19.9954948425293,16.4431114196777,
-6.83922719955444,-22.1378803253174,
23.3351840972900,-26.7085952758789,
34.9005699157715,7.13735151290894,
11.2669324874878,53.9152679443359,
-16.2362022399902,80.9200820922852,
-14.9327802658081,73.2975158691406,
4.14626979827881,39.7852516174316,
3.11527347564697,4.42216491699219,
-26.0380058288574,-6.23359012603760,
-46.7774467468262,13.3498497009277,
-35.1808700561523,40.2480926513672,
-7.21178054809570,46.1931457519531,
5.92783117294312,29.6268997192383,
-2.78379821777344,17.3831863403320,
-19.7209205627441,23.2839374542236,
-34.4456977844238,27.5148220062256,
-47.1500625610352,4.97365713119507,
-51.2343444824219,-32.9795875549316,
-38.8009147644043,-44.6011505126953,
-15.3594188690186,-14.9046707153320,
1.86004602909088,19.9484348297119,
7.29870939254761,18.0235939025879,
12.2554311752319,-15.7422733306885,
17.8152103424072,-34.6690368652344,
12.2896480560303,-12.3922986984253,
-12.6572027206421,30.0680694580078,
-38.5897865295410,50.1514663696289,
-41.4144134521484,31.6893157958984,
-15.3735294342041,-3.52412390708923,
14.5584716796875,-28.1555213928223,
23.1822090148926,-32.9965553283691,
12.6291942596436,-21.7425918579102,
-0.520758688449860,-4.94106769561768,
-2.41947817802429,11.0342044830322,
4.07197189331055,20.6917057037354,
5.11316204071045,18.7607383728027,
-7.06037807464600,3.39435887336731,
-28.4570007324219,-20.2652206420898,
-41.8281097412109,-37.2285232543945,
-41.2386970520020,-33.8872566223145,
-35.4076728820801,-11.5918951034546,
-40.2280883789063,6.74314498901367,
-50.9383544921875,-4.17605447769165,
-44.2233352661133,-37.4546318054199,
-7.38275384902954,-54.8067817687988,
43.8951911926270,-31.0425987243652,
75.1460266113281,18.1036472320557,
67.6292419433594,50.2352371215820,
33.5824470520020,44.9411048889160,
-0.883311271667481,26.6087131500244,
-17.9827308654785,23.4682769775391,
-18.8997650146484,30.3279418945313,
-11.5896797180176,22.1968421936035,
0.348040938377380,-2.06458926200867,
18.5178890228272,-16.0086479187012,
40.4151115417481,-5.72094345092773,
52.2689590454102,8.99064159393311,
36.2746887207031,4.93670225143433,
0.0850623846054077,-8.74186992645264,
-24.5132369995117,-5.98681497573853,
-13.1406116485596,9.35428333282471,
16.9286308288574,10.9461622238159,
32.8560295104981,-8.22699737548828,
20.2887630462647,-23.4091320037842,
1.11815261840820,-10.9070291519165,
-3.19982361793518,12.2999067306519,
-2.86523771286011,13.9280452728271,
-9.21314144134522,-2.78156328201294,
-15.1377372741699,-10.1278867721558,
-4.34926748275757,5.85308837890625,
11.8978643417358,23.3141059875488,
9.28419208526611,22.1425514221191,
-13.2272396087646,9.64553165435791,
-24.6692104339600,9.14690113067627,
-7.77476882934570,28.7254505157471,
13.7279052734375,49.4933242797852,
3.85751175880432,50.2555656433106,
-36.3877296447754,29.2408008575439,
-70.2069702148438,-0.0802018418908119,
-67.7107086181641,-18.9024658203125,
-35.0710105895996,-17.1573638916016,
0.548156619071960,0.391855508089066,
23.8469734191895,17.2352504730225,
29.1129341125488,22.8835716247559,
14.7834224700928,14.9228372573853,
-17.2797622680664,-0.882970154285431,
-52.7946166992188,-18.7083568572998,
-66.9162216186523,-25.5405750274658,
-49.9142990112305,-13.0230474472046,
-20.6580467224121,12.4817590713501,
-5.05419301986694,29.2796554565430,
-5.93179702758789,18.6076202392578,
-7.06660985946655,-9.42801666259766,
1.03614044189453,-29.2445526123047,
6.01875448226929,-28.1494064331055,
1.43041849136353,-14.6922330856323,
3.98413085937500,-8.41939353942871,
25.8241729736328,-13.8453035354614,
49.2761650085449,-28.1931991577148,
37.0000991821289,-43.9425048828125,
-6.01362991333008,-46.5401687622070,
-34.4255561828613,-21.6488456726074,
-23.3767890930176,21.9613647460938,
1.81611061096191,54.5255393981934,
3.54707288742065,52.8890953063965,
-11.1874179840088,25.5830078125000,
-7.08335638046265,-2.06488132476807,
19.0154991149902,-22.4511756896973,
33.1860694885254,-40.3004035949707,
20.6147499084473,-46.9574623107910,
7.59571266174316,-25.9096565246582,
17.0793247222900,23.8426246643066,
26.1996994018555,64.1399536132813,
0.326937198638916,64.3298950195313,
-43.2151718139648,33.9938774108887,
-56.8795242309570,7.92901134490967,
-24.1818504333496,5.33795928955078,
18.7069225311279,12.5162563323975,
35.1996421813965,11.5541191101074,
25.9705371856689,2.86790657043457,
11.4663639068604,-4.94734239578247,
-3.29308700561523,-3.28812861442566,
-26.0979003906250,9.57238578796387,
-48.5484008789063,19.4077720642090,
-54.3143157958984,10.4105377197266,
-45.3202476501465,-21.3703422546387,
-36.5426254272461,-58.3310890197754,
-25.0072937011719,-73.1961746215820,
7.14498090744019,-58.3027572631836,
50.1221733093262,-26.9572544097900,
65.8386840820313,7.71294546127319,
34.8554306030273,46.8955535888672,
-10.2169198989868,71.6745910644531,
-24.4157886505127,57.3381042480469,
-0.0712192505598068,12.0797653198242,
27.5363140106201,-18.9173564910889,
35.4978675842285,-4.11250495910645,
34.6747474670410,27.1212482452393,
36.5654029846191,23.2989768981934,
33.3700942993164,-11.6310214996338,
16.9190273284912,-23.8184032440186,
1.61279785633087,10.5518503189087,
1.61652028560638,41.6130371093750,
4.70993614196777,21.6818523406982,
-3.08328270912170,-19.3640708923340,
-19.3153572082520,-15.4536209106445,
-28.1397762298584,38.9334983825684,
-26.7304363250732,74.1004867553711,
-21.9073543548584,40.4984474182129,
-21.3848934173584,-28.5298500061035,
-18.6331233978272,-64.5842895507813,
-13.6694173812866,-50.3064041137695,
-15.2381439208984,-15.8298053741455,
-13.2913808822632,9.80433845520020,
6.25517463684082,25.8490371704102,
29.8430099487305,30.8103866577148,
26.7711715698242,13.3581628799438,
-2.54627656936646,-21.8795890808105,
-15.2763767242432,-38.6712989807129,
10.5239076614380,-14.6070938110352,
36.3279953002930,20.9577045440674,
17.3512516021729,25.6950187683105,
-24.9528408050537,-3.02474951744080,
-24.2618503570557,-31.9981479644775,
29.3690834045410,-33.6484298706055,
64.8147201538086,-14.9532165527344,
28.3749351501465,1.92640542984009,
-42.0075531005859,10.3675708770752,
-70.7475585937500,18.2270355224609,
-46.0449333190918,22.4648914337158,
-17.8831939697266,25.8189239501953,
-15.0378961563110,32.7876625061035,
-15.3952980041504,37.3828048706055,
3.42640972137451,30.7593517303467,
23.6347713470459,14.5407247543335,
22.8016242980957,10.5539703369141,
11.6244258880615,30.0366458892822,
13.9966545104980,45.0173606872559,
29.2956180572510,21.7638950347900,
34.1499633789063,-29.8231925964355,
18.6608695983887,-59.1129837036133,
2.37206530570984,-41.4995727539063,
-2.43901252746582,-17.2458667755127,
-2.48076963424683,-33.3041229248047,
0.731350541114807,-73.0982742309570,
11.3727245330811,-71.2684249877930,
26.0604972839355,-4.12117671966553,
35.4085578918457,68.9906387329102,
28.0856113433838,77.6123352050781,
9.95355319976807,22.4512462615967,
-3.01797437667847,-25.6311950683594,
-0.444852709770203,-20.1897277832031,
16.1391563415527,16.3513107299805,
36.4628295898438,32.2490196228027,
40.9861106872559,15.2770862579346,
14.7023830413818,-1.61648356914520,
-29.2512054443359,2.70944595336914,
-52.3909072875977,14.9220323562622,
-27.6763286590576,13.4296035766602,
17.5050773620605,-2.45227169990540,
32.6698760986328,-13.0467538833618,
2.74522972106934,-9.24077606201172,
-33.6356239318848,2.75624799728394,
-33.3253326416016,13.1962060928345,
1.87072670459747,24.2072238922119,
30.5908756256104,35.3049697875977,
20.9047870635986,35.7743873596191,
-9.99579048156738,18.3331775665283,
-29.4467964172363,-11.1070384979248,
-20.5448551177979,-28.0283031463623,
5.67417144775391,-10.5886716842651,
24.8987045288086,37.5866737365723,
18.7190151214600,79.0190200805664,
-9.89628219604492,73.9564056396484,
-38.5357246398926,18.2756938934326,
-40.3247261047363,-48.5895843505859,
-14.6567344665527,-76.7417602539063,
5.81767272949219,-52.4423065185547,
-5.66258192062378,-4.60552597045898,
-33.9893875122070,23.4866104125977,
-31.6240539550781,12.1176490783691,
18.7253417968750,-18.7224178314209,
72.5892333984375,-31.2009162902832,
77.2094802856445,-11.6525592803955,
32.3578186035156,19.1369686126709,
-13.8203716278076,21.2409191131592,
-28.1666221618652,-12.4195890426636,
-18.2208862304688,-44.0036354064941,
-9.03746986389160,-36.3204460144043,
-3.81635332107544,-0.776662349700928,
4.36109590530396,18.7271556854248,
5.19895315170288,12.6851606369019,
-12.0064849853516,14.5057411193848,
-28.3296318054199,35.8656692504883,
-17.1860580444336,44.1448287963867,
13.8542327880859,13.8677396774292,
26.2943553924561,-22.6262741088867,
3.88915467262268,-12.3438291549683,
-24.4689483642578,34.7533378601074,
-34.6479415893555,56.6593360900879,
-37.9413833618164,29.4248332977295,
-50.4158439636231,-1.27651381492615,
-59.5291404724121,1.55487227439880,
-33.7068557739258,9.42121791839600,
14.1609191894531,-13.4210653305054,
39.0741653442383,-39.7272071838379,
25.8178710937500,-20.9090461730957,
10.5487327575684,31.5114097595215,
17.2574081420898,54.5352172851563,
26.8213272094727,23.9306201934814,
11.4156951904297,-14.7470684051514,
-15.5976066589355,-18.7973308563232,
-24.2344493865967,-7.83013010025024,
-17.3273601531982,-13.0255088806152,
-18.4655075073242,-19.1716365814209,
-28.6222305297852,5.33174943923950,
-21.2620334625244,36.8068466186523,
15.5269737243652,26.5911483764648,
53.5371932983398,-15.8103828430176,
65.4968185424805,-28.8165149688721,
52.2514190673828,16.6316204071045,
29.7535705566406,68.8358383178711,
-4.88990545272827,66.5496215820313,
-48.9240188598633,22.2770919799805,
-76.7768249511719,-8.98640727996826,
-72.3958969116211,-6.04945611953735,
-46.4716606140137,0.0891063958406448,
-22.2621097564697,-9.89445400238037,
-6.11979818344116,-15.7634410858154,
5.61707210540772,-5.13510799407959,
7.47015523910523,-2.48879981040955,
-11.8170576095581,-25.4737186431885,
-32.9675102233887,-46.8930511474609,
-24.7141323089600,-30.6213169097900,
5.11066293716431,15.4462604522705,
9.87638187408447,45.1947326660156,
-25.1109046936035,24.4219188690186,
-46.5900802612305,-25.8701725006104,
-10.5090236663818,-55.4804992675781,
53.3671989440918,-44.0866165161133,
73.7638092041016,-7.65085029602051,
37.5378112792969,25.2378501892090,
3.73581814765930,34.6643104553223,
12.3796167373657,24.3932476043701,
32.5169448852539,18.2716770172119,
9.90788269042969,25.7403907775879,
-44.2529067993164,29.1187648773193,
-70.7640380859375,4.42041635513306,
-44.5587005615234,-30.8511772155762,
-3.21618652343750,-30.6728725433350,
12.5305137634277,13.8736572265625,
9.73353004455566,54.3880577087402,
12.5230398178101,35.5591049194336,
19.1052589416504,-31.7596855163574,
11.7976436614990,-80.5308761596680,
-6.30032920837402,-72.5720443725586,
-9.58017158508301,-37.8171501159668,
15.2078094482422,-14.2633514404297,
45.5314750671387,-1.31231594085693,
47.9644317626953,17.7353744506836,
23.5051403045654,38.5674743652344,
-4.49685382843018,48.1994781494141,
-17.9043922424316,48.3485488891602,
-11.3958187103271,47.1729316711426,
7.10220432281494,32.4463920593262,
15.4268274307251,-7.63305616378784,
3.81789112091064,-43.2899208068848,
-12.8759346008301,-31.6979007720947,
-9.09273910522461,12.3685302734375,
15.4624691009521,20.9850711822510,
27.4885807037354,-30.6019058227539,
8.02146053314209,-70.5861740112305,
-16.7113456726074,-29.2884445190430,
-6.96144866943359,48.4182662963867,
22.3906383514404,63.8026008605957,
21.1157417297363,-3.55952310562134,
-14.8636875152588,-65.2340927124023,
-28.4153938293457,-47.5472030639648,
6.69268894195557,16.2766761779785,
41.5525360107422,47.3804397583008,
13.5434522628784,28.6907176971436,
-55.8215599060059,7.78896427154541,
-91.8085327148438,3.76543474197388,
-67.0915222167969,-1.50568580627441,
-26.2605895996094,-16.8376159667969,
-10.7622280120850,-17.4404544830322,
-1.84010803699493,0.467583298683167,
28.0889472961426,7.55999660491943,
55.9720916748047,-9.77008056640625,
44.4971084594727,-23.0525321960449,
7.70065402984619,-10.0942945480347,
-7.54863882064819,14.7886762619019,
11.6076602935791,20.9033412933350,
31.5912113189697,15.3642673492432,
23.7388992309570,25.9356040954590,
-4.30066537857056,43.4520034790039,
-33.2305870056152,27.5972347259522,
-53.4515762329102,-21.3875255584717,
-54.2022705078125,-56.3181076049805,
-21.0475540161133,-50.7343559265137,
33.8315620422363,-32.6917381286621,
66.4378280639648,-34.2763328552246,
38.6751861572266,-41.4684715270996,
-18.1812419891357,-22.5646247863770,
-39.6068572998047,7.21086883544922,
-8.63964843750000,0.858620762825012,
26.6693134307861,-49.3237342834473,
22.2563896179199,-91.8366699218750,
-11.8385114669800,-75.6277313232422,
-30.8940792083740,-19.8911552429199,
-16.6903533935547,15.1036357879639,
4.89609241485596,4.93399572372437,
2.33567333221436,-22.7399044036865,
-18.6385955810547,-29.5131759643555,
-26.7526187896729,-12.5246448516846,
-3.35565090179443,7.72018337249756,
41.7063789367676,16.9962081909180,
71.8249053955078,21.0836429595947,
62.1647033691406,34.3209304809570,
20.7678012847900,49.8468704223633,
-17.2757759094238,47.6373443603516,
-22.3445701599121,15.9385166168213,
-5.27982425689697,-28.0894145965576,
4.62515354156494,-52.7928886413574,
-3.59587407112122,-38.7546653747559,
-10.1941070556641,-1.19098067283630,
2.05865955352783,24.3967666625977,
18.3387622833252,26.0986022949219,
7.35371541976929,17.2472305297852,
-28.9970455169678,11.2438163757324,
-50.6642227172852,5.02495479583740,
-29.0033950805664,-1.97947072982788,
14.3137893676758,-0.404771327972412,
35.1296501159668,15.6352796554565,
15.7298555374146,28.8855876922607,
-14.5151672363281,18.5998115539551,
-19.6072311401367,-5.86423015594482,
-2.47778654098511,-9.72481441497803,
12.2574253082275,17.3617534637451,
7.61322402954102,41.7811317443848,
-10.5645694732666,37.1429405212402,
-28.1958999633789,19.9097938537598,
-32.8374633789063,20.2076511383057,
-18.0252189636230,24.9422016143799,
6.59803009033203,4.68071174621582,
17.4714431762695,-34.4987945556641,
-1.18067741394043,-52.8940200805664,
-25.2348899841309,-36.2874526977539,
-15.7637901306152,-23.2353115081787,
25.2197399139404,-38.9121017456055,
53.7326927185059,-48.6203269958496,
34.5337677001953,-11.8526229858398,
-9.04504585266113,42.6152572631836,
-22.6860294342041,47.2412376403809,
1.99167668819428,-3.50578069686890,
24.6148738861084,-41.1044349670410,
15.7824821472168,-22.9333057403564,
-7.48846054077148,5.20505046844482,
-13.0395059585571,-11.0334014892578,
10.0915966033936,-53.0307807922363,
39.5418205261231,-55.4553604125977,
54.0132713317871,-6.78535938262939,
39.6797752380371,35.6204681396484,
3.89660024642944,32.2528381347656,
-26.9639549255371,13.0624771118164,
-26.0545825958252,21.6874294281006,
3.79155874252319,47.1983413696289,
23.1826801300049,51.9049263000488,
2.28680300712585,31.1459674835205,
-36.3179168701172,14.5570735931396,
-45.1166305541992,15.9561243057251,
-17.0784130096436,23.8396606445313,
3.33678674697876,28.7733993530273,
-12.5270557403564,30.8454418182373,
-45.7590751647949,29.4240226745605,
-64.0881118774414,15.2336015701294,
-63.5313186645508,-8.84439182281494,
-63.0571403503418,-21.5052833557129,
-59.0662117004395,-7.22422409057617,
-30.1153507232666,13.1466903686523,
15.6232357025146,22.1981601715088,
38.3820838928223,23.0294914245605,
14.1299304962158,24.9077568054199,
-29.2241878509522,21.6265659332275,
-42.7017059326172,5.70223093032837,
-13.8622932434082,-9.34391021728516,
29.6869850158691,-7.05003595352173,
58.5560379028320,5.47775030136108,
65.3986511230469,2.03086805343628,
49.5523452758789,-18.4756011962891,
16.3990192413330,-26.4603595733643,
-23.0237770080566,-5.88285827636719,
-47.7961006164551,8.32698249816895,
-44.3567504882813,-17.8177032470703,
-24.2498283386230,-68.6020355224609,
-7.40771245956421,-91.6430282592773,
-4.32835006713867,-70.1717224121094,
-5.56527519226074,-37.5514755249023,
-3.46167087554932,-26.3144149780273,
0.845201373100281,-29.0960655212402,
6.85475015640259,-16.9704494476318,
10.8133239746094,10.4316902160645,
13.2116365432739,29.7843475341797,
21.1693992614746,30.2742710113525,
38.2220687866211,23.9166889190674,
52.6693038940430,16.1455707550049,
46.9770507812500,-2.75564670562744,
19.6025009155273,-34.6157455444336,
-4.41757869720459,-58.2588806152344,
-4.17987632751465,-54.0990829467773,
8.08038425445557,-34.8169021606445,
2.98622083663940,-23.5520935058594,
-15.5768775939941,-17.5323467254639,
-11.7458219528198,-1.75239646434784,
23.0673217773438,24.5724754333496,
51.1856155395508,32.0918960571289,
42.1419143676758,10.6526031494141,
15.9497079849243,-8.22581386566162,
12.0171880722046,8.52688980102539,
24.8813953399658,42.9464302062988,
15.9724903106689,46.6715927124023,
-17.0620365142822,6.06613302230835,
-28.7236652374268,-35.9408340454102,
8.83082008361816,-33.0005722045898,
52.2985305786133,6.20916271209717,
50.9210128784180,34.0261650085449,
14.1825141906738,19.9981040954590,
-1.79605865478516,-17.1453857421875,
25.9443187713623,-40.1506423950195,
52.2046356201172,-36.0115890502930,
35.0575370788574,-13.0307302474976,
-9.00082683563232,11.7473745346069,
-35.1272125244141,26.7171726226807,
-29.4290866851807,22.7725582122803,
-13.5864238739014,2.61075019836426,
-6.82117223739624,-19.1251525878906,
2.70757555961609,-22.0962600708008,
23.2203941345215,0.500306606292725,
36.7422409057617,33.5293426513672,
15.1940212249756,47.8600692749023,
-28.1797866821289,28.4265270233154,
-49.0913848876953,-10.9724731445313,
-17.8471527099609,-40.4234352111816,
42.1759719848633,-40.0171737670898,
78.7393569946289,-12.2582244873047,
61.9976844787598,19.9444713592529,
16.0004997253418,40.0341300964356,
-15.5734262466431,42.5362129211426,
-15.2376432418823,32.3872032165527,
1.60222482681274,15.3876476287842,
14.9495601654053,2.88352966308594,
22.3392200469971,5.97847700119019,
34.3290824890137,14.6569328308105,
45.5008392333984,14.8333644866943,
36.9278335571289,6.40678930282593,
-3.23243975639343,7.04115962982178,
-54.5284347534180,25.1787776947022,
-79.1491241455078,37.2377548217773,
-58.4464797973633,10.5541400909424,
-16.4808826446533,-40.8404045104981,
8.29164505004883,-66.8692779541016,
-3.41726207733154,-41.5924491882324,
-32.2136878967285,-0.439703226089478,
-43.8849678039551,2.46066141128540,
-28.6962451934814,-30.5056552886963,
-3.77461838722229,-42.4508323669434,
4.78134775161743,3.88853788375855,
-8.68048286437988,66.6307678222656,
-28.2049102783203,79.9317703247070,
-38.1802482604981,36.1568031311035,
-36.3112792968750,-5.25523328781128,
-38.8016128540039,-3.04638981819153,
-53.4861373901367,15.0240087509155,
-61.4591369628906,-0.311780571937561,
-35.7982101440430,-44.1058006286621,
14.5048103332520,-64.2623138427734,
43.9319267272949,-35.8748245239258,
26.9269008636475,-0.895984113216400,
-9.89365196228027,-1.02765238285065,
-20.2188167572022,-17.8918952941895,
0.765910923480988,-9.33245372772217,
13.6024818420410,26.7709465026855,
1.69353294372559,48.5864601135254,
-0.846728086471558,36.1440124511719,
28.4921627044678,18.5191860198975,
50.2215538024902,23.1686458587647,
22.4042167663574,27.8419361114502,
-32.3352928161621,7.19117927551270,
-44.3581504821777,-23.4846534729004,
4.28957843780518,-26.3651752471924,
57.9784774780273,0.402932882308960,
58.2951545715332,16.4824428558350,
23.4441738128662,-2.77819538116455,
-1.51291525363922,-32.0920410156250,
-10.9819316864014,-31.1314239501953,
-26.9664802551270,-4.35567617416382,
-43.5842437744141,13.7923603057861,
-27.9971904754639,8.01007652282715,
13.0304574966431,-2.03858613967896,
23.3660964965820,7.16072416305542,
-23.9262237548828,33.1775245666504,
-76.9312438964844,46.1310272216797,
-68.4361877441406,26.0297698974609,
-14.9561882019043,-12.1422119140625,
11.5493288040161,-30.8745803833008,
-24.2269325256348,-17.8164730072022,
-70.0944976806641,4.78097009658814,
-57.9175987243652,1.37346994876862,
3.45851302146912,-30.9583034515381,
46.5991058349609,-60.5051879882813,
39.4630393981934,-62.1975555419922,
11.4721517562866,-47.2401542663574,
3.37706398963928,-38.2230186462402,
13.3959655761719,-30.8038635253906,
8.64571857452393,-12.9143695831299,
-17.0015048980713,7.97914600372314,
-29.8584194183350,7.11037826538086,
-3.44398665428162,-15.1363668441772,
48.4217300415039,-23.9386711120605,
80.5146179199219,4.71375894546509,
66.8303756713867,48.4383010864258,
22.2065811157227,68.7040939331055,
-10.2949228286743,57.9897308349609,
-6.92658376693726,38.1307182312012,
12.9177198410034,27.1451644897461,
7.45690631866455,17.2305622100830,
-34.0637588500977,-1.18902313709259,
-73.0134124755859,-19.2063274383545,
-60.0952301025391,-14.9823675155640,
0.205504179000855,9.63905620574951,
43.5728874206543,37.6879997253418,
15.9914150238037,46.3751869201660,
-53.6013641357422,29.6620140075684,
-85.7361831665039,-0.720198094844818,
-45.4294700622559,-17.8459796905518,
16.3918590545654,-13.4600524902344,
30.3310890197754,-3.46848535537720,
-8.16024208068848,-7.48342561721802,
-35.2521667480469,-21.0528011322022,
-13.3018264770508,-25.2622013092041,
30.4947490692139,-13.9047098159790,
42.0922737121582,-12.8889398574829,
15.9794616699219,-33.2475585937500,
-8.18124389648438,-48.7624397277832,
0.518362045288086,-25.4058494567871,
33.0467720031738,19.0527019500732,
57.6677093505859,34.2082290649414,
61.7724189758301,8.92246246337891,
47.4789772033691,-9.64089870452881,
24.2141799926758,19.0284976959229,
4.97914314270020,67.5292739868164,
-3.38997793197632,78.1114501953125,
-0.143920540809631,41.0778808593750,
9.86505126953125,3.88677072525024,
20.9129295349121,3.15528464317322,
38.3166732788086,21.5939865112305,
58.3849449157715,27.0654239654541,
62.3426017761231,20.0217170715332,
38.9210166931152,23.8770847320557,
1.08036708831787,35.6053237915039,
-28.4795284271240,37.5453567504883,
-40.4002990722656,25.5312042236328,
-42.6787147521973,18.1571960449219,
-38.6463356018066,22.2414760589600,
-26.1777286529541,28.0484981536865,
-12.5110473632813,28.3852901458740,
-16.6193637847900,34.3533668518066,
-36.9884872436523,46.6227912902832,
-49.6260681152344,44.2124176025391,
-29.8364124298096,15.3506221771240,
9.30487632751465,-16.9074440002441,
32.8908309936523,-18.7016925811768,
25.0518436431885,-3.64954280853272,
-2.59581398963928,-14.4853153228760,
-23.8164520263672,-52.5545654296875,
-24.8857460021973,-71.5196685791016,
-2.14982056617737,-43.0718269348145,
24.0163612365723,-2.84850597381592,
26.0382537841797,-1.79768931865692,
0.921893835067749,-37.4531631469727,
-22.1272830963135,-51.0113067626953,
-14.2380361557007,-12.9297561645508,
9.13563156127930,40.7155838012695,
9.70984840393066,59.8422279357910,
-23.7725811004639,36.9130668640137,
-48.8074302673340,-1.44359731674194,
-32.6699943542481,-24.9922256469727,
3.91580939292908,-19.0629520416260,
21.2188205718994,14.5456571578980,
21.4595508575439,43.6550102233887,
31.0199127197266,32.9940795898438,
45.6904983520508,-13.7852277755737,
34.5549964904785,-41.1048011779785,
-2.17040824890137,-9.56002807617188,
-19.4018421173096,49.9148521423340,
4.20508480072022,60.6227645874023,
27.5345478057861,3.45867037773132,
8.49131393432617,-57.1837806701660,
-28.3468017578125,-67.1962051391602,
-23.2057285308838,-44.5732955932617,
28.0888519287109,-27.0679149627686,
60.5674018859863,-18.6881408691406,
33.5704956054688,-3.02136898040772,
-14.5321817398071,9.67842388153076,
-28.1114883422852,-11.4510507583618,
-6.68017959594727,-50.9273490905762,
9.56978988647461,-59.3483467102051,
2.93828272819519,-29.0904502868652,
-7.52283668518066,-10.0859594345093,
-6.19608402252197,-28.1094474792480,
0.821525216102600,-40.5290489196777,
1.67564797401428,2.71593213081360,
1.30658650398254,66.8488388061523,
3.31315183639526,69.5417098999023,
0.307512402534485,6.68546485900879,
-7.20750093460083,-42.1616058349609,
-4.19720649719238,-18.2680778503418,
10.9320325851440,40.7903709411621,
13.9042139053345,50.1689224243164,
-10.4440908432007,-3.59489727020264,
-39.4148597717285,-54.7100601196289,
-44.2117156982422,-52.8538932800293,
-26.7257270812988,-20.0089969635010,
-11.4818849563599,-8.93077087402344,
-9.38707828521729,-36.7363929748535,
-3.87864518165588,-68.9173202514648,
16.0522632598877,-68.1110763549805,
33.6338081359863,-25.7483501434326,
27.6947650909424,35.5586547851563,
4.73593044281006,74.2661666870117,
-12.5160655975342,63.2831344604492,
-12.1709547042847,12.9746379852295,
-0.371900737285614,-34.6648254394531,
9.29956722259522,-40.3994750976563,
6.16557264328003,-13.7012767791748,
-10.7220163345337,-4.52181911468506,
-23.7331848144531,-32.3465957641602,
-10.3465833663940,-60.0557479858398,
22.4652748107910,-41.7277679443359,
40.3008766174316,14.9204740524292,
23.4524078369141,54.3276290893555,
-7.92504978179932,41.0633392333984,
-11.6799898147583,-0.923603415489197,
14.2041168212891,-29.2724552154541,
33.0018882751465,-34.0534629821777,
21.8462829589844,-32.1858444213867,
1.99721062183380,-29.9191989898682,
-4.90264749526978,-17.6358585357666,
-5.75878381729126,0.672261714935303,
-15.7003736495972,-3.93191170692444,
-22.4728679656982,-36.6753921508789,
-8.18005371093750,-64.3446502685547,
12.7618427276611,-50.7600517272949,
6.16309499740601,-4.83395338058472,
-27.1208782196045,23.6489353179932,
-40.5617256164551,6.04952383041382,
-5.36113214492798,-35.7495994567871,
45.5144462585449,-50.0713005065918,
60.1202049255371,-19.3321857452393,
31.2768096923828,29.2514820098877,
2.78842568397522,53.8429718017578,
5.63114070892334,33.5030326843262,
23.6381149291992,-6.74550628662109,
30.2503681182861,-25.8062877655029,
27.1026134490967,-3.66629147529602,
29.7347640991211,38.2461090087891,
32.6998977661133,59.0303115844727,
18.1430625915527,39.6105690002441,
-7.25739574432373,-0.464471578598022,
-9.65863609313965,-30.9681148529053,
27.6315593719482,-33.4697151184082,
70.0378265380859,-14.9926614761353,
65.5010986328125,10.5639686584473,
13.1024990081787,31.1103210449219,
-33.3729362487793,37.4325256347656,
-30.4661140441895,25.2818565368652,
5.61624765396118,0.525205552577972,
24.8237514495850,-24.1407852172852,
3.34613060951233,-32.0769805908203,
-23.9525070190430,-13.7629356384277,
-20.5666027069092,19.1495780944824,
6.97979545593262,36.4924774169922,
26.0406436920166,14.1030235290527,
16.4759445190430,-29.6470260620117,
-1.85589933395386,-47.3997650146484,
-1.95625603199005,-24.4717960357666,
18.8477783203125,1.63529896736145,
36.5768890380859,-11.0505504608154,
30.4450016021729,-51.4844169616699,
4.96493434906006,-62.8471603393555,
-13.4513254165649,-25.3668441772461,
-10.2123069763184,17.1322822570801,
2.06205415725708,17.7561264038086,
-6.80474805831909,-11.1170063018799,
-44.2056236267090,-22.3840255737305,
-69.9845733642578,-8.72105312347412,
-44.9318313598633,-3.51796221733093,
18.5211811065674,-19.8691139221191,
63.3481178283691,-28.2132530212402,
51.5300025939941,-6.55940532684326,
8.57037258148193,13.9661664962769,
-13.2363090515137,-4.49438524246216,
1.61549103260040,-47.0659255981445,
23.5270023345947,-60.1685409545898,
29.1707553863525,-20.9042396545410,
23.8794326782227,31.7205333709717,
20.0288219451904,51.2192039489746,
17.2762660980225,35.1014328002930,
10.0665063858032,14.0836105346680,
8.65885162353516,2.93646955490112,
23.9957447052002,-2.78509902954102,
43.0862007141113,-4.63030004501343,
43.5131340026856,1.38888669013977,
21.4447402954102,12.3859338760376,
-1.41604363918304,19.3349151611328,
-10.1711626052856,18.4448223114014,
-8.62921714782715,18.1837253570557,
-17.1459045410156,24.8358421325684,
-36.8617324829102,25.8983898162842,
-50.0833129882813,10.6883420944214,
-40.3699417114258,-9.63767242431641,
-12.5164623260498,-13.0703420639038,
12.0444650650024,5.35411500930786,
11.9842948913574,32.5473976135254,
-8.65359020233154,50.8920707702637,
-22.7364501953125,44.1407012939453,
-9.34928798675537,16.3424873352051,
17.6757907867432,-15.4130277633667,
27.5144195556641,-23.5984954833984,
14.9221200942993,0.616729259490967,
4.64446878433228,32.0275573730469,
13.5016736984253,31.8750820159912,
27.3347778320313,-5.52029037475586,
21.6421298980713,-36.7539176940918,
4.34691095352173,-29.3932476043701,
2.07433915138245,1.03042840957642,
21.2660732269287,15.7839584350586,
30.3971939086914,13.4873571395874,
11.5117053985596,24.4276618957520,
-19.2722740173340,54.4303779602051,
-35.4212188720703,68.9499130249023,
-37.7840805053711,40.4518089294434,
-35.4738388061523,-6.95787334442139,
-21.3480377197266,-27.0404129028320,
9.19998359680176,-21.2271518707275,
36.2935714721680,-20.2315406799316,
34.1643981933594,-26.8094043731689,
11.1854524612427,-9.87329578399658,
-3.55918765068054,34.5749435424805,
-3.51292634010315,64.0727233886719,
-17.0524406433105,48.1713600158691,
-49.3526000976563,16.2104015350342,
-60.9205169677734,7.07240819931030,
-31.7995605468750,9.80657958984375,
-3.41454052925110,-9.43789863586426,
-18.4165477752686,-38.6755409240723,
-47.2714233398438,-29.1429080963135,
-33.3920288085938,20.7724685668945,
17.5840320587158,47.3336486816406,
41.7918128967285,5.42008399963379,
11.3175468444824,-54.2795982360840,
-22.6228351593018,-63.3437576293945,
-14.6385946273804,-27.0478019714355,
4.35392236709595,-2.37187218666077,
-15.3433904647827,-14.5069408416748,
-52.2727432250977,-31.1521759033203,
-44.1485404968262,-19.4841403961182,
5.46573066711426,9.95727920532227,
30.8853416442871,27.6635932922363,
5.48052501678467,26.8707637786865,
-18.8560142517090,10.9698095321655,
0.721725702285767,-13.7811536788940,
35.1723289489746,-28.4424228668213,
30.8487110137939,-4.61707305908203,
-0.870165288448334,48.8263931274414,
-11.2002210617065,78.6540298461914,
10.0814285278320,58.3053321838379,
18.9609909057617,27.9670352935791,
-2.30878615379334,32.4962387084961,
-15.3688364028931,50.1662559509277,
5.33662319183350,28.0366077423096,
26.5453910827637,-32.5686187744141,
10.9042186737061,-58.5611457824707,
-21.6650886535645,-13.7061071395874,
-23.9840660095215,51.1262779235840,
6.54291963577271,64.4459609985352,
23.8204441070557,34.6014747619629,
1.61497640609741,19.3717365264893,
-36.2025566101074,33.2399139404297,
-52.2748947143555,36.3317489624023,
-45.5423278808594,7.51132297515869,
-41.3414459228516,-22.4461765289307,
-43.8606185913086,-20.8840332031250,
-34.8995971679688,-1.60080826282501,
-6.99763727188110,5.97547388076782,
22.4104576110840,-1.94832193851471,
36.7574386596680,1.35226500034332,
31.4354343414307,22.7557201385498,
15.2982816696167,44.0727386474609,
-1.15551531314850,53.2127227783203,
-15.7415752410889,56.0248718261719,
-34.1487808227539,53.8470840454102,
-53.7575798034668,32.9713668823242,
-56.0289268493652,-2.04480695724487,
-29.8816375732422,-19.6044692993164,
11.5677108764648,-1.55250620841980,
29.2037696838379,27.4727287292480,
6.47781467437744,29.5872650146484,
-18.5818862915039,5.84992074966431,
-0.309561252593994,-4.51995229721069,
51.5651473999023,14.4271879196167,
69.6685104370117,28.3619480133057,
27.0476150512695,9.12674236297607,
-26.2020244598389,-19.6030158996582,
-35.7280082702637,-14.1057376861572,
-10.5767936706543,22.5625114440918,
0.977624297142029,42.8459854125977,
-10.7005290985107,25.0462684631348,
-5.10018730163574,-4.87904167175293,
32.3265266418457,-11.4479789733887,
60.2651710510254,0.473575562238693,
49.1379013061523,2.96010112762451,
27.0797233581543,-8.71521854400635,
23.5805282592773,-12.6729831695557,
15.1330480575562,-3.51559019088745,
-28.6162548065186,3.44909429550171,
-70.8081130981445,-3.07394957542419,
-42.9317703247070,-18.2004051208496,
43.3594055175781,-28.1270351409912,
85.8114624023438,-22.8487091064453,
28.9612102508545,2.26196908950806,
-53.7236633300781,32.0742568969727,
-57.0482864379883,36.1287002563477,
14.4978971481323,3.98892068862915,
54.4368019104004,-28.2118377685547,
12.5157375335693,-14.7406702041626,
-40.8441619873047,41.7030448913574,
-26.1998748779297,73.2108001708984,
28.4729766845703,34.6458663940430,
41.9954414367676,-36.0579147338867,
-1.75720286369324,-66.2462005615234,
-39.7297439575195,-38.9674301147461,
-22.1249504089355,3.28325319290161,
20.7717323303223,25.7428054809570,
26.6827411651611,29.0512924194336,
-17.2913208007813,23.1967811584473,
-63.6948585510254,8.41522979736328,
-69.0666198730469,-9.44173049926758,
-35.3800926208496,-11.3520889282227,
7.54163885116577,2.82763099670410,
22.4278755187988,-0.172748774290085,
2.14121580123901,-37.9675865173340,
-16.9739742279053,-74.4308776855469,
5.92711687088013,-65.3177185058594,
53.4549751281738,-23.7277011871338,
68.2574920654297,-0.838022768497467,
22.9915332794189,-10.1932964324951,
-32.7953453063965,-7.73954439163208,
-30.6958503723145,23.3681449890137,
19.3980827331543,45.7939414978027,
40.8054771423340,24.5306720733643,
3.64324760437012,-14.4711284637451,
-33.2082481384277,-15.4373331069946,
-9.48552608489990,21.0587711334229,
45.9381484985352,43.7957916259766,
62.3152618408203,26.0256156921387,
22.3261013031006,1.69279801845551,
-20.4173736572266,8.89999008178711,
-29.0644207000732,33.3686561584473,
-26.7415084838867,34.3095588684082,
-44.9585456848145,5.47460842132568,
-65.6741638183594,-25.0305023193359,
-55.0797348022461,-37.7325019836426,
-16.5625629425049,-30.5337104797363,
10.9239091873169,-10.2140007019043,
9.41920566558838,17.1313533782959,
-3.37089180946350,40.1465492248535,
-14.6290855407715,46.1129875183106,
-28.9502601623535,32.4934539794922,
-39.6898231506348,15.1501922607422,
-29.9664764404297,4.71922683715820,
-2.94764542579651,-2.81886458396912,
16.9071884155273,-3.31778597831726,
13.2145767211914,18.5358619689941,
1.98354351520538,50.3369140625000,
10.0189132690430,54.7524452209473,
31.4129047393799,21.9218578338623,
40.4152488708496,-12.0698547363281,
41.2942199707031,-11.6578712463379,
49.8233108520508,7.19024658203125,
62.0798301696777,2.55005764961243,
47.8165473937988,-24.9672470092773,
12.2768783569336,-25.4869651794434,
-3.50110054016113,11.5217380523682,
13.1164331436157,33.5717430114746,
23.7243022918701,4.43450212478638,
-4.70704221725464,-30.4675083160400,
-46.7280387878418,-13.7858152389526,
-51.7212524414063,31.1748886108398,
-14.3562564849854,30.3255290985107,
16.7642803192139,-27.0331859588623,
16.9479618072510,-66.5387268066406,
11.5516901016235,-37.4740219116211,
27.4607295989990,14.4961786270142,
53.8237304687500,22.2704830169678,
69.9326477050781,-2.87882566452026,
74.4411773681641,1.82173645496368,
60.4804725646973,43.2092361450195,
16.2954196929932,58.1272544860840,
-43.2305297851563,20.1289100646973,
-60.8095054626465,-22.9319324493408,
-11.0974073410034,-21.4807472229004,
51.6271514892578,3.18284988403320,
50.7938194274902,4.42059516906738,
-14.4755325317383,-15.8805532455444,
-67.6656417846680,-16.6531677246094,
-61.8600120544434,3.07878947257996,
-36.0567855834961,2.66396117210388,
-27.6997871398926,-30.7787933349609,
-15.2603940963745,-54.4002380371094,
29.1912822723389,-31.9721546173096,
73.7561264038086,5.01224517822266,
65.9806900024414,13.4214248657227,
16.0146961212158,8.21860694885254,
-19.9171733856201,29.5743865966797,
-16.8896045684814,69.0433883666992,
-8.14305973052979,72.4747009277344,
-14.8785343170166,21.8968372344971,
-11.3812112808228,-30.1492309570313,
19.0852451324463,-19.9165496826172,
40.4742813110352,38.9962615966797,
13.4294843673706,76.5307769775391,
-37.3354721069336,53.5627403259277,
-53.4691085815430,-2.22423768043518,
-30.1373329162598,-42.7477111816406,
-7.55521726608276,-42.1631050109863,
-10.3306913375855,-13.1810922622681,
-20.8964900970459,11.5374975204468,
-21.5390319824219,5.23064994812012,
-18.2456970214844,-21.3822898864746,
-14.8766832351685,-33.3602066040039,
-0.668193101882935,-8.75141334533691,
30.8687877655029,25.3042240142822,
52.0791320800781,19.3861770629883,
33.8340492248535,-26.1377124786377,
-3.32855463027954,-54.8027381896973,
-26.0601654052734,-25.9280700683594,
-32.5084114074707,21.7884140014648,
-42.9753341674805,18.6177444458008,
-50.5221481323242,-33.6077804565430,
-28.0957794189453,-68.8752059936523,
16.1309967041016,-44.0006065368652,
36.6870689392090,-0.267433404922485,
11.7366046905518,0.542136967182159,
-18.6332283020020,-35.2508392333984,
-9.61492824554443,-51.2200393676758,
22.6253623962402,-17.4218120574951,
27.1200675964355,29.0031223297119,
2.35915732383728,35.9217758178711,
2.40009522438049,6.24806594848633,
49.2289962768555,-16.9260692596436,
94.0609893798828,-5.56931591033936,
78.5673522949219,25.0355587005615,
16.9828109741211,41.1637039184570,
-31.5580368041992,29.0925064086914,
-31.5255279541016,7.12791728973389,
-5.96177053451538,8.18616104125977,
11.2357721328735,29.8144531250000,
11.7599401473999,35.6129302978516,
7.19166469573975,-0.796052455902100,
2.20861887931824,-52.8401756286621,
-1.39925551414490,-58.7972259521484,
1.58896589279175,2.13177824020386,
7.29760456085205,70.8592453002930,
-1.81565320491791,72.8383941650391,
-30.2905158996582,12.3742790222168,
-51.3342933654785,-37.7902641296387,
-44.5751304626465,-30.1529064178467,
-24.3874874114990,3.75173091888428,
-24.6178359985352,12.4873285293579,
-44.7985534667969,-2.62036871910095,
-52.5800056457520,-2.12914609909058,
-25.4264106750488,30.2737312316895,
8.06613922119141,61.3180694580078,
8.16181087493897,58.3271217346191,
-18.5722751617432,30.0058078765869,
-37.4889678955078,8.59507083892822,
-30.7476711273193,10.8168210983276,
-12.3334207534790,24.1821575164795,
6.86463451385498,27.5086994171143,
28.6975727081299,11.8107833862305,
51.3087539672852,-13.0880203247070,
58.8266296386719,-20.3631706237793,
40.1948242187500,10.6677122116089,
12.8618335723877,52.5801506042481,
-4.53716897964478,53.2882575988770,
-12.9290981292725,0.345860958099365,
-20.4711227416992,-56.8849830627441,
-12.8985052108765,-64.1513595581055,
24.6002044677734,-27.4278182983398,
67.9431915283203,0.647681176662445,
71.9127197265625,-4.42593383789063,
35.2720298767090,-12.0029621124268,
9.48154926300049,5.37897491455078,
27.7845954895020,28.8677768707275,
55.1092529296875,27.3530368804932,
29.5955123901367,9.06381034851074,
-39.8758430480957,3.55070137977600,
-81.3037719726563,14.9028091430664,
-56.0651588439941,24.1731929779053,
-3.45502686500549,23.4754142761230,
13.7649965286255,19.1293010711670,
-2.99694538116455,11.7285652160645,
-14.4785099029541,-4.48763132095337,
-10.3674459457397,-19.9796772003174,
-13.1715526580811,-16.4658088684082,
-32.7593994140625,-0.402075260877609,
-40.8327217102051,-3.58809971809387,
-22.5302200317383,-31.4329414367676,
-1.03183031082153,-41.7665481567383,
-9.16312503814697,-10.6742296218872,
-38.5010299682617,21.1933593750000,
-51.1408615112305,1.55671119689941,
-28.5440101623535,-44.6429710388184,
11.1342887878418,-48.4239273071289,
43.4382133483887,7.14274454116821,
55.5392990112305,53.7788276672363,
39.2410774230957,34.1028671264648,
9.30590057373047,-16.0073146820068,
-5.03844308853149,-23.3286972045898,
12.9596166610718,16.7692794799805,
46.0499267578125,36.9526100158691,
61.6101531982422,4.73613214492798,
48.1894378662109,-37.1922073364258,
23.2726917266846,-39.1642189025879,
3.00371360778809,-9.55721092224121,
-12.5162410736084,14.1531019210815,
-22.3790607452393,25.3441772460938,
-14.5633935928345,43.0813865661621,
3.90698862075806,63.4385185241699,
-3.24040961265564,57.1497230529785,
-39.1946792602539,16.1760673522949,
-59.5496292114258,-26.1050033569336,
-26.1472320556641,-42.1332740783691,
33.5522193908691,-42.6617393493652,
62.2906837463379,-39.2308807373047,
52.1343383789063,-17.2350997924805,
39.2782516479492,29.8856449127197,
40.7006607055664,63.3442802429199,
27.7569656372070,41.8390769958496,
-8.76469612121582,-13.2007522583008,
-29.0887107849121,-37.3026237487793,
-4.01046371459961,-5.99537944793701,
24.2074317932129,29.9585323333740,
1.14531028270721,22.1089820861816,
-53.9150085449219,-3.58292460441589,
-71.7675018310547,4.94806337356567,
-39.4172477722168,44.3735542297363,
-12.2169237136841,51.2961196899414,
-27.1612834930420,1.12318873405457,
-46.4228820800781,-59.0007743835449,
-22.1118221282959,-73.4182739257813,
25.4911537170410,-43.1457710266113,
37.9001464843750,-12.0819053649902,
2.72693204879761,-3.09626007080078,
-29.3142299652100,-5.03374767303467,
-24.6291007995605,-6.23067617416382,
0.700935006141663,-11.8140745162964,
12.8441524505615,-28.5663051605225,
15.2810144424438,-39.7061882019043,
18.8790645599365,-29.8412513732910,
12.0695838928223,-1.38804531097412,
-17.7062988281250,27.4347515106201,
-48.9536895751953,40.7912330627441,
-45.7771530151367,31.4848594665527,
0.700983762741089,10.5618543624878,
50.3069686889648,-3.03282046318054,
57.4791717529297,0.301131695508957,
26.6897125244141,13.6822471618652,
-4.77312898635864,23.8197555541992,
-11.7584466934204,26.8358955383301,
-4.39900064468384,34.8040809631348,
-8.55674648284912,46.2927894592285,
-36.4535331726074,43.2898483276367,
-71.1537094116211,11.8715972900391,
-80.9573974609375,-32.6111450195313,
-53.3899879455566,-57.7823677062988,
-9.56065940856934,-48.6937026977539,
14.7753944396973,-26.8088264465332,
3.59974741935730,-18.1438961029053,
-16.3438377380371,-29.7545108795166,
-4.98877620697022,-43.0119400024414,
44.8773651123047,-37.5938453674316,
92.4421539306641,-7.13094615936279,
92.9263153076172,21.9882431030273,
47.6346893310547,23.6618995666504,
0.719576358795166,-4.42196702957153,
-9.82168388366699,-34.1164627075195,
9.57186317443848,-37.0110626220703,
25.1919708251953,-19.8601760864258,
22.7398586273193,-11.4956178665161,
14.9171514511108,-16.9961757659912,
11.4680624008179,-12.6945762634277,
2.79766058921814,19.3694057464600,
-15.8839378356934,49.6689949035645,
-28.5449962615967,38.4561080932617,
-13.8095340728760,-3.49632382392883,
18.2104454040527,-20.4685611724854,
33.0953598022461,22.4663391113281,
13.8254642486572,89.3100585937500,
-17.9275798797607,112.700706481934,
-34.6202239990234,69.8488540649414,
-31.4464263916016,-2.92196130752563,
-26.7248668670654,-53.0581092834473,
-23.7289924621582,-57.7157249450684,
-11.9478769302368,-29.0616092681885,
10.8806962966919,9.81085681915283,
28.2913646697998,36.5179901123047,
24.8527584075928,34.1073570251465,
3.25348520278931,6.22706890106201,
-20.5552101135254,-25.1628780364990,
-33.8578605651856,-36.3500022888184,
-31.5890350341797,-25.3808956146240,
-15.1526985168457,-6.38239145278931,
8.21946239471436,9.15284347534180,
23.1772193908691,11.8924016952515,
16.6638069152832,-0.310096025466919,
-2.33294820785522,-19.8401355743408,
-14.3094396591187,-31.6761779785156,
-10.6216316223145,-15.0933780670166,
4.59490156173706,22.1799488067627,
14.8339624404907,48.5950088500977,
11.2145700454712,39.6708297729492,
-7.79173183441162,1.96038889884949,
-30.0639209747314,-35.3827018737793,
-38.5332260131836,-48.3971366882324,
-23.4418029785156,-33.6173667907715,
2.37422060966492,-1.54450213909149,
9.64330673217773,23.8980693817139,
-11.6303672790527,20.9983196258545,
-32.2382469177246,-8.40464687347412,
-20.5261459350586,-36.8333740234375,
14.3425045013428,-33.0239219665527,
28.4143981933594,-4.66371297836304,
0.761223316192627,14.3588361740112,
-39.2861671447754,8.77581596374512,
-52.6238899230957,0.285157799720764,
-36.8523674011231,15.3103256225586,
-22.2961826324463,42.0603027343750,
-27.5958118438721,49.1305122375488,
-35.9860038757324,31.6699409484863,
-28.2968692779541,11.3586578369141,
-6.63208580017090,2.60189509391785,
17.8316078186035,-1.89744532108307,
36.2534828186035,-12.2801151275635,
42.5798530578613,-18.9874801635742,
28.0596332550049,-6.87472963333130,
-0.286096602678299,18.7074508666992,
-16.1868515014648,37.4192619323731,
-4.85875844955444,39.9785079956055,
12.4281415939331,27.2237529754639,
9.04356193542481,6.99747276306152,
-7.78561115264893,-13.8120880126953,
-5.84823274612427,-19.5767860412598,
24.2642440795898,-7.66352653503418,
44.5469017028809,0.880168616771698,
29.0656414031982,-13.5385828018188,
-5.28746509552002,-34.3628654479981,
-20.9368114471436,-27.1312294006348,
-14.6074342727661,14.4485778808594,
-7.80333375930786,43.5101776123047,
-10.0077123641968,22.1667079925537,
-9.48211193084717,-22.4362144470215,
-1.44274747371674,-27.9580993652344,
3.43340921401978,17.5176734924316,
1.78193640708923,62.0692749023438,
2.78987288475037,64.8907623291016,
12.2562036514282,43.0580863952637,
13.4502620697021,31.6072044372559,
-4.73529052734375,29.9630832672119,
-31.8234272003174,11.6391181945801,
-48.2971267700195,-17.5484066009522,
-49.9259262084961,-20.3019866943359,
-42.4601936340332,12.1743822097778,
-24.3641414642334,38.8667602539063,
-2.11093759536743,34.1848487854004,
3.74652957916260,19.5626201629639,
-16.6563796997070,27.1885566711426,
-35.9183082580566,42.9010734558106,
-20.3754577636719,29.5638217926025,
20.7297668457031,-2.13292074203491,
39.0657272338867,-8.85434818267822,
7.19827461242676,20.0942916870117,
-46.4503288269043,36.9571571350098,
-72.9555130004883,11.4822635650635,
-59.6139144897461,-23.4884281158447,
-31.0919265747070,-14.0894737243652,
-7.72358036041260,23.4336547851563,
5.17226219177246,26.0712356567383,
6.21287202835083,-24.8967590332031,
-0.989154338836670,-75.7020568847656,
-1.32855403423309,-70.0114898681641,
21.6112785339355,-22.5290412902832,
49.8891181945801,18.2594146728516,
50.2872047424316,33.9554443359375,
11.5200614929199,45.5430374145508,
-37.6320457458496,55.6104698181152,
-64.4415283203125,40.7671928405762,
-62.1585121154785,-9.27324199676514,
-44.6496429443359,-56.3400688171387,
-23.5186500549316,-63.4782600402832,
0.718189477920532,-40.8646316528320,
24.6595325469971,-25.1148891448975,
38.9715232849121,-24.5495605468750,
43.8331794738770,-13.6020193099976,
40.4505386352539,22.2504920959473,
23.0100212097168,61.8734703063965,
-12.3052167892456,70.8560333251953,
-46.8741836547852,45.6522979736328,
-57.0691413879395,19.1443881988525,
-41.7431335449219,13.0130586624146,
-22.7699985504150,27.7998657226563,
-17.2532024383545,44.8838233947754,
-33.3778686523438,41.7260246276856,
-59.9724845886231,11.9998178482056,
-77.8616333007813,-26.3757476806641,
-66.6003341674805,-39.0177764892578,
-18.7782039642334,-14.4839382171631,
31.8927688598633,18.4096641540527,
34.6711502075195,25.3995780944824,
-12.7085113525391,6.10976314544678,
-46.6345329284668,-4.09353590011597,
-18.2396392822266,9.75980186462402,
36.5433082580566,19.1664581298828,
42.7875862121582,-6.90049743652344,
-2.70915794372559,-43.7475433349609,
-26.0593452453613,-50.3888778686523,
18.1002178192139,-24.3298721313477,
79.2885742187500,-3.35185456275940,
79.6181640625000,-7.07736682891846,
24.2722492218018,-19.5881977081299,
-13.5456037521362,-17.6920280456543,
-3.44648528099060,-9.26826286315918,
5.39658355712891,-6.61505031585693,
-20.9978275299072,-2.85474324226379,
-50.1591224670410,7.77683353424072,
-33.2482757568359,9.55548572540283,
14.1525001525879,-8.48293113708496,
40.8672180175781,-21.0730972290039,
36.3791236877441,4.03142023086548,
36.0592765808106,46.5881500244141,
50.7494812011719,49.4452400207520,
53.7972373962402,8.79588699340820,
30.7451915740967,-20.8953285217285,
11.2449855804443,1.17151272296906,
21.3508129119873,46.2551727294922,
34.6527748107910,58.3768119812012,
16.0223159790039,26.4593353271484,
-14.0097656250000,-14.8026437759399,
-15.3898639678955,-37.5568389892578,
8.15935897827148,-47.5201721191406,
18.2372970581055,-48.5640449523926,
3.49356794357300,-36.5666084289551,
-1.31156671047211,-21.5307064056397,
23.5313072204590,-19.0069160461426,
49.3706741333008,-16.4247283935547,
39.1632461547852,16.3874797821045,
7.76668691635132,71.5372238159180,
-7.01339578628540,97.0816726684570,
-6.97751855850220,69.7505722045898,
-17.8373165130615,29.7782363891602,
-37.3210029602051,23.3944606781006,
-33.6874961853027,35.3862075805664,
-5.81172704696655,16.6423168182373,
6.14079618453980,-36.8391265869141,
-18.5014343261719,-63.6366271972656,
-46.2681198120117,-32.5238914489746,
-36.5556488037109,17.4425468444824,
3.06137752532959,37.8073234558106,
29.5606079101563,27.6889247894287,
26.0690708160400,16.8841476440430,
21.8751335144043,9.50831127166748,
32.0575790405273,-2.51074337959290,
36.9496345520020,-9.03329849243164,
18.2999649047852,8.41402912139893,
-12.5687131881714,35.9190711975098,
-36.2720603942871,38.5872726440430,
-44.9684257507324,15.7722129821777,
-41.6117134094238,9.12109184265137,
-24.8449420928955,40.0549468994141,
-7.76127433776856,70.5588836669922,
-9.88647842407227,56.2483749389648,
-33.7182922363281,10.7803344726563,
-38.6245193481445,-17.2808952331543,
7.07381772994995,-14.5416946411133,
71.7785949707031,-3.75839996337891,
83.9356307983398,-1.95034217834473,
27.6970272064209,0.387300223112106,
-31.0900249481201,10.8894824981689,
-27.3470802307129,13.1059961318970,
20.1193618774414,-2.02062344551086,
41.1698722839356,-12.0484142303467,
10.1086788177490,2.45914649963379,
-35.4646186828613,20.8151760101318,
-49.9900131225586,11.5238780975342,
-38.7494468688965,-20.2164058685303,
-39.0186576843262,-32.7964668273926,
-59.8626937866211,-13.3548641204834,
-72.0549163818359,6.85889863967896,
-50.6545829772949,-1.04041361808777,
-8.68998432159424,-23.5122528076172,
16.3946475982666,-25.8483791351318,
4.80736446380615,-5.11068820953369,
-23.7786483764648,13.3473377227783,
-29.2503013610840,16.7951869964600,
5.37721014022827,20.9969253540039,
42.2680358886719,36.0468444824219,
35.0476264953613,42.4130401611328,
-12.3445816040039,18.0231876373291,
-47.8318786621094,-21.6021881103516,
-32.5897521972656,-42.0221672058106,
12.8908615112305,-33.4176139831543,
36.5162467956543,-22.5200691223145,
20.8879375457764,-33.1360702514648,
0.828069329261780,-55.7442131042481,
7.39007520675659,-53.1217308044434,
22.0418682098389,-11.5399284362793,
17.7539558410645,37.3976402282715,
-3.06371784210205,54.2913932800293,
-10.9666442871094,33.8499603271484,
3.79618406295776,4.38874340057373,
22.7788658142090,-0.168696522712708,
26.9300689697266,18.4328575134277,
22.0983505249023,25.7470798492432,
17.6610145568848,-0.623412847518921,
10.4552097320557,-34.5290985107422,
-0.389364600181580,-36.4733276367188,
-0.389422059059143,-8.41091060638428,
19.7299499511719,4.29502916336060,
36.3206481933594,-20.9123516082764,
17.7348175048828,-46.2320785522461,
-20.7351913452148,-21.8719902038574,
-36.6869087219238,35.7524299621582,
-18.9723434448242,52.6473350524902,
-4.20717620849609,6.63262033462524,
-20.9569454193115,-44.9871597290039,
-48.9434852600098,-44.7340164184570,
-48.0463066101074,-18.0068874359131,
-17.9836997985840,-25.4503860473633,
8.95000839233398,-63.6091270446777,
25.2863903045654,-70.1925277709961,
47.5144577026367,-21.8407955169678,
62.4908981323242,33.7033576965332,
36.3617935180664,45.8629112243652,
-19.8650627136230,28.1215000152588,
-42.9211120605469,17.5584259033203,
-1.63500988483429,16.1355915069580,
47.7050819396973,-1.75119829177856,
35.9254150390625,-29.5810413360596,
-15.0058393478394,-42.0383987426758,
-24.9974002838135,-43.3462638854981,
20.4676742553711,-54.9408378601074,
48.2215881347656,-65.9181594848633,
10.5539379119873,-49.6414031982422,
-41.1423606872559,-16.7276306152344,
-36.8021011352539,-11.1355361938477,
-1.64526724815369,-42.9263229370117,
-2.82864189147949,-60.0189094543457,
-41.2579231262207,-29.1957969665527,
-50.8522567749023,17.9181938171387,
-0.884625911712647,24.5103969573975,
47.2686767578125,4.92385578155518,
36.8102302551270,15.4952268600464,
-9.20580673217773,52.1077308654785,
-23.1793022155762,55.3059806823731,
10.7426319122314,4.42354249954224,
48.8973350524902,-42.0214805603027,
57.0102577209473,-31.2364063262939,
42.6553153991699,17.2595233917236,
13.0332288742065,44.8507843017578,
-29.4742317199707,33.4914245605469,
-62.1875991821289,1.14007580280304,
-53.9308815002441,-33.1822814941406,
-8.83262443542481,-66.2444534301758,
26.1803379058838,-75.7539520263672,
17.9717292785645,-37.5379791259766,
-15.6526317596436,22.5196876525879,
-35.3268394470215,39.4509735107422,
-33.6898078918457,0.706225156784058,
-34.8189239501953,-34.5470962524414,
-39.5421066284180,-23.9116115570068,
-30.1843509674072,4.17717361450195,
-17.5067558288574,5.56285762786865,
-27.9963912963867,-10.6213569641113,
-53.2295913696289,-7.34329986572266,
-56.1572380065918,7.34806680679321,
-24.4668483734131,-8.33834171295166,
9.38949775695801,-52.9505691528320,
21.3748416900635,-60.4683189392090,
31.4182052612305,-8.33587646484375,
54.3000717163086,40.5517158508301,
68.3085174560547,27.3820705413818,
43.2163658142090,-24.5669593811035,
3.12869811058044,-45.6376495361328,
2.63679742813110,-30.6564884185791,
36.9042816162109,-25.0607547760010,
45.7640419006348,-38.4540176391602,
8.94447040557861,-27.4163532257080,
-25.4469032287598,24.0369625091553,
-11.1832342147827,65.4049682617188,
24.0727787017822,50.9043350219727,
28.3289661407471,18.2575263977051,
2.29613232612610,30.2506694793701,
-16.4557743072510,77.4657135009766,
-17.9255065917969,87.4246063232422,
-29.3100070953369,30.0975074768066,
-51.6305427551270,-38.6505928039551,
-44.5123977661133,-62.7221679687500,
6.97945404052734,-45.4694595336914,
55.0374679565430,-25.6552715301514,
45.8836631774902,-19.6624622344971,
-0.562799215316773,-11.4520978927612,
-22.6841449737549,4.70209693908691,
1.48606407642365,13.7168245315552,
35.2631301879883,10.9078931808472,
38.6256294250488,10.3933992385864,
11.6135139465332,23.7218227386475,
-14.9775190353394,37.4111442565918,
-20.3676776885986,38.5547103881836,
-9.99380111694336,29.0536079406738,
2.06566882133484,10.0099773406982,
1.49273788928986,-17.5098114013672,
-15.0579347610474,-41.0689582824707,
-30.7864398956299,-45.1754722595215,
-25.8067798614502,-21.2286968231201,
-2.24053931236267,15.9298877716064,
8.78883552551270,39.0510902404785,
-7.05752134323120,44.7319221496582,
-22.4732627868652,42.0918159484863,
-5.64369535446167,37.1938133239746,
33.5669250488281,28.8365192413330,
49.6086807250977,23.2325706481934,
22.6969833374023,31.8436527252197,
-14.3214006423950,48.8264656066895,
-14.2518959045410,46.2891540527344,
22.9144439697266,14.1479187011719,
55.0207901000977,-22.0538196563721,
48.6079139709473,-25.5173110961914,
16.5897140502930,7.93328189849854,
-8.86637783050537,37.8914833068848,
-12.1432037353516,26.8755130767822,
-5.52287435531616,-17.5531558990479,
-7.58475112915039,-48.9234733581543,
-21.0215091705322,-40.3412055969238,
-25.0789146423340,-6.36039495468140,
-4.72788047790527,17.0147972106934,
24.2867202758789,5.75860214233398,
29.2519760131836,-23.1515903472900,
1.69054388999939,-33.4951858520508,
-25.9393081665039,-2.15049433708191,
-20.4982795715332,51.0785293579102,
8.06002712249756,80.9691162109375,
10.7480077743530,58.6652717590332,
-32.1821975708008,9.31013107299805,
-72.1590576171875,-16.0559501647949,
-57.0408706665039,-0.176687955856323,
-5.07188034057617,17.9280815124512,
22.3509197235107,-4.53319072723389,
-1.46831357479095,-46.4761238098145,
-33.2249565124512,-50.5988540649414,
-26.8226871490479,-6.03899192810059,
6.45144462585449,38.7861938476563,
23.0564746856689,36.0747833251953,
14.3347845077515,7.92249107360840,
7.13282728195190,6.46039867401123,
8.60648250579834,42.1007766723633,
0.631256818771362,70.1253967285156,
-16.5718574523926,59.9651107788086,
-9.15164375305176,27.9738426208496,
31.2916164398193,5.54693078994751,
58.0419082641602,1.75749063491821,
30.8808040618897,6.79557180404663,
-24.4161148071289,15.7535943984985,
-45.3108634948731,18.9736347198486,
-21.2855930328369,1.32272875308990,
1.44431757926941,-31.3702259063721,
-6.35321903228760,-52.8208351135254,
-14.9619369506836,-49.4876518249512,
4.55787515640259,-40.3241882324219,
30.1987857818604,-50.8375091552734,
28.8803272247314,-68.6890258789063,
15.0902433395386,-57.4165687561035,
18.6357192993164,-16.9694442749023,
29.5601882934570,12.9966106414795,
13.0903587341309,12.0987644195557,
-22.9671058654785,7.86500072479248,
-27.6449470520020,17.2378711700439,
17.0819911956787,25.3288688659668,
54.6928367614746,13.8698749542236,
34.7395324707031,2.77040052413940,
-14.1924610137939,14.3528108596802,
-25.8575439453125,33.2654266357422,
8.79946517944336,27.6462955474854,
37.6842269897461,-0.218456983566284,
32.3523521423340,-12.6272830963135,
21.7971458435059,0.300528407096863,
27.2229881286621,2.59613204002380,
31.6078624725342,-17.5246505737305,
12.5904655456543,-24.4370975494385,
-13.1935396194458,12.3778190612793,
-18.5943145751953,54.9877014160156,
-16.7431545257568,58.2841033935547,
-37.8057250976563,28.0065574645996,
-74.6382293701172,3.67202615737915,
-79.9952087402344,-6.37832069396973,
-32.9694519042969,-26.6251525878906,
26.9715213775635,-51.8110046386719,
56.2489547729492,-36.0513687133789,
52.0141792297363,28.9770393371582,
25.7513389587402,79.7071151733398,
-14.9306907653809,59.1669807434082,
-58.1664352416992,-0.789803028106690,
-81.0293884277344,-27.6987342834473,
-68.9219055175781,-16.7213039398193,
-37.6636886596680,-22.9048080444336,
-12.3107509613037,-66.7657470703125,
6.40057945251465,-92.1058959960938,
33.5719833374023,-54.1214332580566,
60.5730552673340,15.2924947738647,
63.4079475402832,50.3645896911621,
48.3148422241211,36.5597839355469,
44.6361732482910,20.6753864288330,
53.2301864624023,30.2173023223877,
34.5366821289063,43.8148002624512,
-17.1528854370117,37.2006225585938,
-57.3400077819824,17.9838371276855,
-44.1170272827148,5.85487318038940,
-2.16298627853394,-6.35830211639404,
8.02789306640625,-22.5888462066650,
-19.6295127868652,-38.4594078063965,
-36.0298843383789,-46.4772033691406,
-11.9039869308472,-48.9434776306152,
13.9875631332397,-49.5532112121582,
9.74713802337647,-40.0559883117676,
-5.16381454467773,-15.8372364044189,
2.22897100448608,12.7313480377197,
17.2413196563721,20.0704154968262,
1.49217176437378,8.69526672363281,
-29.1932334899902,-1.76155567169189,
-23.9343414306641,-4.52766799926758,
29.2582073211670,-7.14909410476685,
68.7577743530273,-2.11597800254822,
47.4241905212402,27.5615119934082,
-5.19476652145386,64.6224136352539,
-23.1207141876221,68.6316375732422,
-0.260331481695175,31.4418678283691,
7.13270521163940,-4.09049320220947,
-24.6713905334473,-0.686589241027832,
-57.6891136169434,23.0866088867188,
-55.1633949279785,15.5981788635254,
-25.4929389953613,-26.8951110839844,
0.876776278018951,-62.5944557189941,
13.9672079086304,-68.0360565185547,
25.5463714599609,-62.9353981018066,
31.7383937835693,-58.0422897338867,
20.9146709442139,-31.5690078735352,
0.0608549416065216,12.7403640747070,
-12.5237522125244,32.6356315612793,
-19.4843025207520,2.23178148269653,
-34.4914588928223,-32.3141670227051,
-45.0357589721680,-12.3704462051392,
-20.6824893951416,41.5247306823731,
25.5835342407227,50.9718284606934,
38.5944747924805,-4.11014938354492,
-1.08362674713135,-54.0061607360840,
-42.4216766357422,-36.0073394775391,
-24.7942657470703,15.9668369293213,
37.2748222351074,29.4884433746338,
73.1015548706055,4.83303928375244,
50.1865997314453,3.93575906753540,
5.30128955841064,47.7889556884766,
-14.9152307510376,83.8905105590820,
-11.5599088668823,57.6567115783691,
-13.4874181747437,-6.63132619857788,
-23.7276210784912,-48.0404701232910,
-25.7094306945801,-40.2908248901367,
-12.8853254318237,-12.0106582641602,
4.87560939788818,5.04032611846924,
16.6675662994385,6.75900411605835,
23.0533771514893,2.26166486740112,
27.8431968688965,-6.51039743423462,
36.2218360900879,-17.8304691314697,
46.9226913452148,-13.4455881118774,
48.8123130798340,9.99948215484619,
30.6441268920898,34.3022651672363,
-3.49228429794312,37.5160026550293,
-28.2178249359131,16.4434318542480,
-17.6012058258057,-9.35420608520508,
15.4452028274536,-25.6429805755615,
38.6033782958984,-37.4312744140625,
37.0789222717285,-53.6225700378418,
25.5605545043945,-58.7376136779785,
20.4012966156006,-35.1236534118652,
16.5525398254395,8.33245658874512,
5.80274534225464,37.7119789123535,
-4.88457059860230,24.3935241699219,
-2.27677011489868,-21.4162788391113,
9.90719318389893,-57.3590011596680,
16.5220947265625,-52.1993446350098,
10.6052703857422,-12.1342649459839,
4.55041265487671,24.8551902770996,
6.17647171020508,31.8287277221680,
14.1866731643677,10.8763751983643,
21.5873680114746,-11.1580514907837,
26.8166790008545,-12.8230171203613,
23.3428573608398,-0.132246613502502,
-0.348793745040894,3.69073891639709,
-42.1018562316895,-7.14348793029785,
-73.0830230712891,-16.6198844909668,
-70.5997772216797,-10.7893342971802,
-40.9144477844238,-3.04163074493408,
-12.5168418884277,-9.09799194335938,
0.510133981704712,-24.7415275573730,
10.8282756805420,-29.1230049133301,
30.5231914520264,-18.0765266418457,
46.8106765747070,-16.1508369445801,
40.6545104980469,-36.7262878417969,
21.9597244262695,-55.3046646118164,
13.7819433212280,-49.8619537353516,
19.1330642700195,-30.8846836090088,
25.0766696929932,-26.0574398040772,
27.6246051788330,-32.0242195129395,
33.9709205627441,-21.9642410278320,
40.2135963439941,5.95802164077759,
30.1266956329346,18.5006275177002,
4.30185985565186,-1.61071681976318,
-4.02033615112305,-27.7635345458984,
19.9917831420898,-29.6674194335938,
43.4079208374023,-12.6159114837646,
24.4249973297119,-6.97219467163086,
-12.4492568969727,-15.0567770004272,
-10.0987796783447,-12.3829860687256,
36.1460151672363,9.21539306640625,
61.8293228149414,25.0369243621826,
22.4420948028564,19.0514411926270,
-33.0329399108887,3.57640910148621,
-38.0016021728516,-4.50117826461792,
-1.22501957416534,2.12536454200745,
3.65506434440613,16.7922534942627,
-44.3813056945801,28.0153026580811,
-78.5299758911133,20.2593460083008,
-45.1353874206543,-11.0275411605835,
19.9317321777344,-40.6813240051270,
44.0265083312988,-32.9127960205078,
24.0281238555908,13.7507152557373,
15.3199739456177,49.8677253723145,
41.4250831604004,34.5757980346680,
61.1770782470703,-3.36006069183350,
38.7215881347656,-7.47924995422363,
-9.52417755126953,21.4168376922607,
-44.1143798828125,29.0955162048340,
-57.6768722534180,-6.94050407409668,
-67.7417068481445,-41.4585113525391,
-71.8571319580078,-31.2820415496826,
-54.2610359191895,5.20492839813232,
-22.0079021453857,22.8988113403320,
-1.58229327201843,16.3132266998291,
1.84428620338440,18.9102878570557,
9.26719856262207,33.9497718811035,
23.2303867340088,32.8718986511231,
27.5031261444092,5.59599399566650,
10.4846143722534,-14.3418445587158,
-12.8167448043823,-4.59782743453980,
-23.4605197906494,10.7447032928467,
-26.1221370697022,0.346028864383698,
-33.2350120544434,-21.3656406402588,
-32.7458801269531,-25.1684703826904,
-3.76593375205994,-13.3256540298462,
37.6294059753418,-12.2363328933716,
57.0986824035645,-22.0164489746094,
46.2085380554199,-15.8642807006836,
27.4125499725342,16.9863548278809,
13.8667840957642,48.7907066345215,
-2.51262855529785,51.2062988281250,
-28.9469413757324,39.4931869506836,
-44.5810699462891,41.6184654235840,
-34.9111747741699,56.4163475036621,
-18.8875408172607,59.9431076049805,
-19.4639492034912,45.8914718627930,
-25.0507545471191,26.1674365997314,
-3.04429316520691,12.6455173492432,
41.1407127380371,2.59201121330261,
56.6110229492188,-5.92638683319092,
18.7892742156982,-10.8203420639038,
-34.5624923706055,-13.1547870635986,
-48.7970733642578,-19.5911369323730,
-20.9991607666016,-23.2354640960693,
1.91185402870178,-8.37633705139160,
-13.0848884582520,25.6438064575195,
-46.7975349426270,47.4662208557129,
-60.6137924194336,29.3752403259277,
-41.3196067810059,-8.51119327545166,
-7.35450172424316,-24.2499389648438,
15.8712072372437,2.59044647216797,
19.0200710296631,43.2331771850586,
0.979137957096100,61.0345687866211,
-28.9270324707031,47.9786758422852,
-53.0449523925781,23.2464866638184,
-58.8155136108398,3.47023701667786,
-52.6910934448242,-9.01958370208740,
-48.5661239624023,-22.5495433807373,
-48.8203735351563,-38.4102668762207,
-40.6648254394531,-52.5303535461426,
-16.2084732055664,-60.2901115417481,
14.0223951339722,-51.2084617614746,
29.1780090332031,-23.8556632995605,
20.6838264465332,11.9037876129150,
0.348346590995789,40.8974380493164,
-19.9481544494629,51.5171546936035,
-26.2000579833984,36.8785476684570,
-14.3121376037598,-2.79850244522095,
10.9288940429688,-47.9244155883789,
28.2323360443115,-63.8928070068359,
21.0968608856201,-31.5126228332520,
-2.79257082939148,25.5354690551758,
-14.0932579040527,51.2610244750977,
2.05576086044312,21.5692138671875,
34.4519309997559,-20.5511703491211,
52.3353080749512,-15.6935348510742,
44.3031349182129,34.5908851623535,
14.8899288177490,68.4781723022461,
-18.9731082916260,44.2010650634766,
-47.0645599365234,-12.2082958221436,
-55.2801055908203,-43.1122131347656,
-43.9382514953613,-34.7804069519043,
-33.0715904235840,-17.7227401733398,
-36.6770248413086,-14.2967052459717,
-48.9233703613281,-10.4074916839600,
-48.4887390136719,2.60952520370483,
-36.3669967651367,1.85289049148560,
-27.3999958038330,-24.1409339904785,
-21.4176311492920,-51.4941177368164,
-0.585846185684204,-44.8186721801758,
39.2381706237793,-14.5495910644531,
65.0164566040039,-3.31001591682434,
51.7278099060059,-18.0410003662109,
25.5787963867188,-27.6001815795898,
35.6271286010742,-13.7115545272827,
72.3342056274414,0.836102128028870,
77.3656463623047,-8.55026245117188,
26.7056045532227,-26.3169059753418,
-35.9748077392578,-20.0588264465332,
-59.2929573059082,-0.104378342628479,
-52.4154548645020,-1.82804656028748,
-51.8502197265625,-29.1403045654297,
-55.1419906616211,-50.9629287719727,
-31.1117172241211,-46.5234375000000,
18.3843784332275,-26.9801025390625,
45.7408256530762,-5.01716184616089,
37.3169059753418,21.0435543060303,
32.2867813110352,40.7084350585938,
53.1736831665039,34.5735664367676,
65.4595336914063,5.31731891632080,
34.9034271240234,-12.0468063354492,
-4.54027652740479,9.60884380340576,
0.788794577121735,39.6415290832520,
41.2034530639648,29.1012935638428,
50.7428512573242,-14.9940338134766,
12.6405591964722,-43.1986274719238,
-17.6879673004150,-29.2143669128418,
3.97666501998901,3.20126175880432,
32.0112724304199,25.9853935241699,
10.4681358337402,30.5157985687256,
-41.4413490295410,17.1980972290039,
-49.2062110900879,-9.22116947174072,
0.879863262176514,-28.6577529907227,
40.5360908508301,-10.8099784851074,
23.8985843658447,35.3092155456543,
-16.5797863006592,48.7063293457031,
-23.3438816070557,-7.54086637496948,
1.49070250988007,-81.5291366577148,
14.5802755355835,-86.6487274169922,
-1.13271141052246,-16.3085498809814,
-15.2975959777832,47.2064704895020,
-6.42094087600708,43.5536117553711,
1.62779438495636,10.3650598526001,
-18.4899253845215,7.89401197433472,
-53.2427864074707,34.6731109619141,
-68.3500366210938,39.7621421813965,
-47.4576416015625,9.60047435760498,
-2.31239080429077,-11.2025165557861,
38.1778640747070,4.10758638381958,
46.8282318115234,24.5496330261230,
24.6430168151855,12.5695896148682,
-2.68565750122070,-19.5645217895508,
-13.3356027603149,-36.4997749328613,
-6.24892711639404,-34.5649032592773,
0.0532192364335060,-42.6340560913086,
-1.11188650131226,-62.5691795349121,
8.21732234954834,-66.3894271850586,
33.9671897888184,-47.4345817565918,
48.8003730773926,-32.9167175292969,
30.2625694274902,-43.9851417541504,
0.129999458789825,-60.6687164306641,
-5.62648153305054,-46.9563903808594,
7.16081237792969,-10.8211469650269,
0.289384722709656,10.4607696533203,
-30.3211917877197,1.97420799732208,
-38.9303283691406,-8.88472747802734,
1.76149368286133,3.26417970657349,
52.6193084716797,31.2439422607422,
54.7946662902832,49.8641357421875,
9.38755226135254,45.3524360656738,
-24.9762096405029,20.1606025695801,
-13.7857637405396,-16.9394321441650,
15.4370660781860,-53.0017814636231,
23.2705669403076,-68.6767272949219,
7.94768762588501,-54.9258270263672,
-4.57351779937744,-24.4650688171387,
-5.57211112976074,-9.25860595703125,
-3.03958916664124,-18.4875831604004,
2.95480060577393,-36.6510887145996,
17.5206851959229,-44.0130195617676,
28.2551269531250,-39.7980690002441,
13.2613363265991,-29.8811511993408,
-25.2723693847656,-19.2867374420166,
-52.4071578979492,-13.2836542129517,
-36.5386314392090,-11.0929698944092,
4.55016756057739,-3.87232542037964,
23.8944149017334,16.2293872833252,
5.61026573181152,42.0652236938477,
-30.2937412261963,43.2267417907715,
-53.1755065917969,8.33272933959961,
-49.2570037841797,-35.1222000122070,
-23.3591823577881,-46.3085517883301,
8.16886138916016,-20.3923835754395,
29.6471405029297,4.64866304397583,
32.9742965698242,7.71449232101440,
25.8784465789795,0.903267085552216,
25.3911495208740,0.0806511640548706,
29.5994167327881,-4.22351837158203,
16.6110477447510,-22.8067493438721,
-15.5656118392944,-39.9173202514648,
-35.6797790527344,-29.1694717407227,
-12.5364913940430,4.62649917602539,
29.5560092926025,28.1086082458496,
46.2491035461426,28.9368724822998,
27.9321651458740,27.0781040191650,
11.6780757904053,37.9344406127930,
24.6098918914795,42.9531364440918,
43.7141914367676,24.9172325134277,
36.7528839111328,3.10928845405579,
14.2937641143799,4.53357505798340,
9.36308956146240,21.7363033294678,
26.2505607604980,24.4951343536377,
32.7202453613281,3.78086376190186,
10.3076343536377,-12.7473983764648,
-21.5643272399902,-6.30274868011475,
-38.5970535278320,6.94161558151245,
-42.3605499267578,5.58166551589966,
-50.1826820373535,-5.62981081008911,
-59.3786735534668,-10.7195177078247,
-54.0818023681641,-16.0834407806397,
-28.1774482727051,-39.1070861816406,
9.76571846008301,-65.7469940185547,
40.2878150939941,-57.3768997192383,
51.0944175720215,-6.06533765792847,
38.4622230529785,41.9459762573242,
9.89087295532227,39.3311691284180,
-20.5920333862305,-5.79913711547852,
-29.7553558349609,-36.1627922058106,
-12.4386978149414,-18.2416667938232,
16.7902851104736,20.1407146453857,
34.7650947570801,30.4144363403320,
25.3874359130859,9.50394821166992,
-9.57015037536621,-10.7938070297241,
-43.0014266967773,-3.67543697357178,
-39.0091667175293,22.5602741241455,
5.31334209442139,34.4600219726563,
48.5766677856445,15.1632385253906,
44.2157630920410,-20.9150524139404,
-2.28137207031250,-42.3943367004395,
-27.4356613159180,-32.1860847473145,
9.97080039978027,-5.06701660156250,
70.3516387939453,11.7407608032227,
76.9999542236328,8.03084659576416,
12.6744003295898,3.74225640296936,
-53.7336235046387,16.3487758636475,
-57.4215812683106,24.3073005676270,
-12.6066331863403,-6.85084009170532,
18.4538021087647,-64.5847015380859,
12.0333080291748,-87.9203796386719,
2.28915500640869,-43.1248168945313,
20.2045459747314,30.5936298370361,
45.5564651489258,65.4214019775391,
41.9232788085938,44.4302330017090,
12.5309638977051,15.5209159851074,
-14.6320428848267,18.8100051879883,
-25.8347129821777,36.6571998596191,
-32.3029212951660,33.5072937011719,
-34.1658859252930,2.87668895721436,
-19.2754116058350,-23.3508987426758,
9.91881179809570,-20.9666347503662,
21.8730792999268,5.01617813110352,
5.39028835296631,31.5448169708252,
-18.4125862121582,34.1944274902344,
-22.7773666381836,4.96331071853638,
-9.91911506652832,-34.7320213317871,
-6.29602718353272,-44.3439369201660,
-8.83185291290283,-9.81022167205811,
7.48494338989258,34.2937355041504,
39.7300796508789,42.1620254516602,
53.9822998046875,5.13350915908814,
31.7883033752441,-40.9826202392578,
2.01764678955078,-59.2303390502930,
3.91671395301819,-49.9975547790527,
36.4711608886719,-33.2750930786133,
61.6017532348633,-15.2412776947021,
61.3174667358398,0.548370480537415,
45.0355453491211,6.82483959197998,
23.5489711761475,-2.48591279983521,
-7.25337886810303,-18.7438507080078,
-36.2911224365234,-29.2699241638184,
-32.6279449462891,-35.4683227539063,
8.40159606933594,-44.0301437377930,
41.3519859313965,-48.5094261169434,
21.5736846923828,-40.4320297241211,
-30.0806941986084,-27.0846004486084,
-47.1177024841309,-19.9084930419922,
-6.08628749847412,-18.5081844329834,
38.3891410827637,-8.08831977844238,
30.4111766815186,16.5662708282471,
-16.7707366943359,35.5884475708008,
-45.8928680419922,38.3172187805176,
-35.3773345947266,36.1463737487793,
-21.2741260528564,36.3780937194824,
-26.7459297180176,25.1462993621826,
-33.9105148315430,-5.24766635894775,
-17.7048206329346,-33.2415733337402,
7.19654226303101,-35.5731239318848,
8.50350189208984,-20.1190567016602,
-12.5830669403076,-15.7364425659180,
-25.3509941101074,-24.3745956420898,
-14.3292274475098,-14.9754390716553,
0.514220714569092,18.7420196533203,
-6.94421768188477,39.6422615051270,
-28.4791164398193,18.6676921844482,
-33.3996620178223,-16.5106105804443,
-11.1423168182373,-13.6927347183228,
21.9849338531494,29.7060031890869,
41.6366310119629,55.6240463256836,
36.4874191284180,31.2078876495361,
13.6481208801270,-11.0503225326538,
-11.9237375259399,-11.3857707977295,
-26.6042346954346,33.7458000183106,
-25.1770458221436,67.4156494140625,
-9.95549774169922,50.7280731201172,
6.01559782028198,9.78334236145020,
5.63596057891846,-6.37566518783569,
-15.9882469177246,5.73080348968506,
-37.1436347961426,9.79423046112061,
-31.4394454956055,-17.8175563812256,
-0.477912873029709,-50.7866935729981,
23.8434963226318,-53.5594367980957,
18.0425796508789,-25.4033641815186,
0.151073932647705,13.3245334625244,
8.50581359863281,46.7709770202637,
36.7189559936523,64.4672927856445,
44.4551811218262,50.2010269165039,
16.0611972808838,-0.519849300384522,
-6.15652465820313,-49.5639762878418,
7.52723550796509,-46.4392089843750,
25.5948009490967,1.89837074279785,
5.69241476058960,31.4772472381592,
-35.4770393371582,9.44884204864502,
-37.7015113830566,-27.2906303405762,
5.34035015106201,-21.6321964263916,
29.7348308563232,18.7332725524902,
-7.79625606536865,36.1412467956543,
-53.3804092407227,8.89028263092041,
-35.3624000549316,-21.6009826660156,
30.2955894470215,-20.6414394378662,
64.4086685180664,-4.74337720870972,
39.6169738769531,-1.35520637035370,
14.9673604965210,-12.5718364715576,
32.2043876647949,-23.9501438140869,
52.8399620056152,-28.1661891937256,
27.3423213958740,-22.2295532226563,
-22.8188877105713,1.43298995494843,
-37.0916519165039,33.6299934387207,
-17.6452770233154,47.4856681823731,
-22.9733409881592,24.5546894073486,
-68.6812744140625,-11.3271570205688,
-90.6748962402344,-25.2522869110107,
-42.7756767272949,-22.7277336120605,
26.0753631591797,-35.3232841491699,
38.1446189880371,-60.8486671447754,
-5.42176723480225,-58.4236984252930,
-38.7850875854492,-18.3322544097900,
-30.2401409149170,16.7018966674805,
-14.8854198455811,11.6358528137207,
-21.5009117126465,-12.9087810516357,
-27.1272583007813,-20.1500320434570,
1.70301163196564,-7.77182722091675,
40.8479881286621,-5.58679676055908,
43.0957527160645,-22.7145919799805,
15.7374000549316,-40.4654388427734,
8.21331977844238,-39.3204231262207,
32.3885498046875,-20.8843517303467,
48.1356391906738,3.11672139167786,
23.7652130126953,28.9113292694092,
-17.5027046203613,41.1475143432617,
-41.1924934387207,26.7853832244873,
-40.7354698181152,3.94552969932556,
-38.4519042968750,2.18458271026611,
-40.0817718505859,15.8507308959961,
-33.1750946044922,4.22953891754150,
-23.9796581268311,-38.5207557678223,
-30.2589702606201,-66.6239395141602,
-40.2944107055664,-46.0223007202148,
-29.0185146331787,-10.1866989135742,
-0.364120483398438,-14.9586114883423,
11.4103116989136,-48.3068504333496,
-3.16346788406372,-44.0872840881348,
-15.6901378631592,16.6717624664307,
-2.92537927627563,69.2133255004883,
8.62941741943359,58.9997711181641,
-12.2660551071167,15.0463743209839,
-52.1148033142090,-3.53849005699158,
-66.1078262329102,5.98088884353638,
-48.2729110717773,-1.16239202022553,
-37.3072891235352,-31.9582672119141,
-46.7530822753906,-43.7487487792969,
-43.7056922912598,-15.7906188964844,
-5.23197555541992,16.1687240600586,
38.3142852783203,12.6477851867676,
42.3049201965332,-12.3399772644043,
13.0360298156738,-19.9749641418457,
-4.26755189895630,-3.32894539833069,
10.2542734146118,5.88873481750488,
33.7328948974609,-0.821642458438873,
42.6125602722168,-0.218752086162567,
38.1405525207520,19.4480075836182,
29.9022712707520,35.3822402954102,
13.6164999008179,25.7839298248291,
-6.10197210311890,-1.96948027610779,
-3.58373069763184,-16.7101917266846,
37.8246498107910,-3.36101412773132,
81.0752334594727,24.2856426239014,
73.8308944702148,41.5008392333984,
7.71494245529175,36.7440948486328,
-61.9825820922852,19.3376865386963,
-78.5676574707031,4.30507040023804,
-43.5674362182617,4.69626569747925,
-6.50472164154053,22.1277198791504,
-6.20251417160034,39.2556953430176,
-28.9255237579346,42.6298637390137,
-42.4339599609375,34.9616584777832,
-34.3760833740234,22.5708103179932,
-18.7274761199951,7.67981195449829,
-16.0518608093262,-4.71949672698975,
-26.7865295410156,-6.32434225082398,
-38.3420028686523,4.42464733123779,
-37.2752037048340,14.3171138763428,
-27.9496650695801,0.952993631362915,
-24.2497730255127,-28.5502738952637,
-31.1146430969238,-37.0746879577637,
-35.2475814819336,-7.42214632034302,
-31.1440925598145,25.1304931640625,
-23.7118053436279,10.8184814453125,
-24.4191036224365,-42.9871101379395,
-34.4085922241211,-70.4214172363281,
-35.4646110534668,-32.7574424743652,
-21.7120056152344,26.7318477630615,
-7.05841493606567,34.7546463012695,
-0.0380263924598694,-16.4672145843506,
7.06289720535278,-57.7254753112793,
24.4707164764404,-34.2152290344238,
34.6899566650391,28.1021862030029,
24.7193889617920,64.3175506591797,
7.67036628723145,47.9385528564453,
9.47350311279297,0.590498328208923,
23.7683448791504,-45.1473350524902,
18.1843757629395,-71.8024673461914,
-15.2556724548340,-65.4919586181641,
-33.4662704467773,-26.2738628387451,
-6.76422405242920,17.1451377868652,
32.0065956115723,23.5329494476318,
28.4333820343018,-5.36968708038330,
-11.7185850143433,-21.0157852172852,
-35.9546470642090,3.22366762161255,
-25.5183582305908,34.3174743652344,
-24.4379787445068,25.2939720153809,
-59.0633888244629,-10.5197706222534,
-89.5716552734375,-21.3070850372314,
-62.6943855285645,7.03842926025391,
3.77678728103638,34.9679718017578,
37.3244552612305,35.5294456481934,
7.37454843521118,29.4032039642334,
-40.9202880859375,40.8967628479004,
-56.8889007568359,47.8716964721680,
-41.4932594299316,13.3160114288330,
-28.5352859497070,-42.9142494201660,
-26.2909297943115,-64.4408264160156,
-17.2314071655273,-26.7248744964600,
-0.886649191379547,21.9737777709961,
7.20750617980957,27.1014556884766,
7.97682666778564,-4.66806840896606,
15.1306934356689,-22.2770996093750,
30.1852283477783,-0.107887744903564,
30.9195671081543,38.4994621276856,
0.428954601287842,53.6897392272949,
-40.8399238586426,28.2760601043701,
-51.4422988891602,-13.6131744384766,
-17.5458431243897,-38.8057746887207,
31.2117481231689,-38.6323661804199,
54.3388862609863,-26.2103557586670,
32.6312522888184,-23.0038719177246,
-19.7410678863525,-30.9801616668701,
-60.6371345520020,-32.3057708740234,
-64.0964584350586,-12.1103916168213,
-40.8509902954102,12.8642616271973,
-24.0312442779541,18.6475048065186,
-29.4138469696045,11.3675327301025,
-36.7051239013672,15.9932403564453,
-23.7382755279541,30.6902332305908,
3.21932601928711,25.1314964294434,
22.1865673065186,-16.2936115264893,
28.3922653198242,-54.5156860351563,
39.5032997131348,-36.5904273986816,
55.0071144104004,22.0397205352783,
41.4275779724121,51.1448402404785,
-9.20513820648193,19.7816772460938,
-55.7489242553711,-24.0661582946777,
-55.8482551574707,-16.9184818267822,
-16.2655143737793,29.1292037963867,
10.2394742965698,47.2753715515137,
-4.85752296447754,11.5238828659058,
-35.7954788208008,-29.5440216064453,
-51.7141609191895,-33.6884918212891,
-50.8877601623535,-18.4657154083252,
-42.9245033264160,-25.2967281341553,
-16.9980545043945,-51.7493515014648,
28.6522121429443,-52.8670845031738,
59.1889610290527,-12.9679355621338,
31.4722366333008,26.0516014099121,
-36.5184974670410,19.4795932769775,
-68.2102203369141,-22.4137420654297,
-20.2687873840332,-47.6068038940430,
51.9286613464356,-26.6270446777344,
64.8355484008789,17.8311252593994,
12.9865493774414,36.5893211364746,
-31.2160949707031,7.85192489624023,
-14.5719251632690,-38.3236732482910,
26.8439044952393,-58.0386276245117,
25.9377765655518,-40.2358055114746,
-18.2453479766846,-12.6933813095093,
-40.7468070983887,-5.60911989212036,
-9.59056377410889,-18.3914394378662,
33.8877410888672,-22.1664505004883,
32.8593406677246,-2.06724357604980,
-5.62690353393555,24.6530036926270,
-24.7066783905029,33.4732933044434,
1.59168338775635,26.0807247161865,
33.7239456176758,14.7450895309448,
18.6258239746094,4.67698383331299,
-25.1995639801025,-7.66752052307129,
-35.3498115539551,-23.8978939056397,
4.41165542602539,-33.7462387084961,
46.2147407531738,-30.6756896972656,
32.7820091247559,-22.8664321899414,
-20.7371921539307,-15.5865907669067,
-46.1836242675781,-0.605953454971314,
-15.6048431396484,25.6806697845459,
19.2676715850830,44.7211227416992,
4.01071548461914,30.8343944549561,
-39.6644477844238,-10.8735580444336,
-48.6609954833984,-38.3293418884277,
-8.01377487182617,-18.7265682220459,
24.5381603240967,24.1466197967529,
2.15969824790955,39.1871414184570,
-40.5397300720215,9.82987880706787,
-34.2009239196777,-22.8043708801270,
27.6274909973145,-18.7633342742920,
80.4863815307617,8.24895954132080,
73.0988388061523,16.1918048858643,
28.8754787445068,-0.623363375663757,
4.29856967926025,-4.58716821670532,
11.6962375640869,23.8277053833008,
13.9454965591431,58.8920440673828,
-15.9381999969482,61.4222488403320,
-60.2131423950195,31.9152927398682,
-81.1368179321289,3.18076729774475,
-61.2695999145508,-5.88344430923462,
-14.4423294067383,3.03383708000183,
26.3287868499756,19.5052375793457,
31.8412513732910,38.1075744628906,
4.37316942214966,46.2592964172363,
-24.9443817138672,32.2810478210449,
-19.8241882324219,7.27142858505249,
16.8323650360107,-0.588143944740295,
39.7483024597168,13.2919569015503,
16.2030010223389,20.2418212890625,
-27.6077213287354,-0.439264297485352,
-41.9049377441406,-30.7548065185547,
-10.3470792770386,-37.7393112182617,
31.5366878509522,-13.2493801116943,
44.4935760498047,16.2794857025147,
27.1855068206787,22.4197235107422,
4.49524974822998,7.56046056747437,
-7.15579700469971,-14.9894752502441,
-12.2143478393555,-33.6124763488770,
-6.71160125732422,-41.8980789184570,
14.5727424621582,-38.8340377807617,
39.6677474975586,-26.7382202148438,
43.9116592407227,-10.2375087738037,
18.3593959808350,11.4696350097656,
-13.1265687942505,34.2696723937988,
-22.9679107666016,38.2184257507324,
-11.8744211196899,9.17450046539307,
-1.38049697875977,-35.8973159790039,
0.415646344423294,-55.4875259399414,
1.21873486042023,-28.2784538269043,
3.01403379440308,17.9890880584717,
-4.53263759613037,36.2238388061523,
-19.1876335144043,15.7833595275879,
-17.2088966369629,-14.9943809509277,
10.5501852035522,-27.3441181182861,
34.9952583312988,-20.4027843475342,
22.9579086303711,-2.37846398353577,
-14.2752628326416,21.6842918395996,
-29.9605598449707,47.2933273315430,
-6.18220043182373,53.3570213317871,
19.4786357879639,32.0707855224609,
5.78962326049805,-2.02244400978088,
-35.3539848327637,-22.4255123138428,
-53.6797485351563,-18.6337547302246,
-27.9513359069824,-1.35931527614594,
13.0202903747559,11.5780124664307,
27.7057132720947,12.5051002502441,
7.84544563293457,-0.229715585708618,
-23.1893386840820,-25.7269935607910,
-37.8245353698731,-51.6184883117676,
-23.9742088317871,-59.0128593444824,
12.5264616012573,-46.8351936340332,
48.3996238708496,-26.7486820220947,
56.0024185180664,-4.13286876678467,
30.6283721923828,25.6186180114746,
-2.12182283401489,57.7931289672852,
-7.38402557373047,66.0594863891602,
14.3793907165527,32.7538719177246,
29.5177154541016,-12.0112161636353,
17.7869529724121,-22.6725463867188,
-6.74631977081299,13.1799802780151,
-19.0356521606445,53.4671478271484,
-15.6739740371704,51.6735458374023,
-11.3907995223999,14.6085290908813,
-13.4100027084351,-9.61779594421387,
-11.6328582763672,4.53905200958252,
0.103699445724487,33.4470787048340,
9.98170948028565,34.7713317871094,
7.78604030609131,0.614641666412354,
-4.57348442077637,-38.5232925415039,
-18.7944717407227,-42.4193267822266,
-29.8908519744873,-11.9273843765259,
-36.9158325195313,11.2577428817749,
-29.0683727264404,-6.39928865432739,
-5.54797220230103,-48.9342689514160,
22.7470207214355,-59.8829536437988,
40.0125160217285,-17.0495815277100,
42.5674705505371,39.0576744079590,
38.6297416687012,47.4531784057617,
29.8616771697998,0.0770401954650879,
8.18126296997070,-45.7633361816406,
-20.4260768890381,-44.2058639526367,
-32.5310134887695,-14.6860179901123,
-15.8879108428955,-2.19715523719788,
8.57468032836914,-13.0581245422363,
16.6739273071289,-13.4337759017944,
10.8964147567749,16.9048652648926,
6.28698253631592,55.7039489746094,
0.617741525173187,66.2753143310547,
-22.3622188568115,43.4866485595703,
-55.9014472961426,7.07795381546021,
-60.5046157836914,-22.0359477996826,
-21.5047950744629,-30.8115959167480,
26.4326438903809,-15.5217437744141,
35.2782325744629,8.72669029235840,
10.8633308410645,14.8677730560303,
-4.60055828094482,-11.4345560073853,
4.41567993164063,-41.9337081909180,
6.31452560424805,-40.0849037170410,
-14.5177936553955,-11.9799089431763,
-30.0708160400391,2.12073302268982,
-11.3981132507324,-18.7620124816895,
23.4517459869385,-48.8690948486328,
28.9201240539551,-50.1266708374023,
-4.46071910858154,-26.5776920318604,
-36.4275779724121,-11.5995645523071,
-32.9811820983887,-18.6599712371826,
0.173789262771606,-23.7556419372559,
34.3596420288086,-15.1311292648315,
50.7976646423340,-2.18111324310303,
52.8530769348145,1.11270868778229,
44.7509078979492,2.10937142372131,
37.0353088378906,13.2946395874023,
40.8334655761719,22.0527820587158,
51.6513519287109,11.9130191802979,
52.4310073852539,-4.35257673263550,
30.7261543273926,4.26229000091553,
-3.69423985481262,39.6074752807617,
-22.4036045074463,61.7807693481445,
-8.09877490997315,41.8314018249512,
26.2604694366455,7.18184852600098,
45.8613357543945,6.15263795852661,
27.8176746368408,38.9666557312012,
-17.6524791717529,55.9615402221680,
-51.5752220153809,24.7122421264648,
-38.5098571777344,-24.5059223175049,
9.75921821594238,-39.8940124511719,
44.3231620788574,-14.3316001892090,
32.1956748962402,15.0327224731445,
-10.0725975036621,21.4868736267090,
-32.3915519714356,18.9823513031006,
-17.9079380035400,25.3990230560303,
10.8130817413330,32.5104713439941,
29.0144367218018,23.5366363525391,
30.6610412597656,7.70392370223999,
29.0799274444580,11.4642314910889,
25.2433300018311,33.8171958923340,
10.3346481323242,50.6393775939941,
-9.03445720672607,40.7303276062012,
-17.8094520568848,15.0416898727417,
-10.1662445068359,-1.54013311862946,
4.90840911865234,-4.51429128646851,
16.8824920654297,-9.64130401611328,
20.6787967681885,-21.4246234893799,
11.8311929702759,-31.9054508209229,
-16.1077251434326,-33.3462333679199,
-49.6183090209961,-27.1161460876465,
-54.2004814147949,-19.6990642547607,
-11.2516908645630,-16.7398452758789,
51.5639305114746,-9.98204135894775,
82.9376373291016,11.0364780426025,
56.3583641052246,40.3657531738281,
0.193489551544189,55.6213264465332,
-43.6886024475098,35.0150032043457,
-58.3349037170410,-11.3830595016480,
-52.6147079467773,-44.9394035339356,
-34.3216781616211,-34.2612113952637,
-10.2270622253418,4.20948934555054,
7.15145587921143,34.5490608215332,
6.14899492263794,42.0756874084473,
-5.98817777633667,41.6807327270508,
-6.65503120422363,36.0230140686035,
9.74416732788086,7.98899555206299,
21.5261821746826,-40.3974876403809,
15.2095394134521,-69.6984176635742,
7.91581439971924,-43.0066223144531,
22.2823333740234,17.8806533813477,
44.2133903503418,54.1018447875977,
38.3640174865723,40.4442863464356,
5.25236129760742,8.93706989288330,
-14.6079711914063,1.15128898620605,
5.77735233306885,15.4654750823975,
40.4760665893555,26.5233078002930,
44.1693496704102,30.0334014892578,
10.8280315399170,39.7565460205078,
-24.4548397064209,50.7286071777344,
-30.4827251434326,46.4311523437500,
-11.7371902465820,27.0003166198730,
5.97016620635986,8.56509590148926,
7.66942453384399,3.90658998489380,
-7.87134742736816,5.34617137908936,
-32.9323196411133,2.97711586952209,
-52.1380844116211,1.38453948497772,
-51.8415756225586,-3.83898806571960,
-38.2408523559570,-27.0685825347900,
-25.8101158142090,-67.4479522705078,
-10.0357179641724,-82.6366195678711,
17.8264579772949,-46.7767219543457,
47.9497299194336,4.67299985885620,
53.7837028503418,14.1164045333862,
28.9932212829590,-15.1823549270630,
4.11340284347534,-25.2526016235352,
12.4093275070190,10.4433727264404,
39.2691574096680,38.5355453491211,
46.3756790161133,8.66067504882813,
32.1216278076172,-48.0433959960938,
24.4325294494629,-54.4274711608887,
27.1010150909424,-2.33800053596497,
12.8711690902710,40.5815353393555,
-18.2695083618164,32.1091690063477,
-25.8665180206299,7.66422653198242,
13.1631145477295,10.8822956085205,
53.2816848754883,27.0914154052734,
41.2648124694824,19.7688159942627,
-6.75039482116699,-1.90514862537384,
-22.2996063232422,-1.09926569461823,
10.2099819183350,22.0485324859619,
33.9965095520020,30.7201766967773,
9.41732978820801,11.5327548980713,
-24.1060791015625,-3.24601674079895,
-19.6706218719482,8.84199047088623,
3.31086254119873,20.9427509307861,
-10.4000701904297,0.367183446884155,
-52.1772308349609,-35.2851104736328,
-55.4603958129883,-44.0363273620606,
3.08009147644043,-21.2238082885742,
57.4747467041016,2.44191145896912,
43.5303192138672,3.67547607421875,
-8.79842948913574,-7.94591331481934,
-20.9028892517090,-10.4567794799805,
18.8019599914551,6.41225242614746,
42.4223442077637,28.1210002899170,
7.40024948120117,37.2257385253906,
-36.3390235900879,25.7325286865234,
-24.4261989593506,5.99952650070190,
33.3474388122559,-3.84887814521790,
65.9015045166016,2.44834184646606,
37.1550331115723,10.7052822113037,
-11.4413642883301,5.90763139724731,
-27.4543609619141,-3.19251680374146,
-8.90593528747559,-1.06839275360107,
11.5890083312988,6.05287313461304,
19.1023597717285,0.638836562633514,
19.6700000762939,-7.28247880935669,
13.7369260787964,9.88312721252441,
-4.13908100128174,51.6198616027832,
-20.2644004821777,80.8476257324219,
-22.9504795074463,72.9516983032227,
-22.6714363098145,47.9245452880859,
-38.4180564880371,38.3812141418457,
-60.4092521667481,37.5793838500977,
-55.5092811584473,15.5625181198120,
-8.66223526000977,-23.8157844543457,
43.2099151611328,-42.0056991577148,
56.8831176757813,-26.7455806732178,
42.8444747924805,-12.6224231719971,
33.6942481994629,-20.1258163452148,
38.4480667114258,-18.3622589111328,
36.6588668823242,15.8702278137207,
12.6816186904907,49.5544548034668,
-22.1865272521973,34.2010650634766,
-48.6247482299805,-17.6028633117676,
-51.2811431884766,-36.5283584594727,
-27.4017715454102,3.26144218444824,
4.62853813171387,42.2987861633301,
12.9041881561279,24.5826816558838,
-19.3770751953125,-21.7690715789795,
-58.1471862792969,-30.7466011047363,
-50.4528160095215,-2.83511495590210,
8.91438293457031,4.93156671524048,
56.5470314025879,-20.2839450836182,
48.2386093139648,-22.2871627807617,
14.2982940673828,27.1948280334473,
-4.21607828140259,70.9644622802734,
-13.8307008743286,44.7748603820801,
-39.9104537963867,-21.3519287109375,
-59.0393676757813,-44.1711044311523,
-28.4557533264160,-4.54818010330200,
34.7612686157227,28.9532833099365,
54.8768539428711,11.6258430480957,
1.77689647674561,-13.7591199874878,
-55.7517127990723,2.13799834251404,
-52.9658164978027,35.8341331481934,
-19.9349803924561,32.9965972900391,
-23.0956249237061,-1.42375493049622,
-51.1199684143066,-21.6306095123291,
-38.1099090576172,-7.93434333801270,
20.9237155914307,11.3588113784790,
51.0698165893555,16.0176162719727,
14.5135049819946,15.2419624328613,
-33.1605339050293,10.9238252639771,
-26.8866748809814,-15.0914964675903,
11.6815919876099,-59.3428611755371,
13.4821434020996,-72.0282211303711,
-25.0793399810791,-27.5115566253662,
-44.9706802368164,27.3476467132568,
-18.8200073242188,34.4153785705566,
8.24252986907959,-4.23667621612549,
-4.79234552383423,-37.6096534729004,
-27.7620830535889,-40.3307113647461,
-13.6192188262939,-36.0213546752930,
27.4042224884033,-47.4262657165527,
49.4073410034180,-57.8882179260254,
32.1999359130859,-43.7034530639648,
1.91161704063416,-15.4524822235107,
-12.3408708572388,3.87704968452454,
-11.7328481674194,12.6533164978027,
-16.4875774383545,20.4299793243408,
-27.5865306854248,20.2244930267334,
-25.0479164123535,0.113557934761047,
-1.65324139595032,-25.8818569183350,
30.9744224548340,-26.9866828918457,
49.0723114013672,-0.868689775466919,
37.8743591308594,23.8122615814209,
4.76881217956543,23.1720352172852,
-18.5329627990723,7.35638952255249,
-9.94042205810547,6.37268066406250,
15.5099992752075,20.9933147430420,
26.8503189086914,28.3779830932617,
20.3055992126465,17.9760589599609,
17.7323226928711,2.75964403152466,
28.9000473022461,-6.31367778778076,
32.2255897521973,-13.7235937118530,
4.73792028427124,-17.8128604888916,
-35.8327598571777,-11.4252920150757,
-51.8334312438965,5.70119714736939,
-38.9132957458496,17.0104370117188,
-30.2504138946533,12.9244537353516,
-31.3743247985840,8.53421974182129,
-13.2866210937500,18.4049377441406,
32.4756355285645,30.2458801269531,
65.6776275634766,15.5395336151123,
45.3619003295898,-22.2633037567139,
-1.36404800415039,-45.4514350891113,
-14.1068410873413,-42.5854682922363,
13.1417284011841,-36.9380874633789,
28.8220138549805,-41.5681266784668,
5.51105213165283,-34.3081016540527,
-18.6572341918945,1.81980741024017,
-0.827805161476135,40.9749183654785,
29.7555255889893,40.3531341552734,
14.5170879364014,5.63282871246338,
-40.4712829589844,-18.9589366912842,
-69.8356323242188,-19.3189983367920,
-40.0822067260742,-21.3349685668945,
14.9441461563110,-37.1167640686035,
44.1121520996094,-36.3619003295898,
43.8298912048340,-6.71093082427979,
36.9890060424805,9.90077686309815,
33.8847579956055,-20.9357490539551,
30.0370903015137,-60.6513442993164,
23.7515945434570,-46.7275543212891,
21.7842884063721,12.7271909713745,
9.48929119110107,45.4559211730957,
-23.8217792510986,12.0369024276733,
-51.4655952453613,-39.3125724792481,
-34.6407890319824,-43.1594924926758,
12.5389537811279,-0.972715377807617,
37.1478462219238,36.2870521545410,
19.0086498260498,45.8079071044922,
-10.2860355377197,38.8785858154297,
-19.0820007324219,23.1781425476074,
-17.9489498138428,-2.77729654312134,
-31.4699077606201,-25.0189647674561,
-36.9761695861816,-20.8864707946777,
2.63078689575195,1.15561306476593,
58.1631164550781,13.4682178497314,
62.3408317565918,8.25892353057861,
7.70784568786621,5.66706895828247,
-36.3437500000000,12.3643579483032,
-24.5004558563232,7.04261064529419,
3.43898820877075,-24.9421367645264,
-10.9094495773315,-52.5965309143066,
-40.8152465820313,-37.6610374450684,
-19.7857151031494,2.80100774765015,
42.9726524353027,26.7082328796387,
64.7146759033203,24.0434284210205,
8.83983325958252,16.9555568695068,
-50.5822944641113,14.7979803085327,
-33.8852462768555,2.27806401252747,
28.7601604461670,-19.9870471954346,
40.8420982360840,-26.9281139373779,
-19.7745323181152,-12.3288202285767,
-71.8793792724609,-1.27019524574280,
-50.5304908752441,-13.7358980178833,
5.82496356964111,-24.8836574554443,
21.5096836090088,-2.95179557800293,
-23.4030952453613,30.2254257202148,
-68.7000122070313,24.7617835998535,
-60.9528045654297,-24.5092697143555,
-18.8332519531250,-66.0970993041992,
5.61756610870361,-63.7397003173828,
-5.84000110626221,-36.5917053222656,
-22.2432327270508,-19.3960437774658,
-10.0115222930908,-17.3176040649414,
30.1767082214355,-12.3552789688110,
56.4673118591309,-9.23470211029053,
37.5229644775391,-24.4186172485352,
0.653633356094360,-48.3888778686523,
-4.13890314102173,-47.9243736267090,
25.3546848297119,-15.2972545623779,
37.3237800598145,11.9990663528442,
-5.24266386032105,5.71156978607178,
-68.8028030395508,-15.4578313827515,
-78.8197097778320,-15.7634992599487,
-21.5623359680176,-3.01737761497498,
33.7636528015137,-9.43494796752930,
28.9389133453369,-38.9314956665039,
-6.63722085952759,-53.0841407775879,
-8.44890022277832,-25.1963825225830,
29.8698253631592,21.8257942199707,
47.9022560119629,43.1851577758789,
12.2481298446655,28.7986068725586,
-33.8665351867676,8.04813003540039,
-30.4820251464844,2.61620330810547,
10.9613456726074,2.85187697410584,
33.6187934875488,-8.11061286926270,
8.01595401763916,-26.1820755004883,
-30.5023841857910,-34.9000892639160,
-39.9439315795898,-21.4625663757324,
-24.6540393829346,10.3986330032349,
-15.7051668167114,42.6023178100586,
-23.7752914428711,57.8656997680664,
-30.3002452850342,52.6653900146484,
-22.0182304382324,34.2201385498047,
-4.88971185684204,12.1836032867432,
11.0687379837036,-11.4104232788086,
19.0595836639404,-31.7304725646973,
20.1282424926758,-37.8445701599121,
20.0741233825684,-16.1466655731201,
28.2783527374268,15.4282560348511,
50.7970619201660,26.8857612609863,
69.4773635864258,12.6670331954956,
53.6841163635254,0.300021111965179,
1.66182279586792,9.53542995452881,
-45.3046417236328,17.2898197174072,
-48.5351638793945,-3.85904312133789,
-22.4473590850830,-41.8468894958496,
-10.3838176727295,-51.6403007507324,
-28.7042369842529,-20.2056903839111,
-48.0585975646973,15.8866615295410,
-42.0734786987305,20.4346542358398,
-23.6929588317871,4.18015384674072,
-22.1085147857666,5.83107519149780,
-34.5758972167969,29.5041790008545,
-30.2161369323730,46.7624855041504,
0.365286350250244,40.0669746398926,
32.4862365722656,19.2778301239014,
42.3464202880859,-2.77670383453369,
23.3196010589600,-25.9656829833984,
-10.1499013900757,-44.0406379699707,
-39.1892433166504,-44.3386421203613,
-41.1890182495117,-25.2629528045654,
-15.8312816619873,-12.5952434539795,
6.84615373611450,-25.7971935272217,
-1.11833095550537,-43.6203536987305,
-28.9379005432129,-29.7054080963135,
-35.2128677368164,7.15815067291260,
-7.22789859771729,19.8591308593750,
10.0373430252075,-4.53277015686035,
-17.6886215209961,-23.9226226806641,
-52.2246170043945,-8.90345478057861,
-33.7716865539551,13.7123098373413,
29.5817565917969,3.98084926605225,
65.4702529907227,-18.9299716949463,
43.7395629882813,-3.51446938514709,
7.27801799774170,44.4342155456543,
5.79692935943604,59.2127952575684,
23.1426715850830,17.6017837524414,
21.2949409484863,-18.8932685852051,
3.54877424240112,5.49946880340576,
-0.799350023269653,51.9761238098145,
8.18376541137695,44.6236152648926,
-6.22853755950928,-13.9134359359741,
-47.8104438781738,-45.7307319641113,
-76.6094055175781,-20.1141376495361,
-63.3191413879395,9.51214694976807,
-30.7180747985840,-9.22371101379395,
-4.31348609924316,-45.0531349182129,
15.9317283630371,-39.3547744750977,
34.3943939208984,2.85233235359192,
38.4413452148438,21.2524929046631,
26.1279315948486,0.591148972511292,
23.8022594451904,-13.2944192886353,
44.9266662597656,6.24682521820068,
55.3824996948242,33.7892227172852,
16.9838542938232,39.2930755615234,
-49.2016296386719,24.9085464477539,
-78.5969696044922,7.19458675384522,
-56.8732986450195,-12.8076333999634,
-38.9389038085938,-35.5472831726074,
-56.4303283691406,-40.8597793579102,
-67.9577713012695,-15.6752920150757,
-29.2370071411133,17.8110523223877,
30.8792762756348,25.8305492401123,
48.4436874389648,19.7921619415283,
11.0562591552734,35.6275138854981,
-29.0902557373047,60.3834037780762,
-34.6883354187012,43.5692901611328,
-20.7981491088867,-20.0403900146484,
-10.2048673629761,-68.5097885131836,
3.53126597404480,-49.6782302856445,
28.6478137969971,8.10090446472168,
39.0375976562500,32.7468032836914,
6.58071041107178,-0.578115582466126,
-39.3986854553223,-46.8567733764648,
-42.2440719604492,-65.4698486328125,
3.12308979034424,-53.6309509277344,
49.1259918212891,-28.4418201446533,
49.0123939514160,2.44215703010559,
10.4880695343018,25.4471645355225,
-26.3657131195068,13.0279312133789,
-32.2984886169434,-35.4429359436035,
-13.2544250488281,-72.2584381103516,
12.7689914703369,-56.2752265930176,
23.9462471008301,-3.51560759544373,
5.24738216400147,29.7924709320068,
-31.5527820587158,19.6820793151855,
-42.1108551025391,-8.33907032012940,
-6.63792705535889,-11.7348299026489,
34.2578239440918,16.2999553680420,
26.8718605041504,50.3474349975586,
-20.5867938995361,66.1709060668945,
-42.0595436096191,58.8479576110840,
-2.33343744277954,36.4381904602051,
49.2696990966797,17.2038173675537,
45.7161750793457,11.5431451797485,
0.693902730941773,9.91904926300049,
-13.4225835800171,-4.73256921768189,
25.8426971435547,-26.0206604003906,
62.4398536682129,-28.8702812194824,
53.8582572937012,-10.3504295349121,
29.5674934387207,3.45480227470398,
36.3406639099121,-2.89917850494385,
54.4744682312012,-10.6628532409668,
28.0137977600098,1.03861916065216,
-36.8017997741699,15.7751350402832,
-65.6174163818359,-0.704109668731690,
-19.8348426818848,-36.7840347290039,
45.4647026062012,-37.1842308044434,
50.8896598815918,12.8264636993408,
-5.30700349807739,59.6592369079590,
-55.0539131164551,47.1512908935547,
-55.2105751037598,-6.70308828353882,
-30.4418144226074,-43.2759819030762,
-12.0395107269287,-39.5591583251953,
-2.71661043167114,-27.3821048736572,
9.52474689483643,-32.8166923522949,
21.5024948120117,-42.2973899841309,
20.0016326904297,-36.8707351684570,
4.53704547882080,-28.4539947509766,
-2.18940401077271,-32.2977981567383,
11.1124191284180,-32.0363540649414,
30.7986812591553,-4.42543077468872,
33.0712738037109,32.3631896972656,
12.0932083129883,34.4157333374023,
-14.1735048294067,-2.89992213249207,
-14.1332893371582,-32.4807701110840,
25.4594326019287,-18.1027278900147,
70.9817428588867,17.6257286071777,
72.4985961914063,29.1272792816162,
23.2575302124023,11.5800647735596,
-33.5104026794434,-2.14245247840881,
-53.2353668212891,2.97650575637817,
-41.7036705017090,-0.751783967018127,
-32.2697029113770,-25.4326877593994,
-36.3056716918945,-44.8847999572754,
-29.3320789337158,-31.0309581756592,
-2.49297356605530,-4.36064529418945,
17.1118507385254,0.720172882080078,
12.2796936035156,-12.6180467605591,
1.29394936561584,-7.27705955505371,
8.96021556854248,24.2700176239014,
21.9814319610596,44.2643127441406,
8.59750366210938,18.4129199981689,
-20.8991565704346,-31.8436679840088,
-26.3577728271484,-58.5666770935059,
3.07636690139771,-51.5588226318359,
28.6030464172363,-41.0771980285645,
20.5952415466309,-48.5433540344238,
0.522539854049683,-62.9043540954590,
12.4942836761475,-62.1770210266113,
54.9062881469727,-39.5576553344727,
78.6625213623047,-7.49373722076416,
53.2584648132324,16.4606037139893,
-2.67627358436584,19.9723224639893,
-45.9124794006348,6.33415699005127,
-55.2609443664551,-9.22240734100342,
-32.3825912475586,-8.53036975860596,
13.7647848129272,5.24537897109985,
59.5382347106934,12.7199449539185,
66.4430541992188,3.82007646560669,
23.6220054626465,-4.56958723068237,
-31.9169750213623,-0.204447060823441,
-44.4951477050781,3.06301760673523,
-4.24526453018189,-7.56839179992676,
35.6040191650391,-25.7395019531250,
18.5862216949463,-25.7068176269531,
-40.0936012268066,-5.36976718902588,
-75.9772033691406,10.4781932830811,
-50.0002212524414,2.96714425086975,
6.95596599578857,-11.1595706939697,
35.1198577880859,-7.64735126495361,
8.39624404907227,12.2181358337402,
-30.5542068481445,25.3205051422119,
-28.5669555664063,22.6469364166260,
19.2722339630127,18.8381385803223,
65.4821624755859,23.9873371124268,
61.6634521484375,24.0347938537598,
20.1824398040772,-0.0417905449867249,
-9.36265945434570,-37.7132606506348,
6.11598920822144,-55.2529716491699,
45.4424705505371,-34.2781219482422,
60.6204338073731,8.73540019989014,
35.5206832885742,38.4618339538574,
-2.45316600799561,38.3347396850586,
-21.2857627868652,21.1216239929199,
-19.4898109436035,6.80942344665527,
-14.1249933242798,1.85114061832428,
-23.3750114440918,4.57210636138916,
-40.5642433166504,12.8028488159180,
-48.7978096008301,20.8086109161377,
-37.5340080261231,20.1062927246094,
-12.1748008728027,1.73144912719727,
15.3181238174438,-27.9234161376953,
28.7064933776855,-42.8593940734863,
25.9714984893799,-24.5099983215332,
13.7138299942017,15.7982931137085,
4.50386047363281,43.1223678588867,
1.74563956260681,39.9483146667481,
-5.62158060073853,18.1531696319580,
-25.9580898284912,10.3244562149048,
-47.5653877258301,26.5494537353516,
-52.2574615478516,42.1668052673340,
-34.0506553649902,33.4315185546875,
-8.90535831451416,10.7275876998901,
7.05942678451538,7.56114339828491,
16.3741245269775,30.6334571838379,
31.6717967987061,47.5604858398438,
48.4533233642578,31.3479461669922,
48.2292900085449,-3.89909029006958,
31.4151096343994,-22.9707126617432,
15.3666162490845,-18.9867515563965,
8.59644126892090,-20.3377246856689,
1.95719015598297,-39.2257423400879,
-14.6795053482056,-51.2221527099609,
-29.3362865447998,-33.1788177490234,
-23.8534049987793,-6.91626548767090,
-2.69388198852539,-4.77412319183350,
14.2513542175293,-19.7523403167725,
24.3900451660156,-16.0839996337891,
33.4281196594238,18.6373348236084,
34.7148056030273,53.8119468688965,
8.89911365509033,65.6648025512695,
-30.3938751220703,62.1492652893066,
-40.5054931640625,58.1540908813477,
-6.39543533325195,46.5418281555176,
25.9816055297852,17.5083885192871,
7.23579692840576,-12.3829421997070,
-45.7695465087891,-20.5975761413574,
-69.5440826416016,-17.2750244140625,
-36.2115058898926,-35.3846015930176,
9.99213790893555,-72.9887847900391,
15.3013772964478,-86.2243804931641,
-14.4832468032837,-51.6363945007324,
-34.4562492370606,2.33608555793762,
-28.2885189056397,30.3251857757568,
-16.2920570373535,23.8693046569824,
-16.7182712554932,10.4117507934570,
-25.8405685424805,16.4363307952881,
-29.1512794494629,34.3758163452148,
-20.1538143157959,42.5672836303711,
2.60532760620117,38.7064056396484,
32.6635665893555,28.9934425354004,
49.7027778625488,25.8666973114014,
37.2516860961914,34.4246215820313,
8.31943798065186,46.1751060485840,
-3.10811471939087,38.1275825500488,
18.7825374603272,5.69221544265747,
36.8419837951660,-21.5193691253662,
17.8550090789795,-7.76110172271729,
-16.8933105468750,25.7226219177246,
-24.1613292694092,25.6859283447266,
0.536808967590332,-27.2870998382568,
18.2709922790527,-75.7667160034180,
6.04774951934814,-52.1447334289551,
-16.0247688293457,20.9113655090332,
-20.5178775787354,56.4883880615234,
-12.3582429885864,19.2831153869629,
-10.3687391281128,-29.6828804016113,
-10.6736135482788,-27.9286270141602,
-3.09253478050232,10.3066492080688,
-6.61948108673096,23.6327877044678,
-38.6923866271973,-1.80931162834167,
-75.0930023193359,-29.2736968994141,
-65.1112442016602,-38.3907966613770,
-7.95355892181397,-48.0334968566895,
38.9919815063477,-61.2740859985352,
40.5339508056641,-47.8621788024902,
23.8360843658447,4.40858173370361,
31.0277347564697,48.9040298461914,
54.1240615844727,37.9267959594727,
53.2407646179199,-7.29302644729614,
21.7203121185303,-23.8282546997070,
-4.28929376602173,-1.16092967987061,
-7.62288522720337,14.0749645233154,
-14.5271482467651,-4.95488500595093,
-38.6338005065918,-33.8415145874023,
-54.9135856628418,-35.4807167053223,
-42.4813842773438,-9.16561317443848,
-18.6756572723389,13.1242685317993,
-7.65332984924316,18.8808917999268,
-3.29420471191406,17.5388183593750,
14.3528633117676,9.24765014648438,
31.0657386779785,-9.38922119140625,
25.4566783905029,-23.2550067901611,
5.05928039550781,-18.4238395690918,
4.98396825790405,-8.90710544586182,
25.6085815429688,-10.7259788513184,
27.6533946990967,-9.48123931884766,
-8.64135265350342,16.6733989715576,
-40.1271247863770,49.4790077209473,
-24.8020992279053,39.2890014648438,
18.7318592071533,-19.1939792633057,
37.3784866333008,-58.1468849182129,
17.5245075225830,-23.3273944854736,
-3.39994025230408,39.2540435791016,
0.442335724830627,40.3443908691406,
21.9211330413818,-17.1757526397705,
36.4425010681152,-43.1615676879883,
36.5592575073242,6.01282024383545,
28.4531269073486,61.6363105773926,
18.5019607543945,41.9118995666504,
9.81419277191162,-25.9865016937256,
10.2445678710938,-52.9010314941406,
16.4136848449707,-14.1099300384521,
17.4798870086670,21.4050312042236,
12.8718414306641,9.45446777343750,
16.6641235351563,-11.2860069274902,
21.7597351074219,2.03569412231445,
0.779854774475098,23.7492160797119,
-39.3457717895508,5.75985622406006,
-54.0312767028809,-33.8107070922852,
-17.7872409820557,-32.5292358398438,
29.9075546264648,12.3307685852051,
30.2458496093750,39.1161994934082,
-9.49984931945801,13.7287588119507,
-22.9326591491699,-24.2084903717041,
18.4706306457520,-28.7161388397217,
59.7473068237305,-10.5300216674805,
48.2621612548828,-18.4401435852051,
11.4270858764648,-51.4203948974609,
9.20439529418945,-58.0819358825684,
38.7201080322266,-20.1388511657715,
37.6125869750977,21.6574821472168,
-16.8026275634766,23.9856891632080,
-69.9393615722656,-10.9924259185791,
-61.9013519287109,-43.2785949707031,
-5.69057941436768,-44.5354804992676,
38.9161071777344,-18.8191719055176,
43.1209640502930,3.32946562767029,
25.2655200958252,2.90795779228210,
11.4519824981689,-6.77194166183472,
-0.818914830684662,5.05451345443726,
-13.9503202438355,48.5668487548828,
-13.9423875808716,91.7218093872070,
2.13689112663269,80.9313430786133,
14.1360902786255,15.8151988983154,
9.29916286468506,-35.5186729431152,
1.55948328971863,-20.2129783630371,
4.98669147491455,27.7605781555176,
11.2654981613159,46.3575744628906,
6.14545869827271,30.9387283325195,
-5.85458803176880,29.1611099243164,
-7.94299602508545,57.1394500732422,
-6.27524805068970,69.4110107421875,
-27.8495445251465,29.7398929595947,
-63.8012580871582,-22.3523559570313,
-68.3585281372070,-35.4663429260254,
-30.1505088806152,-24.1901760101318,
8.07592296600342,-36.7126083374023,
6.90470361709595,-67.0027236938477,
-12.9709186553955,-57.5342521667481,
-8.44133090972900,-5.31798458099365,
15.7701673507690,23.5182876586914,
19.0175113677979,-8.35774993896484,
-4.69037103652954,-45.8528442382813,
-10.6049442291260,-28.5520553588867,
14.1191339492798,18.4128379821777,
28.2474250793457,24.9736862182617,
5.26050043106079,-21.7974376678467,
-13.5627479553223,-55.7706680297852,
10.3055934906006,-37.2463722229004,
38.8168716430664,-0.376169681549072,
9.89047813415527,8.83919715881348,
-58.4105072021484,-5.61699390411377,
-81.2659072875977,-20.5910644531250,
-30.0753974914551,-38.5546798706055,
24.9303112030029,-61.3960876464844,
16.5528526306152,-60.3790473937988,
-21.8779850006104,-15.6437311172485,
-12.6538372039795,37.0248260498047,
46.2046852111816,48.1025466918945,
81.3366470336914,21.4035644531250,
59.9739227294922,10.8138446807861,
26.1472682952881,38.7520446777344,
21.0193214416504,62.6730041503906,
26.7695980072022,35.8683929443359,
12.3899250030518,-24.2097606658936,
-3.46121168136597,-61.3602256774902,
15.1478815078735,-55.7695541381836,
55.1299705505371,-23.9249248504639,
62.1693267822266,6.96957683563232,
19.2958583831787,17.9385738372803,
-29.7757034301758,2.35046386718750,
-40.0035209655762,-28.9824638366699,
-24.7128868103027,-47.2495613098145,
-11.8652563095093,-31.6619510650635,
1.00749778747559,-0.172723531723022,
25.8795013427734,18.1495971679688,
47.7435035705566,18.1939601898193,
36.4387321472168,19.6928749084473,
-4.50035667419434,29.3181514739990,
-37.8009681701660,17.9234676361084,
-37.7014923095703,-27.4763259887695,
-19.9920425415039,-66.9685058593750,
-16.7913990020752,-57.8209228515625,
-30.4353771209717,-11.2837476730347,
-38.5899658203125,28.8356113433838,
-27.4371452331543,35.0088729858398,
-1.31667470932007,21.8596229553223,
29.7662315368652,9.90424537658691,
47.9265594482422,-0.218279242515564,
36.6716766357422,-7.85913419723511,
5.56268882751465,-0.512928724288940,
-21.0078754425049,17.9066352844238,
-26.8841342926025,18.8055953979492,
-24.5894412994385,-16.7533035278320,
-30.9740200042725,-54.7009353637695,
-34.1086616516113,-45.4136276245117,
-11.6053495407105,-1.45190882682800,
23.7016429901123,18.3286437988281,
27.9366893768311,-13.1843976974487,
-6.64878273010254,-50.0381011962891,
-34.4186744689941,-39.3339233398438,
-22.5122528076172,8.78429222106934,
-3.90505218505859,36.8465347290039,
-22.8554897308350,18.9916419982910,
-63.3236045837402,-12.7539768218994,
-65.5134582519531,-24.5054206848145,
-16.9453582763672,-19.3208103179932,
24.6356029510498,-8.02361679077148,
14.2878074645996,9.31103897094727,
-19.6808395385742,26.7731418609619,
-20.9405345916748,16.3015003204346,
10.7455253601074,-30.0719814300537,
30.8462486267090,-72.0681762695313,
23.8196296691895,-63.9194412231445,
13.5168304443359,-15.1988315582275,
16.9755973815918,23.8048362731934,
15.8778762817383,24.7997627258301,
1.06125974655151,12.0446653366089,
-11.6724920272827,9.28415775299072,
-9.18048667907715,-1.33013391494751,
-0.423087596893311,-34.3288002014160,
5.18188810348511,-63.4542121887207,
21.7346744537354,-54.0861587524414,
56.7231140136719,-14.0817356109619,
79.3518676757813,19.9856777191162,
50.1072769165039,32.6560783386231,
-14.3946647644043,36.9159851074219,
-49.1238136291504,35.9319763183594,
-27.4483089447022,17.9224281311035,
13.4350843429565,-11.4851531982422,
32.4672126770020,-17.1451625823975,
34.4975395202637,15.2302942276001,
39.2821197509766,47.1458244323731,
43.0903434753418,36.1171073913574,
25.5053710937500,-5.96309089660645,
-3.60172033309937,-34.8526344299316,
-11.8316411972046,-35.5011978149414,
8.71366119384766,-25.3103942871094,
32.1944618225098,-15.9725475311279,
38.3305511474609,1.11593401432037,
34.8121910095215,22.7041473388672,
26.1864337921143,28.5126781463623,
4.94969511032105,13.5040321350098,
-28.9301471710205,8.97079086303711,
-44.0128479003906,35.3020896911621,
-24.4509391784668,61.3338050842285,
0.418612897396088,46.8467788696289,
-8.27908611297607,1.54608035087585,
-48.3534851074219,-21.3303966522217,
-74.8747787475586,-5.00452709197998,
-58.2805213928223,6.05402469635010,
-18.0962104797363,-20.0399475097656,
9.26035881042481,-54.5060119628906,
15.3121690750122,-46.6835098266602,
18.2611370086670,2.50227189064026,
28.8565406799316,36.7844848632813,
39.1838912963867,25.4585552215576,
40.9480590820313,-0.0191547870635986,
31.2923679351807,8.47343158721924,
16.0435848236084,46.3939971923828,
2.29602241516113,66.1346511840820,
-2.02343726158142,40.6414031982422,
3.13557386398315,-5.86915779113770,
8.52777385711670,-33.2211189270020,
10.2550945281982,-25.4665679931641,
8.06478977203369,1.37686133384705,
2.35195302963257,18.2164859771729,
-7.70670366287231,14.2900829315186,
-24.6398200988770,0.837054312229157,
-32.6919975280762,-6.33595848083496,
-15.4816856384277,-5.05081510543823,
15.4913892745972,-5.48044061660767,
28.4386520385742,-20.9900779724121,
14.3074169158936,-38.3310546875000,
-1.76584851741791,-32.1532783508301,
3.75574135780334,-0.0834062099456787,
19.3892765045166,31.7264366149902,
17.0418796539307,44.2590522766113,
1.20491456985474,47.7626113891602,
2.71168184280396,52.3410949707031,
26.1387157440186,50.8535728454590,
32.1085433959961,25.8864288330078,
-7.75529623031616,-7.81991386413574,
-56.1348991394043,-15.4780168533325,
-55.8930168151856,5.96698284149170,
-8.52474975585938,15.8840494155884,
23.9333629608154,-10.1825799942017,
1.90216898918152,-45.1109199523926,
-44.7716445922852,-49.3706474304199,
-60.1467514038086,-29.4932956695557,
-38.7253875732422,-21.4454898834229,
-14.4278497695923,-28.7890567779541,
-10.7483596801758,-20.3004608154297,
-16.7102317810059,9.58917808532715,
-21.2042503356934,26.9061660766602,
-28.3940773010254,7.32599353790283,
-32.7885742187500,-26.9853916168213,
-12.4981374740601,-34.6304664611816,
31.8154125213623,-20.2395744323730,
61.1734848022461,-15.3805522918701,
45.5252380371094,-29.5210723876953,
10.3803453445435,-39.1753349304199,
4.08114480972290,-28.5229549407959,
34.6727371215820,-12.3397998809814,
65.4966964721680,0.150468111038208,
66.6448669433594,15.8589620590210,
50.4754600524902,29.1005859375000,
39.4692306518555,21.0321311950684,
27.0480041503906,-8.87651824951172,
4.91899967193604,-26.9272880554199,
-16.0159149169922,-0.923769950866699,
-15.1980466842651,49.9856414794922,
-0.969789981842041,70.8819732666016,
6.38040685653687,42.5543098449707,
3.29129600524902,1.40499615669250,
3.56001114845276,-14.4468669891357,
9.04918193817139,-0.166613563895226,
3.06367540359497,26.3068885803223,
-15.9606904983521,48.6810035705566,
-25.9151496887207,52.7296066284180,
-11.1627531051636,25.5662231445313,
12.4495544433594,-16.4353637695313,
16.0158710479736,-29.1611804962158,
-2.05080556869507,13.9276638031006,
-23.9314365386963,70.6510848999023,
-40.4764060974121,74.2200698852539,
-55.6702957153320,11.0593357086182,
-60.9968338012695,-50.9803276062012,
-39.7070732116699,-42.4020347595215,
5.84147977828980,23.4057540893555,
43.2675666809082,69.6738052368164,
40.2918815612793,51.8374710083008,
2.43140697479248,-3.87647867202759,
-28.3129444122314,-38.0409355163574,
-22.0247726440430,-26.7845916748047,
16.1157321929932,1.26684546470642,
50.4771270751953,13.1141023635864,
51.8136215209961,9.48798084259033,
19.2464122772217,13.1484889984131,
-23.1414642333984,35.0629653930664,
-43.3753547668457,53.8595046997070,
-28.6897659301758,49.7133750915527,
2.78502798080444,25.9619407653809,
21.7357921600342,4.97484397888184,
16.0712108612061,5.41385841369629,
3.91404104232788,17.4691543579102,
6.86985778808594,19.6394176483154,
26.1303787231445,14.3985309600830,
36.3420715332031,17.6014633178711,
13.0458354949951,30.5827198028564,
-31.5109310150147,41.2428436279297,
-62.1269340515137,35.1170043945313,
-55.1299858093262,19.0865154266357,
-20.0659198760986,13.0360784530640,
8.64252090454102,13.1188058853149,
4.96378707885742,-0.0762408971786499,
-17.4578895568848,-31.5411987304688,
-27.1046791076660,-49.7027664184570,
-7.15001583099365,-29.7222862243652,
18.7155380249023,4.78326463699341,
21.7674674987793,5.92516136169434,
4.78866004943848,-29.1008987426758,
-0.282422840595245,-47.7463836669922,
26.0747604370117,-12.5714817047119,
49.7412414550781,40.0725860595703,
27.3679885864258,46.4563598632813,
-28.0312576293945,-2.07076716423035,
-57.4540367126465,-46.5008583068848,
-35.7992553710938,-40.9885749816895,
-4.32183218002319,-0.487305164337158,
-9.26295280456543,37.7279701232910,
-38.4281463623047,59.9629783630371,
-41.7168731689453,65.9457702636719,
-16.1806411743164,48.1156501770020,
-9.28880023956299,5.26806545257568,
-34.4032211303711,-33.3502960205078,
-41.2483024597168,-34.5726661682129,
8.05860328674316,-6.31291961669922,
70.1498336791992,13.8281850814819,
70.2428054809570,13.1371145248413,
6.98129892349243,10.8729295730591,
-47.7544784545898,20.4448833465576,
-47.1737403869629,22.2170429229736,
-24.0337219238281,2.72970223426819,
-24.2082042694092,-8.34125423431397,
-38.7628746032715,14.8500919342041,
-28.9785041809082,48.3803443908691,
4.75737953186035,49.6604804992676,
19.3757152557373,11.3014678955078,
-3.11357498168945,-23.7159233093262,
-29.8454685211182,-16.6913585662842,
-24.5075836181641,18.8948974609375,
-0.663958847522736,42.8426246643066,
12.1573247909546,27.9612274169922,
7.86510181427002,-12.0908803939819,
2.93235611915588,-45.4918594360352,
2.85337138175964,-42.8511886596680,
1.43673753738403,-1.17224633693695,
-6.28618812561035,44.6415214538574,
-6.47541666030884,47.8360214233398,
9.86036491394043,1.41351413726807,
27.2253532409668,-50.5428009033203,
25.2808475494385,-63.0272979736328,
4.23207855224609,-37.3932952880859,
-15.7405948638916,-9.13164234161377,
-17.8027381896973,0.0636593624949455,
2.49014163017273,-1.63073301315308,
33.1690902709961,0.183131277561188,
52.0902786254883,-4.16789197921753,
47.8654022216797,-20.3498668670654,
33.7157821655273,-31.2647361755371,
26.2669086456299,-19.6147060394287,
30.6884765625000,0.0523121356964111,
30.6689910888672,-2.50870990753174,
15.8864583969116,-27.4549598693848,
5.57124900817871,-38.9842758178711,
18.1958141326904,-19.4722747802734,
39.7591819763184,5.93768882751465,
37.5731315612793,7.51346206665039,
6.62659502029419,-9.23755264282227,
-15.9013195037842,-14.1954345703125,
-8.94724082946777,1.25459086894989,
5.73228406906128,6.40553140640259,
-3.54298329353333,-15.6315393447876,
-23.9696235656738,-46.5646438598633,
-12.7262487411499,-53.9604339599609,
37.0093421936035,-32.9010848999023,
76.0137939453125,-0.952544689178467,
58.6004638671875,21.8124923706055,
-2.64868307113647,24.5499343872070,
-52.1407546997070,6.08149385452271,
-56.7532272338867,-19.5328350067139,
-26.1617660522461,-28.8742027282715,
16.5714817047119,-13.3189029693604,
50.8951873779297,10.7386608123779,
60.4750709533691,15.5159730911255,
39.0174102783203,0.848555207252502,
3.60442709922791,-6.63565158843994,
-19.9862613677979,7.29896306991577,
-21.1039714813232,27.6585426330566,
-15.0748004913330,38.6283340454102,
-13.2801866531372,41.8364639282227,
-4.25672435760498,42.0993270874023,
17.3481025695801,34.6114578247070,
21.5158348083496,21.7531795501709,
-14.2670383453369,15.4546566009521,
-57.6433868408203,22.8409786224365,
-50.2406005859375,22.5960140228272,
2.87100219726563,-2.77320909500122,
34.1186256408691,-32.8578910827637,
4.26431798934937,-33.9186477661133,
-37.1711959838867,-4.92319154739380,
-20.3321456909180,14.0122451782227,
37.5593452453613,2.43598270416260,
58.1635513305664,-7.46965885162354,
13.5446109771729,16.3332328796387,
-35.7411460876465,50.9685134887695,
-36.0062675476074,55.8563919067383,
-13.7045669555664,26.4669456481934,
-19.7940635681152,-1.79963815212250,
-47.2708969116211,0.263853192329407,
-49.2632331848145,20.1550750732422,
-18.4385166168213,33.9599266052246,
9.34974575042725,29.6084613800049,
13.4711570739746,5.48418045043945,
13.1715211868286,-31.1377506256104,
30.0268363952637,-54.4256515502930,
43.2111091613770,-31.4154319763184,
23.8183650970459,20.8336143493652,
-14.1882572174072,34.2579612731934,
-30.0117969512939,-21.0558967590332,
-8.66114997863770,-83.5702209472656,
32.1850738525391,-71.2796325683594,
67.5315322875977,6.76873683929443,
68.6109313964844,57.4017791748047,
26.7233657836914,27.0614376068115,
-22.3655433654785,-29.8428802490234,
-25.4294509887695,-34.9635200500488,
27.1269512176514,3.92679882049561,
72.8512573242188,19.6551055908203,
48.7411422729492,3.67400312423706,
-21.7717895507813,7.88424444198608,
-52.7011184692383,45.9896202087402,
-16.0335655212402,64.5073852539063,
21.8613109588623,25.8849334716797,
2.93896698951721,-23.7447357177734,
-28.5506000518799,-24.7420177459717,
-7.92132949829102,8.34401988983154,
42.6103782653809,12.3338060379028,
49.9535522460938,-26.2194290161133,
1.62907361984253,-57.9250106811523,
-37.2255325317383,-44.9429702758789,
-22.2321987152100,-12.7939653396606,
3.97800683975220,9.01018905639648,
-5.94464588165283,33.5330276489258,
-32.0265998840332,67.1491165161133,
-28.5404968261719,75.8805923461914,
-5.76850032806397,39.0851745605469,
-1.76472020149231,-9.98630142211914,
-10.2454710006714,-20.1217021942139,
15.5143566131592,3.34074974060059,
60.9185028076172,12.3479766845703,
61.5291328430176,-10.6227960586548,
-0.926535606384277,-29.0291385650635,
-53.9375762939453,-19.1243553161621,
-32.0527458190918,-6.51634693145752,
28.9759769439697,-13.8123607635498,
43.3983993530273,-19.7096595764160,
-8.15435218811035,-0.582887887954712,
-58.0894393920898,20.7826328277588,
-54.8210983276367,12.2483386993408,
-27.0487155914307,-12.2009696960449,
-21.8245849609375,-6.40439414978027,
-35.8392677307129,33.5804443359375,
-40.8675842285156,61.3963890075684,
-35.8947601318359,44.2336692810059,
-41.6664619445801,2.24273490905762,
-58.0523071289063,-16.8357143402100,
-61.6751060485840,-2.60038638114929,
-41.5200881958008,13.7113943099976,
-9.74218750000000,11.2172231674194,
11.8424768447876,-2.22855401039124,
18.2435722351074,-10.1865158081055,
14.1437253952026,-1.59005308151245,
-1.26119756698608,18.5055541992188,
-16.7791118621826,27.4744033813477,
-8.88127517700195,9.43506145477295,
18.5772914886475,-16.7239685058594,
29.8208026885986,-12.9509716033936,
9.47990226745606,28.6463851928711,
-22.4983062744141,63.6071243286133,
-32.5997467041016,43.7298622131348,
-23.4423274993897,-12.0260410308838,
-19.6048927307129,-34.3975105285645,
-20.9005298614502,6.32279586791992,
-4.24508380889893,48.6847381591797,
24.3308658599854,29.4247341156006,
26.8542289733887,-25.7867374420166,
-9.26401710510254,-37.9107131958008,
-35.7458381652832,11.2174816131592,
-10.3072605133057,53.5636062622070,
35.4048805236816,30.8860054016113,
32.0914993286133,-27.0324707031250,
-26.0756912231445,-47.7003746032715,
-70.9107589721680,-20.7748908996582,
-49.7264633178711,2.51760005950928,
8.57523155212402,-7.08355855941773,
38.4959373474121,-22.4543228149414,
13.2008285522461,-16.5535030364990,
-31.0028114318848,-5.79611778259277,
-47.6605758666992,-15.9853191375732,
-24.4149799346924,-31.0723953247070,
21.6849822998047,-25.5419445037842,
56.3444938659668,-9.55559349060059,
54.6230697631836,-10.7683048248291,
21.2166385650635,-23.7440547943115,
-2.83164334297180,-11.9954490661621,
7.95688867568970,28.0836524963379,
29.9903526306152,51.5658912658691,
28.7453632354736,28.1219444274902,
10.9660081863403,-7.40060806274414,
12.5461063385010,-11.0328149795532,
38.1124382019043,3.58195114135742,
51.8930397033691,1.02509331703186,
24.7472152709961,-16.3557777404785,
-12.5940265655518,-15.4857406616211,
-16.0579051971436,2.93092656135559,
7.47606897354126,2.49180269241333,
19.7546539306641,-29.9915027618408,
19.2195339202881,-52.1244735717773,
31.6350135803223,-27.7017669677734,
54.5026435852051,17.6279525756836,
51.3351440429688,34.1006126403809,
13.4244365692139,22.8454551696777,
-18.3864231109619,14.8665704727173,
-16.3865756988525,13.7558584213257,
-8.12202835083008,-1.63534712791443,
-31.5912361145020,-25.7029457092285,
-66.6853179931641,-31.8851699829102,
-57.0098457336426,-18.3886909484863,
-1.19993281364441,-13.9838476181030,
42.0479469299316,-25.3739185333252,
39.5741958618164,-18.8770275115967,
25.9002780914307,20.2756614685059,
35.1900634765625,47.3834152221680,
44.1442108154297,19.7701606750488,
17.9491882324219,-26.0900611877441,
-22.4922180175781,-20.5785064697266,
-33.4990997314453,36.2751693725586,
-15.4476499557495,67.6875991821289,
-11.8645153045654,37.1110649108887,
-38.0376014709473,-10.3203191757202,
-50.2560729980469,-16.8938331604004,
-16.5828380584717,5.81697607040405,
26.4279003143311,13.5397186279297,
24.8717994689941,-2.22101449966431,
-15.7243099212646,-8.68203926086426,
-42.6660690307617,9.58485794067383,
-30.9762554168701,25.5548820495605,
1.41716265678406,22.6720466613770,
27.2437095642090,16.4811229705811,
28.0788688659668,19.5158863067627,
3.52380776405334,19.5378780364990,
-37.7082824707031,12.2302999496460,
-62.6462135314941,15.3842353820801,
-43.3291015625000,30.7071743011475,
4.29483318328857,36.3596801757813,
28.2537250518799,20.7176628112793,
7.83895492553711,13.1543912887573,
-13.5720586776733,35.9001350402832,
4.85103416442871,61.6504020690918,
35.7773208618164,39.3470230102539,
31.4075336456299,-21.2097187042236,
1.46469354629517,-50.3178863525391,
-0.826409876346588,-15.3260641098022,
35.7644309997559,32.7936859130859,
59.7528076171875,41.3762817382813,
28.8405151367188,27.6904544830322,
-25.7255096435547,32.5848388671875,
-45.8866348266602,47.5413856506348,
-25.2537536621094,25.7909164428711,
-3.18406677246094,-32.5543174743652,
-0.843707323074341,-70.8517227172852,
-0.884576022624970,-58.8737297058106,
9.06100368499756,-37.8361091613770,
13.4633388519287,-44.9675865173340,
4.76114416122437,-55.8793144226074,
-6.50226593017578,-31.0311813354492,
-11.1506776809692,6.54274749755859,
-13.8665008544922,3.14083385467529,
-16.1461944580078,-34.4332237243652,
-14.2930107116699,-44.4941329956055,
-7.71515560150147,-8.04777812957764,
-12.1833820343018,21.7795982360840,
-28.3105545043945,1.14336836338043,
-31.5254783630371,-36.9766616821289,
-2.05190587043762,-31.3306903839111,
25.5784358978272,9.80768775939941,
9.21991920471191,27.2333259582520,
-36.9095535278320,-3.18886041641235,
-50.9879875183106,-37.7870445251465,
-11.1391925811768,-36.8657531738281,
31.0176181793213,-22.5057353973389,
24.5466289520264,-26.0706577301025,
-8.88052558898926,-39.3218727111816,
-8.14313793182373,-34.3139076232910,
34.2495613098145,-8.53508949279785,
66.3158721923828,10.9928541183472,
52.5531425476074,4.95979261398315,
23.8162212371826,-8.07175827026367,
30.6510467529297,-1.47560381889343,
65.7577209472656,22.8767471313477,
74.3097076416016,41.3111267089844,
28.7492637634277,37.5024566650391,
-36.1607856750488,14.3312063217163,
-67.9188079833984,-8.19799041748047,
-52.2216377258301,-5.48125505447388,
-17.7557888031006,23.2967052459717,
0.829013764858246,43.7777099609375,
3.42039489746094,24.5747337341309,
15.1398792266846,-19.9620265960693,
43.0988311767578,-36.7030639648438,
63.8974609375000,0.00838851928710938,
47.1101455688477,58.0494308471680,
-1.39788627624512,76.0171279907227,
-35.7987136840820,41.1579933166504,
-18.8023643493652,0.633945584297180,
24.1904964447022,-1.12862062454224,
32.5135993957520,29.5350856781006,
-11.5521411895752,59.3985595703125,
-59.6866264343262,69.5222549438477,
-61.7192192077637,61.4411048889160,
-26.2793006896973,38.3969841003418,
-7.47240257263184,7.41268920898438,
-27.3847675323486,-18.1707324981689,
-44.3871459960938,-24.3600444793701,
-21.0918273925781,-24.6274738311768,
22.0233039855957,-42.1918029785156,
37.4460144042969,-68.7766418457031,
16.8038005828857,-69.1426696777344,
-5.97873449325562,-31.7700138092041,
-9.52677345275879,8.29919433593750,
-14.9104890823364,10.4479331970215,
-40.6774063110352,-14.6916666030884,
-64.6700744628906,-30.0433139801025,
-58.3005332946777,-31.4415149688721,
-24.1154785156250,-43.9661979675293,
7.20808124542236,-66.5786437988281,
18.7852230072022,-62.7830848693848,
21.7430458068848,-9.29059219360352,
24.0720520019531,56.4388618469238,
14.6073837280273,79.1928482055664,
-9.04785919189453,49.1703147888184,
-25.8178138732910,8.85470867156982,
-20.2312450408936,-3.99337887763977,
-3.11464095115662,7.12347555160523,
7.09841442108154,19.9941291809082,
9.48548793792725,15.1909370422363,
5.86688852310181,-12.6553115844727,
-9.37460231781006,-46.2195930480957,
-39.5168380737305,-53.0125160217285,
-60.6159095764160,-21.9070320129395,
-40.6208610534668,15.1188840866089,
14.6888580322266,20.9289207458496,
53.4772377014160,-1.00248730182648,
43.9142532348633,-5.08727693557739,
7.04382324218750,26.6581420898438,
-20.3168163299561,52.4457435607910,
-29.2086925506592,27.8496513366699,
-34.1478195190430,-17.5144100189209,
-36.9785995483398,-18.6674289703369,
-31.1926364898682,21.7788333892822,
-25.8153915405273,41.2914505004883,
-35.3435287475586,13.2609519958496,
-49.7004814147949,-15.2341156005859,
-38.4351577758789,0.558195948600769,
0.745197534561157,25.9317855834961,
29.9524269104004,3.24455547332764,
20.4515647888184,-46.5263137817383,
-6.65925884246826,-48.8829383850098,
-8.05025100708008,10.8395462036133,
13.8510484695435,55.7262496948242,
27.9366111755371,29.6149330139160,
23.3272590637207,-22.9712848663330,
12.6561079025269,-30.6442565917969,
10.6616973876953,-0.746506690979004,
11.3996286392212,9.02235031127930,
7.41647291183472,-10.0144844055176,
3.55789017677307,-8.73889350891113,
3.55079746246338,29.8494606018066,
0.214782267808914,60.1772804260254,
-4.49125289916992,45.2719535827637,
6.22012710571289,11.6004114151001,
28.3503799438477,4.81333923339844,
23.9428615570068,16.9900455474854,
-23.6367893218994,8.24603843688965,
-67.9597930908203,-17.8825950622559,
-53.3855247497559,-24.9551029205322,
11.2409448623657,-12.2027921676636,
59.7314758300781,-10.5975303649902,
56.6199989318848,-24.4452228546143,
33.7518119812012,-26.5049648284912,
30.5347843170166,1.58419346809387,
28.3809719085693,36.0297508239746,
-7.58136034011841,45.9488792419434,
-56.9895744323731,34.0265045166016,
-62.9068489074707,18.1500244140625,
-22.6638622283936,-1.79349315166473,
5.38927173614502,-23.4131813049316,
-12.6489620208740,-22.0695190429688,
-38.6797294616699,16.0999584197998,
-22.6647357940674,51.0702056884766,
20.7240085601807,32.8720741271973,
38.6870346069336,-17.1776771545410,
21.4134254455566,-31.1475448608398,
4.34415912628174,15.0251235961914,
11.4650058746338,66.5968246459961,
18.9636669158936,65.5061798095703,
5.25789880752564,21.1291332244873,
-5.53086900711060,-16.5500431060791,
5.84225177764893,-26.6520824432373,
19.0469055175781,-30.9411125183105,
2.84017753601074,-39.7951240539551,
-26.6305522918701,-39.9751358032227,
-26.9561462402344,-27.1440296173096,
6.07846212387085,-12.0075254440308,
30.4312191009522,1.49320983886719,
16.2381362915039,26.0378303527832,
-13.2754917144775,56.0404701232910,
-24.7157325744629,63.4789581298828,
-21.2138500213623,42.2744064331055,
-24.0334339141846,19.4552307128906,
-25.6735000610352,19.9861965179443,
-4.58899021148682,31.0464286804199,
28.2573566436768,20.5733699798584,
40.1243095397949,-18.6210727691650,
24.8686027526855,-51.3408164978027,
10.2571649551392,-47.5949935913086,
14.8575553894043,-14.3493556976318,
15.8231420516968,20.0900535583496,
-10.6202602386475,29.3983612060547,
-43.0004043579102,8.17015457153320,
-41.9854660034180,-29.3020992279053,
-8.11864757537842,-49.3200607299805,
19.8634319305420,-34.3853340148926,
19.4814453125000,-2.16383957862854,
8.17094039916992,11.2736759185791,
0.323702812194824,1.58618640899658,
-13.0477914810181,-3.18916511535645,
-38.1706314086914,15.7581071853638,
-48.1365013122559,32.4809112548828,
-20.0500144958496,14.4092607498169,
28.5605564117432,-27.3527832031250,
55.9389305114746,-41.8465728759766,
46.4071884155273,-9.65149688720703,
31.3333835601807,31.3069610595703,
35.7836532592773,41.9783134460449,
43.2271080017090,25.3712329864502,
27.8432140350342,14.4283428192139,
-7.09367179870606,21.0947208404541,
-31.7612476348877,27.5789852142334,
-30.5777797698975,20.7798137664795,
-11.0790319442749,9.74176216125488,
3.87254548072815,3.06571841239929,
0.0338527262210846,0.816664993762970,
-22.0168132781982,-0.161907196044922,
-43.3875312805176,6.27636146545410,
-37.9936599731445,25.7442893981934,
0.152727529406548,40.9228515625000,
39.8706321716309,31.8877792358398,
38.6183929443359,2.86082267761230,
-11.6069755554199,-22.4910392761230,
-61.8430938720703,-29.4642753601074,
-68.9063491821289,-18.1124629974365,
-37.2192649841309,0.596851050853729,
-3.31900334358215,13.6510372161865,
12.3857250213623,15.4176425933838,
16.2782993316650,6.95011425018311,
23.5789184570313,2.17395353317261,
31.2168025970459,14.5354785919189,
33.4436225891113,33.0729255676270,
30.5978507995605,21.5131759643555,
25.0426406860352,-27.8027992248535,
17.1571464538574,-70.9654159545898,
19.6774044036865,-63.3538970947266,
45.6361618041992,-17.4738712310791,
79.5628128051758,8.95702934265137,
78.0433197021484,-9.98946762084961,
24.5726451873779,-34.5096969604492,
-28.8329219818115,-20.9610881805420,
-21.5716247558594,13.5987386703491,
33.4418449401856,22.7398872375488,
63.8798599243164,3.91979217529297,
23.2911014556885,-2.73679471015930,
-45.9017143249512,17.7044601440430,
-74.8349304199219,25.7234725952148,
-57.5216407775879,-8.39098739624023,
-36.7825736999512,-47.3279380798340,
-35.3086547851563,-35.8680305480957,
-30.4165458679199,20.3874435424805,
-8.64938735961914,52.7840843200684,
13.3884944915771,20.9037246704102,
17.4880638122559,-42.0224647521973,
15.3724317550659,-64.6614990234375,
21.9220981597900,-24.8371105194092,
21.8870773315430,28.9160728454590,
-1.56544172763824,42.8647003173828,
-34.6170883178711,12.9335708618164,
-45.2212448120117,-17.3736572265625,
-27.7268314361572,-10.3843021392822,
-15.5727958679199,26.1698284149170,
-28.8266124725342,46.2864532470703,
-45.6717453002930,23.9602680206299,
-38.8937492370606,-18.2485771179199,
-18.9619026184082,-37.9986190795898,
-11.9124402999878,-29.0243263244629,
-24.9209766387939,-18.6616764068604,
-37.9900398254395,-24.3662872314453,
-38.0554504394531,-26.2486228942871,
-27.7084655761719,2.11402893066406,
-20.3209629058838,45.8924827575684,
-17.0541210174561,63.3914146423340,
-16.6225452423096,45.8161010742188,
-23.9661788940430,27.3594474792480,
-39.2474555969238,29.5201930999756,
-48.2408485412598,34.3360786437988,
-35.8122673034668,8.85194969177246,
-8.36292552947998,-36.3897972106934,
21.0667495727539,-58.1472244262695,
36.6293716430664,-39.9917297363281,
30.6230411529541,-14.0678195953369,
2.89347410202026,-14.3109540939331,
-23.9468879699707,-35.1043586730957,
-21.3937835693359,-46.4233970642090,
21.2745647430420,-33.7441749572754,
65.9388961791992,-14.1802310943604,
63.9890403747559,-1.57543611526489,
13.7907314300537,10.9176540374756,
-30.1368579864502,33.7020721435547,
-26.1952972412109,57.1596450805664,
-1.72467994689941,66.7352981567383,
-8.24704933166504,54.8357658386231,
-49.5022010803223,29.9772357940674,
-73.5801696777344,5.01711225509644,
-47.7862854003906,-10.0779647827148,
4.98248100280762,-15.4282360076904,
39.3602218627930,-13.6182851791382,
45.2269668579102,-6.01139688491821,
46.2306060791016,5.90697431564331,
51.5310440063477,20.6274452209473,
50.8658981323242,29.3957424163818,
40.1727294921875,19.1770114898682,
29.8276653289795,-5.15540695190430,
21.6468772888184,-16.9822483062744,
5.35134696960449,-1.56863105297089,
-16.9578285217285,17.8425769805908,
-28.4323844909668,13.7693023681641,
-21.4707756042480,-9.21544075012207,
-7.65325546264648,-20.0904502868652,
-2.39304542541504,1.27107298374176,
-3.36304497718811,31.7773151397705,
-6.91942119598389,44.8931083679199,
-19.5813331604004,45.5288124084473,
-45.8102836608887,50.4180183410645,
-61.9545097351074,46.2397689819336,
-40.0495681762695,9.03431415557861,
0.488854408264160,-42.3914756774902,
13.0312919616699,-57.4505653381348,
-14.8808021545410,-24.5327377319336,
-37.6718177795410,1.93916130065918,
-20.5429782867432,-30.1257667541504,
14.6041631698608,-86.3872528076172,
23.3365688323975,-87.6600799560547,
-0.484818935394287,-20.3912944793701,
-24.4746589660645,38.6887969970703,
-24.0891189575195,26.6200218200684,
-8.23788833618164,-19.0404548645020,
9.01626300811768,-21.3051815032959,
27.9020843505859,23.6167812347412,
44.5461578369141,47.5347442626953,
42.4935569763184,15.5056381225586,
24.2293071746826,-30.7070693969727,
9.96435928344727,-37.0248756408691,
10.0573406219482,-14.4227981567383,
5.07850551605225,-6.25901794433594,
-9.70888519287109,-18.5922927856445,
-11.9280290603638,-23.2249259948730,
11.8398532867432,-9.96907711029053,
32.9674682617188,-4.10924339294434,
16.8527622222900,-10.9965963363647,
-17.9898567199707,-6.57914018630981,
-21.9850254058838,14.7317733764648,
13.0051355361938,27.3779201507568,
32.7800636291504,11.7606935501099,
1.04464888572693,-12.5999526977539,
-47.1687622070313,-18.4086112976074,
-57.5860824584961,-5.78607988357544,
-29.9436206817627,3.98680543899536,
-4.83694458007813,7.91718912124634,
3.84724140167236,21.7239131927490,
12.5810546875000,34.9152259826660,
30.1568126678467,22.7604560852051,
37.4196090698242,-1.43340992927551,
19.5405769348145,4.06909513473511,
-10.8508586883545,39.3898887634277,
-36.7915344238281,52.2902450561523,
-54.3183212280273,12.6895484924316,
-59.4176788330078,-40.9656867980957,
-38.9985122680664,-52.9794006347656,
1.80170929431915,-33.5481719970703,
24.2266178131104,-32.6572151184082,
4.79863309860230,-54.6564178466797,
-25.9354343414307,-46.0441398620606,
-22.5584926605225,8.51350212097168,
9.60012149810791,48.9750328063965,
26.2343235015869,25.6282482147217,
7.88414192199707,-27.2807502746582,
-13.7649965286255,-43.9419784545898,
-5.34115743637085,-22.7680530548096,
18.0602474212647,-17.1527328491211,
24.1519241333008,-41.1623725891113,
10.9272174835205,-45.4247093200684,
4.38901615142822,-1.52020359039307,
9.83945465087891,49.0534896850586,
7.80150127410889,53.1624374389648,
-8.26047325134277,20.0725326538086,
-20.7982578277588,5.47884845733643,
-18.4365139007568,25.5024223327637,
-9.07743263244629,40.9496803283691,
-2.55252456665039,22.4867382049561,
5.84694910049439,-8.58360004425049,
23.5122909545898,-18.5471534729004,
45.6201362609863,-6.66519880294800,
57.3867225646973,5.98427200317383,
56.2210121154785,5.76782560348511,
47.8649482727051,7.62392091751099,
33.6419639587402,25.4182453155518,
12.3375005722046,48.3444862365723,
-5.72208738327026,52.5836029052734,
-6.16219186782837,29.8311042785645,
3.27506732940674,-0.317181825637817,
-0.586095631122589,-13.3389749526978,
-24.7529640197754,2.65234279632568,
-44.3362426757813,30.4073352813721,
-35.2839469909668,41.5214614868164,
-5.05522966384888,27.2751750946045,
11.1721525192261,13.5374307632446,
-5.49268770217896,23.7601871490479,
-37.0256233215332,49.9639358520508,
-52.8389549255371,65.6792755126953,
-41.0780372619629,51.3089294433594,
-19.2498073577881,15.9801712036133,
-3.05192899703980,-20.7412738800049,
-0.0682814568281174,-45.8487625122070,
-4.15898799896240,-53.4215888977051,
-8.50937271118164,-35.6008224487305,
-6.86086845397949,3.74724245071411,
-2.42419934272766,35.4551124572754,
-2.93331480026245,40.5625190734863,
-9.88861846923828,32.6671905517578,
-16.8773174285889,39.7819290161133,
-16.4331607818604,56.5140342712402,
-9.79324436187744,41.0108337402344,
-1.22319173812866,-19.0672302246094,
9.56078338623047,-75.1499862670898,
27.1109542846680,-71.2443237304688,
43.3937950134277,-24.9904479980469,
39.0658798217773,-4.79500961303711,
16.2500114440918,-34.4097137451172,
-5.12844848632813,-55.5968017578125,
-9.54826164245606,-21.1321315765381,
-8.38502979278565,31.4527111053467,
-15.4046907424927,36.5467147827148,
-21.7286052703857,-9.36319160461426,
-9.36965179443359,-37.9655342102051,
13.6411905288696,-15.1301822662354,
21.3818931579590,20.4765739440918,
8.96970939636231,22.6898365020752,
4.41624832153320,3.99169397354126,
23.5477313995361,3.44101524353027,
37.2868080139160,20.2855072021484,
16.0355281829834,19.6635437011719,
-25.9243850708008,-7.12900543212891,
-46.0922927856445,-22.6297626495361,
-30.0847244262695,-13.2707586288452,
-8.80246448516846,-6.34741926193237,
-9.70321846008301,-27.8170528411865,
-22.1660785675049,-57.1140213012695,
-22.5248794555664,-55.6549606323242,
-9.78539752960205,-15.1344795227051,
-1.20083320140839,28.4503364562988,
2.37683939933777,41.8435173034668,
12.6150550842285,30.9744014739990,
25.8266448974609,20.9065799713135,
17.0419692993164,21.3395805358887,
-19.3520011901855,21.1781349182129,
-52.3521919250488,6.07763195037842,
-46.4912910461426,-25.9386749267578,
-13.0600757598877,-56.1176872253418,
9.40515041351318,-56.8932762145996,
-3.09301710128784,-26.0689640045166,
-30.2154884338379,6.26820945739746,
-40.0740699768066,8.51579189300537,
-29.6244144439697,-15.7083921432495,
-18.3298091888428,-34.3694152832031,
-17.6682052612305,-26.1397590637207,
-16.9734096527100,-0.171982884407043,
-9.19019031524658,14.9442958831787,
0.944813609123230,13.4882221221924,
7.82246017456055,6.80719280242920,
12.6181659698486,-4.23495435714722,
23.3141517639160,-18.5688743591309,
41.3952255249023,-23.2924823760986,
59.5381355285645,-5.20645284652710,
65.3138275146484,21.4786224365234,
59.3166618347168,26.0709590911865,
47.4969253540039,6.67205905914307,
37.9963378906250,1.09511744976044,
31.9096698760986,25.3131618499756,
15.6694002151489,44.5196266174316,
-18.6671791076660,14.8074779510498,
-46.3972091674805,-40.5528907775879,
-38.1282081604004,-55.8366661071777,
-3.59715938568115,-12.1569881439209,
10.8728780746460,26.5796298980713,
-17.7485637664795,9.94026184082031,
-49.9447326660156,-32.9963302612305,
-37.1095008850098,-39.5810012817383,
6.67492818832398,-2.39619588851929,
10.8582601547241,31.0889816284180,
-44.4132461547852,31.9333839416504,
-86.9224853515625,19.0690841674805,
-51.1635665893555,11.1475744247437,
25.5981445312500,-1.24204695224762,
49.6163635253906,-30.1264572143555,
2.47833299636841,-52.9382400512695,
-41.2272491455078,-49.5301742553711,
-19.1857395172119,-37.3704299926758,
33.2219848632813,-47.3838577270508,
51.9483947753906,-69.3261947631836,
38.8036346435547,-64.7091140747070,
36.0535697937012,-29.4024772644043,
44.6656799316406,11.3786716461182,
21.5763759613037,35.9344329833984,
-35.4370994567871,40.5881080627441,
-60.9396820068359,30.2485828399658,
-16.5566291809082,7.89271879196167,
43.9163475036621,-12.2783098220825,
47.8385009765625,-3.88450980186462,
2.44039297103882,30.5786590576172,
-25.5014991760254,50.1579208374023,
-1.68739390373230,36.4657592773438,
41.5500259399414,15.5996608734131,
53.8832015991211,14.4573678970337,
32.3119392395020,8.06958866119385,
5.76833534240723,-31.1433029174805,
-9.79696369171143,-74.0643997192383,
-9.80298519134522,-59.1448097229004,
6.87841892242432,7.60212421417236,
16.8873195648193,53.2524337768555,
-5.72096061706543,29.3747806549072,
-47.0359611511231,-20.9757156372070,
-56.4925003051758,-23.8845958709717,
-16.6378517150879,19.4059448242188,
16.6597175598145,43.4979362487793,
-12.1461048126221,14.1608419418335,
-70.1754455566406,-35.8730506896973,
-72.0174255371094,-57.6247253417969,
-1.88569331169128,-45.7673606872559,
49.7483673095703,-19.6919898986816,
17.3438320159912,-3.09080648422241,
-44.1342353820801,-4.64341974258423,
-42.5689392089844,-21.2925491333008,
20.4923572540283,-32.1948051452637,
52.6419944763184,-14.0968484878540,
8.81837654113770,21.4856395721436,
-45.7458801269531,35.5489501953125,
-36.5441780090332,4.65263319015503,
16.4116592407227,-33.8240318298340,
38.5258827209473,-25.0881462097168,
6.39772415161133,27.9965591430664,
-30.6959037780762,65.3363647460938,
-27.6088447570801,54.9189300537109,
-3.58159255981445,31.1863498687744,
-4.07750272750855,36.1229553222656,
-26.9329319000244,62.3794708251953,
-32.7625427246094,67.2431335449219,
-6.25437164306641,36.8265762329102,
27.2936687469482,6.84878969192505,
28.1799240112305,0.739365458488464,
-6.26213932037354,0.699660181999207,
-30.6168632507324,-17.1917304992676,
-12.7907629013062,-46.7801284790039,
24.6739387512207,-60.6039581298828,
33.0265922546387,-52.0538139343262,
-2.09911847114563,-40.0170745849609,
-41.5021858215332,-30.5746021270752,
-43.8873176574707,-12.8721837997437,
-21.1448535919189,8.89403915405273,
-19.9238357543945,11.3236293792725,
-52.9102401733398,-15.6041040420532,
-74.4182586669922,-43.0356979370117,
-47.0069999694824,-27.6551704406738,
6.38090085983276,26.4923763275147,
28.4418144226074,64.8474197387695,
-0.119949340820313,48.5077056884766,
-42.2377624511719,-3.98361420631409,
-53.2436943054199,-37.4665756225586,
-29.2228679656982,-25.2793922424316,
3.37877035140991,9.76972675323486,
26.6913337707520,28.6903438568115,
38.8680305480957,19.8664779663086,
46.0262947082520,5.73631858825684,
51.4215545654297,6.65072441101074,
53.1273040771484,20.7165966033936,
48.5160789489746,29.1045875549316,
39.0326805114746,20.3065452575684,
26.5423221588135,1.94025957584381,
17.2324390411377,-2.73889636993408,
14.7255458831787,14.0347728729248,
15.4401092529297,37.5318069458008,
11.3085689544678,43.6096572875977,
4.23805570602417,30.5861549377441,
-2.59340667724609,17.4104709625244,
-12.1508159637451,16.5443649291992,
-24.3137550354004,21.2892074584961,
-31.6849689483643,16.5716533660889,
-24.2834014892578,11.7355327606201,
-7.72975254058838,23.6698951721191,
-0.488936722278595,44.3783264160156,
-8.07710456848145,46.5996742248535,
-19.3985538482666,21.9024200439453,
-19.2117652893066,1.84651553630829,
-14.5181941986084,16.3769989013672,
-17.4038887023926,53.3797225952148,
-25.1412887573242,68.3571395874023,
-22.6332244873047,44.6762886047363,
-9.50980472564697,11.5825462341309,
0.399491518735886,-3.04003906250000,
-1.63065969944000,-7.25309514999390,
-3.83423948287964,-22.4215488433838,
4.14584779739380,-46.5295982360840,
12.4870567321777,-51.6861763000488,
7.47592449188232,-27.3412628173828,
-2.64888262748718,1.46335089206696,
2.16985797882080,11.8057317733765,
19.4036731719971,9.03308391571045,
21.3144073486328,12.7621049880981,
-4.62663316726685,21.9072360992432,
-32.4470901489258,20.1766281127930,
-25.1807956695557,-0.409903168678284,
11.3438434600830,-20.4085941314697,
33.8892173767090,-11.1551160812378,
13.5247392654419,23.6284065246582,
-22.9933052062988,44.3689918518066,
-31.9056568145752,22.3997650146484,
-8.53048133850098,-27.3338203430176,
12.7721920013428,-54.3325271606445,
12.2329759597778,-29.9190597534180,
8.19566345214844,15.6156101226807,
21.2145996093750,29.5239353179932,
36.7374916076660,8.99272537231445,
25.1684856414795,-5.55955076217651,
-8.40858268737793,8.58636856079102,
-29.4541835784912,19.5234546661377,
-25.9132213592529,-8.59091949462891,
-20.7831516265869,-52.6800308227539,
-27.6598930358887,-58.0900764465332,
-26.1589775085449,-15.8185253143311,
-1.59879517555237,24.5191802978516,
20.7819709777832,20.0247344970703,
8.41985797882080,-5.92029571533203,
-20.3765125274658,-8.34868812561035,
-21.6109600067139,14.9806022644043,
7.30171203613281,27.4779434204102,
20.3490886688232,8.35667324066162,
-7.00529813766480,-21.1605377197266,
-37.9813117980957,-35.0633773803711,
-29.1032104492188,-30.2358570098877,
2.99532461166382,-17.0687580108643,
10.3400688171387,-1.43426239490509,
-10.1705760955811,7.35037326812744,
-16.2739562988281,-4.13025808334351,
12.2342567443848,-35.2939605712891,
43.3419494628906,-58.9850082397461,
35.9229621887207,-47.9516601562500,
0.365180730819702,-5.65348625183106,
-25.5368061065674,29.4934062957764,
-24.4932289123535,35.4177780151367,
-12.0920486450195,23.3531684875488,
-8.29292869567871,9.68818473815918,
-12.8642196655273,-2.57891464233398,
-16.9949226379395,-19.1216583251953,
-23.7015819549561,-33.6899452209473,
-30.6183128356934,-36.1415367126465,
-27.7025108337402,-30.2059898376465,
-9.89517116546631,-26.6752452850342,
12.6656122207642,-24.0175533294678,
18.1448898315430,-14.3431539535522,
-6.03827667236328,-4.43017244338989,
-43.0659751892090,-12.9258480072021,
-55.2895240783691,-40.6444129943848,
-24.7751197814941,-57.2731590270996,
23.0027122497559,-33.7499618530273,
44.0112190246582,7.45072937011719,
20.2028121948242,20.8028507232666,
-14.7098321914673,-10.7609195709229,
-12.9907493591309,-51.2272911071777,
27.9107284545898,-53.7938652038574,
59.9561538696289,-13.3941888809204,
45.2646903991699,30.7521400451660,
5.75986671447754,41.8318214416504,
-10.9517393112183,21.5169372558594,
4.66421413421631,-0.0274784564971924,
18.8531341552734,0.124125450849533,
5.05318593978882,16.4084682464600,
-20.4958000183105,22.6979846954346,
-22.4158554077148,1.67453765869141,
-1.54209661483765,-32.6261482238770,
13.4682903289795,-47.9075393676758,
11.1893053054810,-30.0809364318848,
6.12053966522217,1.76535797119141,
4.71460247039795,23.8674812316895,
-5.70015716552734,33.0489578247070,
-26.4746856689453,38.4814300537109,
-31.6967029571533,39.9019699096680,
-3.82090520858765,26.5452709197998,
27.6356906890869,-0.639247238636017,
21.0137958526611,-10.6556987762451,
-11.0549173355103,9.73552227020264,
-21.9527568817139,34.8410987854004,
11.1909456253052,33.5946273803711,
49.6262512207031,11.8021621704102,
53.3132553100586,1.74529433250427,
37.3523330688477,14.3021221160889,
36.6056213378906,27.8355293273926,
44.3521461486816,28.2005825042725,
28.3170852661133,27.5790863037109,
-9.77346229553223,31.9518756866455,
-31.8974628448486,24.0996894836426,
-15.9992456436157,-4.54554128646851,
16.3531856536865,-23.1351776123047,
30.5160121917725,4.08602237701416,
19.7110881805420,55.9177436828613,
-6.90012645721436,70.5205383300781,
-46.5602569580078,25.9518508911133,
-82.9735870361328,-26.2346992492676,
-83.5594482421875,-36.1529922485352,
-35.9492378234863,-10.9462852478027,
17.7809543609619,7.18575763702393,
24.9836673736572,-0.140794098377228,
-0.973757982254028,-9.32205390930176,
-8.81792736053467,-0.964608728885651,
15.6496114730835,15.4640140533447,
27.2062320709229,24.4003829956055,
-3.30285167694092,26.9299831390381,
-40.5245933532715,22.9007034301758,
-34.2161521911621,14.0373668670654,
5.21696996688843,9.15069389343262,
18.0770263671875,23.6968345642090,
-18.0606918334961,42.2444267272949,
-60.7742919921875,26.5688037872314,
-66.7628326416016,-31.8639030456543,
-37.0214805603027,-78.2225646972656,
3.92373585700989,-61.6137847900391,
38.5177230834961,3.86083698272705,
53.7765655517578,44.0223083496094,
40.4093475341797,20.9935512542725,
6.70099067687988,-20.5181179046631,
-19.6157913208008,-19.9724159240723,
-19.1229496002197,20.7752532958984,
-10.6609745025635,53.0886192321777,
-21.2333469390869,51.2382278442383,
-48.5973548889160,25.0219459533691,
-62.7259216308594,-6.46568489074707,
-52.7377853393555,-36.1503219604492,
-39.7439956665039,-53.7487335205078,
-32.8018951416016,-49.5125427246094,
-15.6437454223633,-33.2841110229492,
14.8709678649902,-36.2946052551270,
29.6018218994141,-59.6239624023438,
12.4797334671021,-62.2842559814453,
-17.9004993438721,-22.7599716186523,
-24.7065620422363,22.9918460845947,
-3.60828685760498,20.4415626525879,
21.8908252716064,-11.8722877502441,
36.9422836303711,-13.4114809036255,
45.1088752746582,28.6742115020752,
43.2911071777344,58.0160255432129,
21.5343780517578,34.3080368041992,
-6.79273891448975,-9.07282161712647,
-8.35588264465332,-12.7778549194336,
23.4870052337647,13.2116861343384,
47.1494483947754,14.1711177825928,
35.4340820312500,-20.4514217376709,
11.4392566680908,-39.9992675781250,
17.1734218597412,-10.8173894882202,
47.3601722717285,33.5038833618164,
56.8163948059082,50.4050292968750,
24.4297962188721,40.5415725708008,
-17.2504711151123,37.0487174987793,
-28.7035007476807,41.1318550109863,
-11.3615236282349,32.9336280822754,
7.01686286926270,10.7934761047363,
14.7207841873169,2.21374034881592,
17.0888614654541,18.4673614501953,
14.3589611053467,38.0613174438477,
-0.485998988151550,35.3892440795898,
-21.2158145904541,14.0540304183960,
-30.9533252716064,-7.23192405700684,
-23.8157691955566,-25.8721218109131,
-15.2625246047974,-45.0977134704590,
-15.0837726593018,-52.7831764221191,
-17.2616004943848,-27.6208248138428,
-6.20659255981445,20.9284019470215,
13.5385398864746,57.4225311279297,
26.6341228485107,51.6208190917969,
23.4035968780518,14.3202552795410,
15.7740783691406,-7.61951684951782,
8.61153697967529,11.9025077819824,
-3.97963237762451,44.7402076721191,
-23.3240013122559,43.8512039184570,
-36.3063316345215,-0.358541488647461,
-25.8942375183105,-45.7848930358887,
3.75366020202637,-50.9526634216309,
31.6904430389404,-24.7825698852539,
43.0786781311035,-15.2979240417480,
44.4698524475098,-35.1895523071289,
45.2702713012695,-43.7368583679199,
39.9042930603027,-6.96321105957031,
19.5302314758301,49.0849266052246,
-11.2309284210205,60.7167091369629,
-36.8781280517578,16.8054733276367,
-49.3335380554199,-27.6930637359619,
-46.9953079223633,-19.1077289581299,
-32.2104682922363,29.2220859527588,
-7.42532920837402,57.2342681884766,
14.8341674804688,36.5182685852051,
18.3204040527344,-0.753198862075806,
8.44391632080078,-10.8894386291504,
4.12097787857056,11.6587104797363,
17.9593677520752,34.6109619140625,
32.5359458923340,32.0671043395996,
29.5934658050537,6.92969465255737,
18.2665252685547,-24.0627822875977,
13.9512472152710,-40.6197509765625,
16.9686183929443,-34.9896583557129,
10.1739473342896,-12.4548835754395,
-0.794891834259033,9.80329799652100,
4.02802705764771,17.3049049377441,
33.2977561950684,17.5659523010254,
60.9765739440918,21.5907974243164,
54.7661399841309,27.7465190887451,
18.4719886779785,18.8301486968994,
-24.1115550994873,-6.59633636474609,
-54.0125122070313,-18.5527534484863,
-64.2136077880859,7.23456382751465,
-48.7474555969238,44.6558151245117,
-11.0240554809570,43.9409980773926,
24.1712703704834,-3.23338174819946,
36.2185821533203,-48.1626396179199,
35.7265357971191,-39.5785408020020,
45.3181304931641,12.1584167480469,
55.4581909179688,51.2904319763184,
33.6795806884766,50.0890007019043,
-21.6685676574707,23.7584724426270,
-61.0404815673828,1.41911017894745,
-40.3187713623047,-14.1141796112061,
14.2939233779907,-24.4880180358887,
40.9188728332520,-22.2076416015625,
20.8005523681641,-4.11860942840576,
-7.05614376068115,11.4414100646973,
-16.7567920684814,8.43091773986816,
-18.4048080444336,-3.59878134727478,
-28.0020446777344,-1.93017256259918,
-32.5721359252930,14.7606964111328,
-25.6791496276855,20.5856723785400,
-29.4440383911133,-1.00298118591309,
-55.0538177490234,-35.3733825683594,
-71.2365646362305,-57.4506492614746,
-36.2064399719238,-62.5198097229004,
33.1057624816895,-48.4220886230469,
73.1366424560547,-10.8456850051880,
51.0292129516602,36.0059318542481,
5.72398185729981,60.9349555969238,
-12.9731454849243,48.7951316833496,
-7.55984258651733,26.9171867370605,
-6.23814201354981,32.5227928161621,
-17.4686679840088,56.6290016174316,
-26.5334815979004,51.2994117736816,
-22.1006507873535,1.35004556179047,
-4.67052459716797,-43.6981773376465,
18.2014980316162,-40.4953460693359,
34.7797470092773,-13.6518545150757,
30.0779571533203,-13.4980182647705,
-1.43300652503967,-40.6115760803223,
-31.3972396850586,-50.1569175720215,
-25.3952999114990,-26.8759899139404,
11.7877607345581,-3.32328796386719,
34.4332885742188,-6.30938863754273,
23.7357311248779,-10.0532617568970,
9.37120437622070,8.55356121063232,
13.2408475875855,23.9460945129395,
18.5769996643066,1.28485536575317,
8.34595870971680,-38.9554901123047,
1.56251740455627,-36.1704711914063,
25.0384235382080,14.4451227188110,
58.1937332153320,47.8719978332520,
49.8408966064453,19.2370357513428,
-1.82580602169037,-31.1671810150147,
-35.1253051757813,-46.4969978332520,
-13.1224431991577,-19.8358325958252,
24.8849411010742,5.13922595977783,
20.3774185180664,2.73623609542847,
-15.3214435577393,-11.9825458526611,
-30.2427406311035,-18.9625320434570,
-10.3403730392456,-24.0783081054688,
13.8563976287842,-30.4515724182129,
26.4966106414795,-31.3267288208008,
41.4749908447266,-25.0130252838135,
62.5590019226074,-19.5680408477783,
56.3403244018555,-13.5502223968506,
6.97689580917358,5.95961380004883,
-41.7376785278320,28.7234020233154,
-40.7695693969727,18.1631870269775,
-7.18864059448242,-29.8752651214600,
9.78746700286865,-67.3923110961914,
6.78702974319458,-51.6659507751465,
20.2252635955811,3.75105977058411,
54.1648635864258,35.2334785461426,
61.8469772338867,10.2748661041260,
25.1903915405273,-36.2494392395020,
-11.4270982742310,-55.6533241271973,
-3.39326667785645,-37.0675544738770,
23.0742683410645,-5.42497444152832,
13.9750852584839,12.7656383514404,
-23.8609580993652,5.43817949295044,
-28.4582099914551,-18.9261035919189,
12.7474803924561,-29.0643157958984,
41.7239189147949,-1.59075164794922,
11.4229345321655,41.0931015014648,
-36.5225296020508,43.9824905395508,
-35.9683990478516,-15.2809286117554,
10.8959102630615,-80.8368835449219,
53.7069358825684,-77.5645751953125,
58.7889785766602,-6.44994020462036,
43.5955657958984,52.8694877624512,
33.1178054809570,50.6697807312012,
31.0598297119141,22.1745853424072,
27.5901927947998,23.1488609313965,
29.9122333526611,43.0155029296875,
39.2800292968750,42.9216194152832,
38.8898353576660,26.4699077606201,
16.9682674407959,36.3174743652344,
-12.9356575012207,70.9731063842773,
-34.6711311340332,71.2331390380859,
-45.3777389526367,6.05743646621704,
-35.8490943908691,-59.5177345275879,
6.56549167633057,-51.9336166381836,
60.8020935058594,7.82144260406494,
82.2697296142578,35.9923057556152,
50.3008422851563,-1.46446037292480,
3.00948286056519,-50.4180374145508,
2.08929371833801,-60.8005867004395,
40.4821739196777,-49.9608688354492,
57.2649879455566,-49.0793876647949,
27.5676078796387,-47.3349685668945,
-0.727801144123077,-19.5385131835938,
8.81616973876953,10.6987905502319,
29.7337131500244,1.70414698123932,
24.0907211303711,-38.6587257385254,
10.3804626464844,-47.9210662841797,
24.9692173004150,2.01690530776978,
45.9701080322266,59.8355636596680,
15.0378408432007,58.7911033630371,
-62.2084045410156,6.75169754028320,
-95.1466369628906,-35.6902885437012,
-33.6304397583008,-33.3260574340820,
53.4039993286133,-0.896636009216309,
67.9565200805664,21.6090068817139,
9.70083045959473,13.0836219787598,
-25.5765209197998,-8.44625568389893,
7.39606237411499,-13.4289855957031,
45.7981567382813,10.7600908279419,
24.9309616088867,40.5735321044922,
-30.6582965850830,36.3270263671875,
-49.2144737243652,-10.9920959472656,
-16.8163642883301,-53.8685417175293,
11.5193910598755,-39.2770690917969,
-6.58017539978027,19.0033550262451,
-40.8050270080566,53.4401321411133,
-39.1594047546387,37.1554107666016,
-2.13049173355103,10.4789342880249,
22.1530246734619,16.4713745117188,
2.48039245605469,34.6236648559570,
-36.8684577941895,16.4200267791748,
-52.5310554504395,-31.6763153076172,
-24.5468215942383,-47.2688255310059,
18.2194995880127,-4.28030014038086,
27.8046340942383,42.4024353027344,
0.425946831703186,36.2055625915527,
-22.1368236541748,-3.60260486602783,
-7.64766979217529,-14.5118036270142,
26.9229946136475,14.0449790954590,
36.7585105895996,29.2664413452148,
12.1115798950195,1.44338226318359,
-5.40699243545532,-30.5720825195313,
15.8512773513794,-17.6684017181397,
49.9012069702148,30.1434326171875,
48.7159957885742,62.8833732604981,
19.1332397460938,52.9353599548340,
4.91827487945557,22.8530426025391,
19.6722946166992,-0.372480332851410,
27.8496646881104,-14.9276819229126,
2.30559897422791,-25.4866924285889,
-32.0784492492676,-26.6314525604248,
-31.7933883666992,-20.4950962066650,
-3.19335246086121,-20.1279716491699,
16.0737075805664,-24.4395160675049,
14.6884584426880,-20.7634868621826,
17.6061325073242,0.512983202934265,
29.2035827636719,28.2342700958252,
15.4901075363159,43.5884590148926,
-35.2183570861816,39.8427085876465,
-73.0587234497070,18.5813484191895,
-49.4647636413574,-18.4333820343018,
9.97125911712647,-57.3770523071289,
32.8487472534180,-64.0701904296875,
1.95587325096130,-20.7468986511230,
-25.6385459899902,32.0016708374023,
-5.40089988708496,37.2034721374512,
31.9121646881104,-8.63786888122559,
34.0883026123047,-45.0760040283203,
7.87781524658203,-25.6756973266602,
1.77899050712585,25.0894393920898,
24.1806182861328,47.0604171752930,
29.9205627441406,22.7053642272949,
-3.97715735435486,-13.5221691131592,
-38.0790252685547,-25.2646522521973,
-25.3122272491455,-14.1851596832275,
19.9671478271484,-5.44500350952148,
48.5791435241699,-9.25780677795410,
43.5465393066406,-22.8715496063232,
32.3775901794434,-34.5573577880859,
41.8081665039063,-36.3071517944336,
54.2949562072754,-25.0693225860596,
42.0284271240234,-6.30636453628540,
12.9132823944092,3.89129328727722,
-1.94672703742981,-1.08133900165558,
9.72838020324707,-13.5182409286499,
27.3609580993652,-23.0464286804199,
24.7681503295898,-25.7278995513916,
3.05308938026428,-21.2197761535645,
-12.8374061584473,-12.1522350311279,
-4.06570291519165,3.66772508621216,
17.4466361999512,20.0331153869629,
25.4532737731934,29.4764213562012,
13.6740217208862,33.9446029663086,
-4.59444379806519,38.8805885314941,
-16.0969696044922,40.3503227233887,
-23.4735660552979,26.3535633087158,
-37.5514106750488,-2.31414747238159,
-55.2094306945801,-27.7964458465576,
-58.7090263366699,-26.7678413391113,
-39.7205276489258,-5.36064243316650,
-12.7498292922974,11.9546318054199,
7.11928176879883,11.9602203369141,
18.7744159698486,8.76781082153320,
28.2451438903809,20.3475074768066,
29.3092765808105,40.5774345397949,
11.7339916229248,42.3378334045410,
-17.9276561737061,19.0785598754883,
-32.9040145874023,-3.19286870956421,
-19.2197704315186,-0.174564719200134,
2.47038698196411,15.2247934341431,
-4.11835813522339,9.98769092559815,
-41.1075363159180,-23.1818637847900,
-69.1964263916016,-52.0415153503418,
-57.3988990783691,-43.0157089233398,
-19.7640991210938,-1.05722117424011,
8.75716400146484,29.9680423736572,
11.1951236724854,21.9445552825928,
4.27292871475220,-5.13675498962402,
-0.0179711580276489,-12.0642623901367,
-7.02999353408814,11.0394964218140,
-17.7567749023438,34.9588394165039,
-13.8033351898193,30.7327327728272,
4.81945991516113,7.95799446105957,
8.41749000549316,-1.37792003154755,
-24.2735767364502,4.67816114425659,
-58.9290809631348,-3.25569868087769,
-45.5636024475098,-35.4208641052246,
7.01761722564697,-53.8200378417969,
37.4686470031738,-29.1311187744141,
16.7567481994629,16.8616828918457,
-8.11503601074219,31.8244953155518,
7.45564746856689,4.97183465957642,
40.2265014648438,-20.6238689422607,
28.1839561462402,-14.6053962707520,
-23.0274353027344,0.504255890846252,
-43.1723518371582,-3.31949949264526,
-2.02637457847595,-14.5779905319214,
51.1456031799316,-5.90996646881104,
62.1749534606934,13.8051128387451,
44.5505218505859,11.2037029266357,
39.9906616210938,-11.0408267974854,
44.0473518371582,-6.69519138336182,
26.2691116333008,38.2209129333496,
-8.44963932037354,82.1898956298828,
-25.9365844726563,80.3605422973633,
-19.3109645843506,44.9030876159668,
-26.1480598449707,22.1422176361084,
-54.3522148132324,30.4422702789307,
-56.0672836303711,44.3962326049805,
-0.451127648353577,36.2152748107910,
63.6252822875977,12.4570846557617,
67.5528869628906,-6.47479534149170,
12.1677083969116,-11.7260780334473,
-37.3451995849609,-2.84318447113037,
-39.0358963012695,13.9388027191162,
-9.42632484436035,18.8798885345459,
15.5120296478271,-5.22940826416016,
25.1850528717041,-42.9773330688477,
25.9604816436768,-58.2850494384766,
11.5771665573120,-34.6383590698242,
-21.3444442749023,2.59238934516907,
-49.1667213439941,21.9182605743408,
-49.0657730102539,20.1425704956055,
-34.6552009582520,21.1586399078369,
-32.0307769775391,28.9990043640137,
-42.4348602294922,28.2219257354736,
-38.7073554992676,18.1856899261475,
-12.3055305480957,17.5074710845947,
18.1011238098145,26.5019664764404,
31.2588787078857,21.4539108276367,
29.5730876922607,-7.27116966247559,
25.3556232452393,-31.1686477661133,
17.2393722534180,-13.8088932037354,
-0.227819800376892,31.7885704040527,
-15.1435108184814,55.5023689270020,
-7.96608352661133,37.4890213012695,
12.4774179458618,8.64291381835938,
16.2017612457275,2.21503782272339,
-8.13126373291016,10.8739852905273,
-33.3526458740234,1.94462251663208,
-30.8729057312012,-28.1688632965088,
-8.25003814697266,-46.7015075683594,
-3.16206526756287,-31.3135375976563,
-28.0388374328613,-4.37808609008789,
-53.8739318847656,3.86325287818909,
-38.8623580932617,-1.95392525196075,
13.3233127593994,9.16036033630371,
54.1500968933106,42.8535041809082,
44.9696388244629,61.6304969787598,
-6.15710735321045,31.9574203491211,
-51.1916580200195,-19.6213493347168,
-57.2876167297363,-36.6592330932617,
-34.0565452575684,-1.67589688301086,
-8.89466667175293,37.8632392883301,
3.74529123306274,32.0669479370117,
12.2637662887573,-7.30135202407837,
16.6282997131348,-29.0092582702637,
6.17039632797241,-8.37007045745850,
-19.2616157531738,23.1278495788574,
-39.3666419982910,21.7975311279297,
-34.6068115234375,-11.7467432022095,
-11.4334230422974,-39.4454727172852,
0.377161055803299,-35.1009902954102,
-16.9609737396240,-11.3084821701050,
-44.3690986633301,1.44982719421387,
-53.7273025512695,-12.9520778656006,
-34.4437522888184,-45.7309455871582,
2.09117650985718,-68.6513900756836,
31.6818714141846,-59.4391098022461,
45.6992645263672,-13.7938480377197,
48.4944458007813,43.4553146362305,
43.8018035888672,70.7269821166992,
32.4866104125977,46.5917778015137,
16.7144432067871,1.98124790191650,
9.09636592864990,-15.5220775604248,
20.1713008880615,10.6510162353516,
41.1406822204590,41.9174003601074,
44.1104202270508,34.4393348693848,
12.1563634872437,-3.58525943756104,
-30.7398681640625,-24.0711250305176,
-48.2433166503906,-4.59635925292969,
-29.8921127319336,25.1787319183350,
-6.40454292297363,25.4276638031006,
-10.3942871093750,2.54433059692383,
-39.8458480834961,-8.25283527374268,
-57.7202682495117,5.17253780364990,
-45.0657119750977,9.56806182861328,
-16.2012348175049,-16.3162841796875,
3.14204597473145,-54.7154045104981,
2.55914878845215,-65.9486160278320,
0.644063115119934,-41.8315544128418,
9.95527839660645,-16.3433170318604,
18.7459545135498,-12.2579898834229,
4.75444364547730,-17.0097885131836,
-30.1011371612549,-9.26966094970703,
-51.8430709838867,9.89588451385498,
-36.4411773681641,16.7629623413086,
-1.59344291687012,2.87933135032654,
17.5367908477783,-7.26466131210327,
14.1919574737549,5.29126548767090,
17.0963001251221,29.3518238067627,
41.1670951843262,42.3271484375000,
59.1397018432617,41.3587150573731,
36.7994956970215,42.7096405029297,
-13.4539299011230,42.2704849243164,
-48.7771873474121,17.8188076019287,
-50.1522521972656,-31.9079132080078,
-34.1208724975586,-61.9480209350586,
-16.9595642089844,-36.4931564331055,
-3.56183910369873,20.2507972717285,
-0.117945656180382,43.6943359375000,
-16.1491317749023,9.98167705535889,
-37.5600051879883,-39.8649444580078,
-29.4642353057861,-58.4330291748047,
12.6473989486694,-42.6344985961914,
47.0374984741211,-17.0339145660400,
36.0281562805176,13.0306148529053,
5.08065319061279,48.5486259460449,
1.53293514251709,66.8986511230469,
20.2685775756836,42.8896636962891,
8.90736770629883,-10.0521240234375,
-41.3013572692871,-47.4027824401856,
-68.0882263183594,-46.7737197875977,
-30.8978385925293,-31.4983501434326,
30.0813827514648,-27.6698417663574,
46.8898200988770,-29.6313953399658,
13.8046131134033,-16.4247283935547,
-13.9770021438599,4.94839525222778,
-3.41621613502502,16.5853862762451,
16.1048469543457,25.0604953765869,
8.05705070495606,39.3096046447754,
-25.2431144714355,41.6317329406738,
-53.9838523864746,13.5644378662109,
-62.8967590332031,-32.8248481750488,
-51.1931762695313,-55.3555068969727,
-16.2545127868652,-36.2898712158203,
26.4748401641846,-5.61591482162476,
40.9930686950684,12.4614572525024,
13.4767742156982,23.5636749267578,
-25.4181213378906,38.2219696044922,
-36.8325157165527,31.6527118682861,
-21.6999874114990,-18.7774353027344,
-10.6327123641968,-69.2530059814453,
-18.7549571990967,-57.2560310363770,
-26.3301982879639,8.47141647338867,
-21.4061412811279,47.1746635437012,
-20.9941139221191,12.7989082336426,
-26.9519844055176,-45.4020423889160,
-18.5385837554932,-52.1690521240234,
8.08719539642334,-3.81536722183228,
15.6218347549438,40.1393165588379,
-15.8777256011963,47.2495651245117,
-47.7024650573731,38.4715423583984,
-27.1044254302979,34.3441047668457,
28.1973571777344,21.3250007629395,
46.3889160156250,-1.11715257167816,
5.30890178680420,-4.02092027664185,
-37.5027618408203,23.0223960876465,
-26.0893821716309,44.3507156372070,
15.4481115341187,27.8442802429199,
18.0036888122559,-1.83796906471252,
-28.7359695434570,-0.440991133451462,
-69.0890731811523,18.9201583862305,
-67.5535430908203,7.87457418441773,
-42.1369476318359,-41.6334915161133,
-22.9323921203613,-76.5391540527344,
-10.8605813980103,-55.4537086486816,
9.14845275878906,-9.87023925781250,
33.5182342529297,7.12301063537598,
45.0325279235840,-0.523872613906860,
36.9171791076660,3.56125855445862,
16.1256885528564,27.6860160827637,
-4.30300426483154,39.0317077636719,
-12.6720161437988,19.5259723663330,
2.23178434371948,-4.68538808822632,
35.2398452758789,-0.931720733642578,
46.5989227294922,28.3206100463867,
9.42510890960693,48.5360717773438,
-46.0743942260742,34.0930290222168,
-55.1665306091309,-5.80507373809814,
-5.58408498764038,-41.5127067565918,
50.4409561157227,-41.7420387268066,
55.1580390930176,-0.290122747421265,
20.9310359954834,55.2073211669922,
-2.40812492370605,72.2911300659180,
-0.920602679252625,39.2305755615234,
-5.19826602935791,-7.88701820373535,
-33.8073348999023,-24.1502532958984,
-56.2361640930176,-5.28633880615234,
-44.3649101257324,16.4429721832275,
-17.3069076538086,22.7410469055176,
-15.2153053283691,25.0035552978516,
-42.5183753967285,34.6486663818359,
-65.0927200317383,38.4779777526856,
-60.8546981811523,18.6882152557373,
-42.0026283264160,-12.1566104888916,
-31.7063617706299,-28.6668148040772,
-32.4313087463379,-31.4396476745605,
-29.7078781127930,-41.9195289611816,
-13.5988569259644,-63.7866096496582,
9.71500396728516,-72.0176544189453,
31.4722518920898,-47.3289833068848,
36.5423088073731,-5.72928905487061,
14.0707092285156,24.0164566040039,
-17.9742317199707,26.1143169403076,
-27.1084384918213,11.8540563583374,
-1.15614497661591,-1.04263210296631,
27.4809761047363,-0.874522328376770,
27.7522563934326,15.8629360198975,
11.4804801940918,39.8802833557129,
16.2415313720703,50.1682167053223,
44.8537902832031,33.5299797058106,
54.8271789550781,10.2021913528442,
20.1909465789795,12.0135965347290,
-18.8370609283447,36.8271980285645,
-14.1493215560913,50.4891319274902,
18.5357761383057,32.2172431945801,
22.4687385559082,2.71884393692017,
-21.4857540130615,-6.41111564636231,
-67.8607406616211,11.0382499694824,
-69.3816223144531,27.7567825317383,
-36.3737335205078,27.2711982727051,
-8.52226638793945,18.7346553802490,
-2.05323696136475,8.92088699340820,
-5.96367216110230,0.997044801712036,
-13.0262775421143,4.78878307342529,
-26.0882644653320,31.2236480712891,
-38.4603576660156,66.1641082763672,
-30.4737968444824,71.1725082397461,
-4.78946495056152,30.4023838043213,
8.98027896881104,-14.1497659683228,
-4.93549489974976,-14.1109333038330,
-25.9615402221680,20.8401145935059,
-28.3684043884277,33.2697219848633,
-13.7059555053711,-2.72322893142700,
-0.671641945838928,-42.4312362670898,
0.0777193605899811,-27.6532154083252,
-3.97389054298401,30.4102439880371,
0.323375880718231,65.5762100219727,
7.18884372711182,40.8359069824219,
14.0936794281006,-9.82412815093994,
17.1373863220215,-26.7376651763916,
9.19715499877930,4.46025276184082,
-12.4535150527954,44.9430694580078,
-27.0241889953613,50.8531341552734,
-12.0868101119995,21.7309513092041,
28.3930549621582,-8.67516040802002,
52.4028434753418,-10.6327304840088,
35.0134811401367,9.51937389373779,
2.53417110443115,21.0837535858154,
-3.66791415214539,7.85296058654785,
15.4842996597290,-18.4562492370605,
15.7747840881348,-30.4216327667236,
-23.7024631500244,-22.2102661132813,
-67.5151901245117,-14.0877008438110,
-66.3639602661133,-17.1165237426758,
-27.9775905609131,-17.8103981018066,
-4.83759880065918,-2.50170946121216,
-24.1059207916260,19.1319923400879,
-55.0889282226563,21.8932533264160,
-50.2299194335938,0.217313885688782,
-2.67796611785889,-19.3068332672119,
44.7099227905273,-10.6845617294312,
49.6542015075684,20.5561218261719,
12.9317407608032,49.6050262451172,
-25.4970149993897,58.7619056701660,
-31.6224803924561,50.0555076599121,
-9.55963706970215,33.9406967163086,
4.96602773666382,16.8669071197510,
-15.4553737640381,4.24041652679443,
-51.4870567321777,-3.65640044212341,
-56.8220062255859,-10.2405242919922,
-18.8213214874268,-17.6590709686279,
18.9753341674805,-20.8255004882813,
12.2011699676514,-15.3516893386841,
-30.8339233398438,-5.72752952575684,
-57.0291976928711,-5.49683856964111,
-44.3062400817871,-15.0867738723755,
-22.4469070434570,-19.9663829803467,
-26.8129901885986,-9.12399482727051,
-37.5536766052246,7.30748319625855,
-13.9724102020264,8.07819747924805,
35.0527992248535,-3.98494005203247,
57.4635124206543,-2.45423698425293,
27.0008468627930,20.5862216949463,
-18.2807178497314,47.2191734313965,
-22.8671779632568,48.4516410827637,
12.1671504974365,27.9432487487793,
37.7959632873535,15.7595939636230,
25.4555377960205,28.5287971496582,
-10.0960531234741,48.0217819213867,
-35.6483802795410,53.1521148681641,
-40.6350479125977,37.1489715576172,
-35.2495422363281,9.30013847351074,
-26.5226535797119,-22.2265148162842,
-11.3988103866577,-48.1888198852539,
5.24654054641724,-51.4292449951172,
11.1741828918457,-25.4656009674072,
0.558194339275360,4.22610330581665,
-10.1635217666626,-1.91016149520874,
-2.99070477485657,-43.7624053955078,
19.5206985473633,-71.9617614746094,
34.9489402770996,-45.5264892578125,
21.6660995483398,11.3695735931396,
-9.28371810913086,31.9928512573242,
-27.8116226196289,-7.54863834381104,
-24.1974105834961,-61.8786697387695,
-13.7906227111816,-70.9501037597656,
-10.3156118392944,-33.3984069824219,
-5.03996562957764,7.93777751922607,
13.2846889495850,19.8093357086182,
29.3528175354004,17.2570362091064,
16.7533798217773,25.8852214813232,
-21.3933811187744,43.8219947814941,
-47.4947357177734,52.1523513793945,
-39.8236503601074,39.5719718933106,
-21.4776916503906,17.8696632385254,
-24.6516304016113,2.52652406692505,
-39.1818428039551,0.484949588775635,
-29.3039150238037,10.5574893951416,
10.1036472320557,26.6686992645264,
40.8237304687500,33.1365318298340,
27.5482406616211,28.3550014495850,
-9.49325656890869,21.5884933471680,
-21.2699432373047,21.9693756103516,
6.51981544494629,29.3903255462647,
38.2451438903809,27.1750869750977,
39.7625427246094,8.36339378356934,
17.6162242889404,-14.1972465515137,
0.678098082542419,-23.4366874694824,
0.447018802165985,-16.3594169616699,
3.52756738662720,-2.31432604789734,
5.90195798873901,6.64454698562622,
18.2646636962891,0.368238985538483,
35.9016075134277,-13.9658737182617,
32.5411605834961,-16.2437267303467,
-4.79924726486206,11.3480453491211,
-42.9062194824219,50.2637710571289,
-38.2232055664063,60.0444488525391,
7.03637886047363,22.3592376708984,
40.2341842651367,-24.0459728240967,
28.4142360687256,-29.4126205444336,
-5.96806097030640,3.45012474060059,
-20.0036983489990,23.1825904846191,
-5.45621395111084,-1.89137411117554,
15.5740671157837,-38.0052375793457,
23.3812980651855,-42.1045074462891,
23.6737709045410,-18.6833572387695,
22.2216606140137,-3.67850303649902,
15.3555021286011,-12.5195703506470,
2.07377862930298,-22.8917655944824,
-6.87747907638550,-20.1625576019287,
-8.75031471252441,-20.4029006958008,
-9.37993335723877,-36.3114585876465,
-7.68228340148926,-53.8196182250977,
8.30793952941895,-52.0736351013184,
35.5132064819336,-35.4379997253418,
49.5864486694336,-21.5109157562256,
36.0136566162109,-12.5588598251343,
13.5599937438965,9.93301773071289,
12.4507598876953,41.0083007812500,
29.8013496398926,51.7251892089844,
36.1476631164551,25.1874027252197,
22.1308860778809,-19.6702518463135,
13.1543149948120,-46.5496978759766,
28.4630603790283,-34.5715599060059,
51.3880119323731,-0.0268039703369141,
54.8911399841309,24.3610439300537,
42.2615661621094,17.5103454589844,
34.2640113830566,-11.1004953384399,
33.3603553771973,-34.1659545898438,
20.7227725982666,-26.1887855529785,
-9.84293365478516,1.77441930770874,
-33.8444976806641,11.9593992233276,
-27.2096214294434,-13.9791193008423,
1.75985383987427,-45.6888313293457,
25.5016613006592,-43.5542984008789,
27.8562602996826,-9.65227127075195,
13.0594253540039,12.6028633117676,
-4.34156560897827,1.08473670482636,
-16.6019248962402,-18.7556152343750,
-17.7410812377930,-13.3355684280396,
-8.06953239440918,5.47384548187256,
0.983284056186676,0.430351972579956,
-5.63874149322510,-26.8710231781006,
-23.3850517272949,-33.1713104248047,
-34.0378036499023,2.97606611251831,
-20.8075351715088,42.1487159729004,
4.59576272964478,34.3598785400391,
18.0121326446533,-15.0018205642700,
4.13714408874512,-47.4221954345703,
-17.3203468322754,-31.8439979553223,
-17.9396667480469,7.06748819351196,
7.98383045196533,24.6734600067139,
39.1269340515137,10.9556264877319,
42.9218711853027,-8.20803642272949,
10.9042034149170,-8.71076107025147,
-24.4584121704102,6.80690383911133,
-25.6344738006592,22.3956260681152,
4.97518157958984,24.4899272918701,
28.3855857849121,6.52447509765625,
23.6804828643799,-20.9243774414063,
13.8808393478394,-33.3397064208984,
28.4847106933594,-18.0615653991699,
50.9372138977051,10.2584562301636,
31.1630058288574,32.9397506713867,
-36.7282714843750,45.7967834472656,
-83.4016571044922,52.2235908508301,
-49.0955200195313,47.8459472656250,
24.3520832061768,22.5599994659424,
44.6241569519043,-10.2843618392944,
-9.03743743896484,-18.9125003814697,
-57.0800056457520,1.82011938095093,
-33.7663116455078,15.6135511398315,
19.4430866241455,-2.71229171752930,
21.6028156280518,-23.5166282653809,
-22.4748058319092,-10.4797925949097,
-33.0703125000000,20.4686260223389,
15.8762502670288,22.7306556701660,
51.4920616149902,-7.88245582580566,
13.4660282135010,-27.1222076416016,
-51.1236152648926,-10.1406669616699,
-63.1613235473633,13.3020935058594,
-24.8401165008545,6.49812412261963,
-5.16376781463623,-19.6338119506836,
-28.6705570220947,-30.8666496276855,
-49.2704238891602,-28.6304225921631,
-37.2002868652344,-31.8939399719238,
-20.5499019622803,-28.9966621398926,
-24.1236000061035,5.30697822570801,
-26.8864288330078,49.3186340332031,
-2.32560253143311,50.9690856933594,
20.9507102966309,5.02368879318237,
7.08304595947266,-28.3203945159912,
-20.0152854919434,-10.2571115493774,
-13.3690071105957,27.6469993591309,
17.3208427429199,29.8517723083496,
21.8560714721680,-1.59077334403992,
-5.49151659011841,-19.2533645629883,
-17.3054809570313,-10.9585990905762,
8.41523170471191,-10.3768186569214,
33.8338317871094,-21.7933826446533,
14.6465568542480,-8.31094551086426,
-30.4571743011475,34.5684890747070,
-51.6649055480957,53.7884712219238,
-43.9600296020508,18.5970706939697,
-40.1290168762207,-31.6669998168945,
-43.1526260375977,-41.7887573242188,
-31.8683376312256,-27.3301391601563,
-5.53194093704224,-37.3718872070313,
10.6610641479492,-69.3752212524414,
8.58308792114258,-62.9799652099609,
4.33422565460205,-6.89322519302368,
-0.0530546903610230,29.9515438079834,
-14.6892223358154,3.25542688369751,
-33.9814834594727,-36.6624870300293,
-27.9652328491211,-23.2222747802734,
7.52556419372559,22.1841640472412,
25.4677429199219,30.5400466918945,
-11.1164045333862,-3.02252435684204,
-62.9937438964844,-15.6657047271729,
-58.4633865356445,17.9767761230469,
3.70823764801025,47.6709671020508,
51.4358978271484,29.3247470855713,
45.2646751403809,-3.90603971481323,
17.2418098449707,6.46359634399414,
4.14024591445923,46.8380508422852,
-4.28232955932617,56.6832046508789,
-34.7156372070313,17.9850788116455,
-69.2805328369141,-26.0820827484131,
-66.1938171386719,-44.1225013732910,
-27.4793357849121,-36.4711112976074,
-0.131380796432495,-15.9654407501221,
-2.79540753364563,10.1389360427856,
-7.32869482040405,23.9824275970459,
5.84784030914307,6.66749620437622,
14.2653236389160,-25.2030868530273,
5.85030746459961,-25.0405941009522,
5.68860292434692,17.4198055267334,
30.7393779754639,49.6726837158203,
43.1612434387207,23.5937938690186,
5.02009773254395,-26.7603130340576,
-51.5777587890625,-30.2568244934082,
-61.0913734436035,13.1635904312134,
-15.3098754882813,33.1984138488770,
17.2545833587647,-9.17450046539307,
-6.33859252929688,-69.4428176879883,
-42.3392181396484,-80.2433700561523,
-31.3811607360840,-35.3452873229981,
4.22157526016235,10.9954652786255,
7.19696617126465,19.8935527801514,
-24.3960208892822,-2.09704709053040,
-30.3692283630371,-24.2205600738525,
14.8948669433594,-25.5613498687744,
61.6124992370606,-6.70322465896606,
53.9720993041992,23.3812332153320,
3.03118610382080,43.6105918884277,
-37.4478607177734,36.2170524597168,
-43.8969383239746,7.14305210113525,
-34.0654449462891,-17.2754955291748,
-23.1223754882813,-27.0491905212402,
-4.76002550125122,-26.5914516448975,
16.0391731262207,-19.5274009704590,
16.1328086853027,-7.59378242492676,
-10.1840400695801,-1.22793662548065,
-39.5372428894043,-9.17580127716065,
-48.2256622314453,-27.6619510650635,
-36.4443740844727,-24.0863304138184,
-19.3759880065918,18.8765296936035,
-7.22615003585815,61.4806938171387,
-0.296406924724579,52.7029724121094,
0.677284777164459,0.619458675384522,
-4.16992092132568,-35.2267990112305,
-6.96911859512329,-23.1105651855469,
1.94156622886658,-2.10746407508850,
13.2047643661499,-22.0567378997803,
13.2628068923950,-60.9046287536621,
7.92921733856201,-60.9934997558594,
11.0335350036621,-18.1220970153809,
21.5988273620605,5.32769012451172,
24.5473918914795,-27.3161640167236,
15.4913997650146,-66.5811996459961,
10.1733522415161,-41.4114685058594,
16.7821331024170,32.2945098876953,
28.2935581207275,70.5994949340820,
27.6379470825195,33.5574722290039,
16.7936611175537,-21.5892505645752,
5.46423864364624,-18.7966518402100,
-4.71830320358276,37.1923637390137,
-16.1098594665527,78.3487472534180,
-21.1212768554688,58.3432121276856,
-8.56875228881836,1.69514441490173,
13.0685815811157,-31.5179233551025,
18.1456050872803,-21.6809120178223,
-2.77863454818726,3.67801856994629,
-28.3434276580811,9.29918003082275,
-39.8784751892090,-11.3869647979736,
-40.9563751220703,-37.3615837097168,
-47.1713638305664,-44.9331207275391,
-57.6049652099609,-27.9015216827393,
-52.6952514648438,-5.60797214508057,
-27.6522312164307,9.71492481231690,
-2.39384365081787,17.2739830017090,
9.65369987487793,17.8116302490234,
23.1408100128174,9.29094982147217,
46.5886650085449,-3.60612154006958,
65.5062179565430,-4.69768095016480,
59.0299758911133,17.5601062774658,
33.5487632751465,51.6367263793945,
12.2005548477173,60.3757438659668,
-1.34512460231781,29.8701820373535,
-24.9074020385742,-12.9025945663452,
-53.4118957519531,-35.4995117187500,
-52.2672691345215,-39.7198295593262,
-11.6137733459473,-45.8630065917969,
25.1715641021729,-56.4143600463867,
12.3992786407471,-54.4173393249512,
-29.0615425109863,-36.7321815490723,
-31.5914497375488,-26.3474388122559,
18.5767707824707,-33.9303054809570,
63.9839630126953,-35.8826026916504,
56.3515396118164,-5.77318954467773,
17.9563713073730,38.9663734436035,
4.79976940155029,57.7312240600586,
22.5488262176514,44.5582008361816,
29.0422554016113,33.7745018005371,
0.803927361965179,42.6068801879883,
-29.1297435760498,43.2524871826172,
-24.4082794189453,3.78317546844482,
7.98238849639893,-47.3017768859863,
31.2931842803955,-54.8882675170898,
23.9924335479736,-8.83066368103027,
-3.63778018951416,41.7243766784668,
-30.9218654632568,51.8860588073731,
-34.2642250061035,30.2541122436523,
-8.96361160278320,13.7243347167969,
26.4306221008301,14.2955465316772,
42.3794021606445,13.3096876144409,
24.3550834655762,-1.64654254913330,
-9.90040969848633,-14.9310932159424,
-24.4026012420654,-17.7824287414551,
-12.2964468002319,-21.6955814361572,
6.30542325973511,-40.4016876220703,
12.8258075714111,-64.6626434326172,
9.90238285064697,-65.3781356811523,
3.49339866638184,-35.5363159179688,
-6.26629972457886,0.539913594722748,
-14.8123130798340,8.22595596313477,
-9.94139671325684,-12.4605350494385,
16.0370197296143,-22.3518905639648,
42.8415908813477,1.73748946189880,
40.3620986938477,39.0665016174316,
6.98277950286865,46.5583267211914,
-20.3905143737793,12.3245801925659,
-12.1530036926270,-33.3042984008789,
19.5709915161133,-57.0694923400879,
34.4218864440918,-57.3424110412598,
20.7827873229980,-46.4097328186035,
4.41329908370972,-24.2095184326172,
10.2130165100098,10.3791618347168,
27.8172836303711,37.6430397033691,
30.5495662689209,30.7486228942871,
16.7604198455811,3.35102653503418,
9.73410224914551,-5.82821607589722,
21.8470420837402,16.7278118133545,
36.8279991149902,38.4290847778320,
39.3720626831055,30.2833557128906,
34.7185783386231,7.90234470367432,
39.6665344238281,5.04556179046631,
46.3265533447266,16.7447299957275,
38.0192070007324,16.7481708526611,
18.6351127624512,2.09290218353272,
8.89391803741455,-0.0713315606117249,
20.3793888092041,16.2659072875977,
32.4237747192383,17.0719165802002,
23.6801071166992,-10.5215148925781,
4.04077196121216,-35.0420303344727,
0.718028247356415,-16.9732799530029,
21.4473171234131,26.2490863800049,
40.5754356384277,34.9470329284668,
36.9943542480469,-5.83750438690186,
20.3177490234375,-44.4294013977051,
18.6545047760010,-30.5237827301025,
42.5200576782227,22.1454086303711,
70.6371612548828,52.8964004516602,
65.2804336547852,34.7623748779297,
20.9687995910645,4.66535139083862,
-30.2376823425293,2.79942035675049,
-57.5553169250488,16.4773559570313,
-57.6110076904297,5.21015691757202,
-46.0573577880859,-37.0843200683594,
-29.4616565704346,-61.3357849121094,
-2.62527418136597,-30.3788013458252,
29.4565277099609,28.7137966156006,
36.7953147888184,55.3432235717773,
10.0502891540527,31.1474876403809,
-15.1902866363525,-3.11398267745972,
-3.10751891136169,-3.94322776794434,
25.3051300048828,26.5336284637451,
16.5537300109863,51.5632781982422,
-35.5909385681152,50.1620750427246,
-66.5790786743164,25.7138023376465,
-32.1828346252441,-5.04498815536499,
27.0187053680420,-18.5360260009766,
34.7213745117188,-0.902193009853363,
-12.9140539169312,39.1461257934570,
-45.6947135925293,59.8948554992676,
-14.5255365371704,35.4173049926758,
42.2718887329102,-4.60248088836670,
57.9437332153320,-6.75550746917725,
22.3804397583008,26.0675392150879,
-20.4341735839844,37.6541252136231,
-30.1518077850342,-1.00887846946716,
-12.1210823059082,-47.5252799987793,
10.2442111968994,-37.5680122375488,
19.1714687347412,19.8335628509522,
8.67716121673584,52.5785636901856,
-14.1823444366455,25.8089370727539,
-27.9246025085449,-25.3385143280029,
-17.1444244384766,-52.0470733642578,
9.59884548187256,-47.2750358581543,
29.6524639129639,-35.2586212158203,
28.9235248565674,-28.6306571960449,
21.1964969635010,-22.1697139739990,
27.2610244750977,-19.3560256958008,
42.8208656311035,-18.6739101409912,
54.0812873840332,-5.41928100585938,
57.4408569335938,28.1138229370117,
47.3737106323242,56.8168754577637,
19.3192081451416,44.1252899169922,
-19.7241668701172,-7.18509292602539,
-49.1650733947754,-41.5286483764648,
-50.3634071350098,-14.1847457885742,
-33.3878898620606,43.9513816833496,
-23.7278156280518,72.0669250488281,
-23.0538635253906,48.1778450012207,
-10.7832307815552,6.24752330780029,
14.3139209747314,-5.65659046173096,
19.3527603149414,21.3224887847900,
-16.6112442016602,49.7495307922363,
-54.9101257324219,43.8258247375488,
-41.4858093261719,2.03226208686829,
15.3976831436157,-34.5583648681641,
51.6104736328125,-27.5669593811035,
27.5051002502441,16.0503768920898,
-24.1771106719971,40.9316978454590,
-43.3654098510742,2.05657243728638,
-18.9363899230957,-70.3057403564453,
16.5934944152832,-96.9619140625000,
37.1403236389160,-48.5234222412109,
43.5581436157227,16.2505798339844,
38.5623588562012,33.3366966247559,
13.4323835372925,6.74531793594360,
-14.4343147277832,-10.4369087219238,
-12.4368619918823,5.60247087478638,
20.9214744567871,21.3461894989014,
40.4086875915527,17.6447315216064,
14.2417507171631,22.9434032440186,
-32.3841514587402,52.6289215087891,
-53.8577880859375,66.8935699462891,
-40.9280853271484,24.3183574676514,
-22.6132774353027,-44.5787200927734,
-14.0011234283447,-69.8138351440430,
1.68126082420349,-39.3729362487793,
28.8051929473877,-14.3602266311646,
39.1704025268555,-32.6814041137695,
27.7323989868164,-53.9456901550293,
23.7572689056397,-33.1463813781738,
42.4896278381348,11.8232498168945,
54.6762428283691,23.3755722045898,
30.7047672271729,-8.13109493255615,
-2.66246914863586,-29.0025043487549,
2.46257042884827,-7.63937854766846,
35.3812599182129,24.8993415832520,
42.1522750854492,32.3183975219727,
5.59260749816895,20.4689826965332,
-28.5382595062256,14.5105743408203,
-17.4581356048584,18.4537849426270,
6.72963285446167,18.4393768310547,
-6.44232559204102,7.23207759857178,
-48.0037956237793,-9.25572109222412,
-66.6084899902344,-17.0733203887939,
-44.7558860778809,-14.2876319885254,
-12.8199119567871,0.105739414691925,
5.33396720886231,10.6651172637939,
14.5950632095337,-5.09906959533691,
29.7447090148926,-51.4359893798828,
43.5264663696289,-81.7252044677734,
50.2924728393555,-49.6878204345703,
52.8719291687012,22.1109371185303,
49.6599540710449,57.4216232299805,
20.6760902404785,28.0836601257324,
-31.8650321960449,-15.4499578475952,
-62.8209419250488,-15.9792079925537,
-31.9007129669189,10.7009267807007,
24.8200912475586,6.11882781982422,
38.3707580566406,-36.3878173828125,
0.313644886016846,-65.5432891845703,
-27.9959831237793,-54.4767494201660,
-0.830251693725586,-39.0347557067871,
51.2864074707031,-47.8618812561035,
63.5007972717285,-48.3976974487305,
26.8858261108398,-2.83890008926392,
-14.8556909561157,63.2748718261719,
-30.4675540924072,88.2973327636719,
-28.9642639160156,60.6816749572754,
-27.5631370544434,33.8878669738770,
-23.5811653137207,38.9410400390625,
-16.3044166564941,49.7870101928711,
-17.7962207794189,30.8541793823242,
-30.1523647308350,-7.46430444717407,
-28.8303947448730,-26.6362838745117,
1.33037281036377,-22.4835128784180,
38.4575653076172,-22.3042888641357,
47.9462699890137,-26.0063591003418,
23.3515644073486,-8.45456504821777,
-9.73529148101807,26.9488048553467,
-21.9288272857666,48.7948532104492,
-14.5445365905762,31.4157638549805,
-5.32316780090332,-2.01650619506836,
-0.185214832425118,-18.4667968750000,
-0.352320343255997,-10.9073476791382,
2.33252263069153,5.70669651031494,
14.6693658828735,15.5990352630615,
34.0672149658203,20.4824790954590,
44.1341476440430,11.2581110000610,
26.6317920684814,-12.1968736648560,
-9.31861305236816,-23.2085151672363,
-34.6527519226074,5.08454084396362,
-38.0677375793457,48.7461738586426,
-35.4921188354492,53.5957603454590,
-45.8023223876953,2.99312877655029,
-62.1237335205078,-57.9067039489746,
-56.1722183227539,-80.0444107055664,
-17.8185672760010,-61.9190025329590,
32.1312065124512,-30.4963378906250,
65.9289093017578,1.30158257484436,
69.0999526977539,39.6341018676758,
41.9245948791504,64.1904602050781,
0.298494815826416,43.1188430786133,
-25.4844646453857,-6.99663448333740,
-13.7677154541016,-27.3796634674072,
16.8185081481934,1.72267961502075,
20.9274692535400,34.9154930114746,
-19.6857547760010,24.3626899719238,
-65.2805023193359,-9.95896530151367,
-65.7502288818359,-18.9003372192383,
-23.2554569244385,-2.86427330970764,
8.57945537567139,1.56825065612793,
2.23059678077698,-11.9973545074463,
-17.0769081115723,-6.60831212997437,
-7.99975824356079,32.6742858886719,
20.2324085235596,55.4938430786133,
29.8892879486084,28.1063461303711,
14.7819366455078,-11.6361417770386,
0.356697380542755,-8.15441131591797,
9.18003273010254,31.4931316375732,
26.4646339416504,44.3291091918945,
30.2735061645508,10.5122966766357,
24.3069858551025,-29.5859909057617,
24.6301593780518,-34.5965919494629,
25.3623580932617,-13.1085271835327,
11.6189279556274,5.14395046234131,
-17.7946319580078,8.34997558593750,
-43.0861206054688,7.01702117919922,
-52.4932823181152,-4.12826681137085,
-51.6382141113281,-30.2075157165527,
-38.5430221557617,-49.7029418945313,
-3.58020305633545,-32.9660224914551,
42.0254478454590,12.9989395141602,
60.9620857238770,49.3141555786133,
30.1304035186768,57.2065505981445,
-22.0529270172119,49.3396949768066,
-46.0731201171875,47.1680870056152,
-31.9012813568115,53.4753265380859,
-19.8764095306397,54.6167221069336,
-38.4428825378418,41.5682907104492,
-68.2111129760742,13.3227157592773,
-73.2980880737305,-27.2390213012695,
-50.2033195495606,-67.1807327270508,
-29.9602108001709,-80.8765945434570,
-27.1409187316895,-57.1083793640137,
-27.3778152465820,-22.2391395568848,
-14.4458265304565,-7.56906414031982,
2.60590028762817,-11.9157295227051,
3.45157313346863,-6.62212610244751,
-15.8955774307251,18.1269245147705,
-35.4288482666016,35.1459960937500,
-38.3018302917481,18.4056415557861,
-39.3739471435547,-22.6882553100586,
-53.0084114074707,-48.7249221801758,
-67.0470581054688,-45.6382217407227,
-50.0225753784180,-28.0051860809326,
3.96746134757996,-16.3177661895752,
51.2424774169922,-8.83823585510254,
44.3990783691406,-3.82051348686218,
-8.00022792816162,-10.1794471740723,
-42.5196990966797,-32.6790199279785,
-23.9942836761475,-53.3848915100098,
15.2255363464355,-42.2623329162598,
21.6793212890625,-3.84940934181213,
-4.03336000442505,31.4879627227783,
-14.7901506423950,36.9786796569824,
10.8642625808716,25.4440422058105,
43.5500068664551,22.4587192535400,
46.8585700988770,33.1901893615723,
31.2107143402100,39.9097328186035,
24.5319786071777,31.1565628051758,
31.9495792388916,16.0687408447266,
28.8111267089844,2.77126979827881,
13.2380352020264,-6.50353574752808,
2.00773715972900,-12.3754911422730,
4.09172534942627,-8.26430702209473,
5.25127792358398,7.60180282592773,
-8.47888946533203,22.5153236389160,
-20.8114032745361,25.5363979339600,
-16.9487991333008,23.8839397430420,
-10.7843103408813,32.3761520385742,
-20.8684158325195,51.4216690063477,
-43.0792198181152,56.5694656372070,
-52.1868515014648,33.8117256164551,
-39.2183113098145,-4.52304601669312,
-25.8281173706055,-32.1602783203125,
-34.7289543151856,-38.6684608459473,
-54.6124534606934,-28.3657760620117,
-59.3512611389160,-12.6027803421021,
-37.7398223876953,4.16687679290772,
-8.16235065460205,21.6258163452148,
5.45134449005127,32.3150444030762,
-6.24327421188355,24.4958019256592,
-31.7718238830566,-1.56750607490540,
-47.4722099304199,-27.0659122467041,
-35.7036590576172,-29.5520477294922,
0.713046550750732,-3.79370999336243,
39.2208518981934,24.8403015136719,
50.0820770263672,22.1056480407715,
28.5146522521973,-7.33264732360840,
-0.725850939750671,-20.9247055053711,
-10.4190845489502,6.90744304656982,
2.78933000564575,40.7276000976563,
18.3789882659912,27.8727035522461,
17.1814098358154,-27.9991989135742,
5.73293685913086,-60.9699974060059,
-4.62678956985474,-31.1420307159424,
-11.9612102508545,22.4655685424805,
-25.4907493591309,34.1804771423340,
-38.9010658264160,4.10224771499634,
-35.4104309082031,-12.2396812438965,
-17.2059478759766,8.01059532165527,
-14.4622268676758,28.2034683227539,
-41.7473831176758,12.8364686965942,
-72.6941986083984,-16.5329399108887,
-60.2683334350586,-15.9733743667603,
-2.38073062896729,7.84626054763794,
46.5225830078125,15.1881980895996,
42.0914154052734,-5.17490911483765,
0.0178995132446289,-20.0657539367676,
-30.9839649200439,-6.01012516021729,
-29.6979312896729,15.6772699356079,
-14.5087518692017,6.72151184082031,
-4.00216484069824,-32.5692062377930,
-0.868140816688538,-56.3827781677246,
-3.56395506858826,-38.0602111816406,
-16.3313179016113,0.647792816162109,
-31.3512058258057,18.4454345703125,
-22.4712333679199,-1.64145147800446,
14.0478410720825,-31.5148468017578,
43.5651855468750,-26.0672092437744,
32.0813713073731,19.9111557006836,
-3.45391130447388,62.9460334777832,
-14.0880041122437,62.7242469787598,
12.5589752197266,30.7896823883057,
33.4308700561523,10.8011503219605,
18.4731502532959,19.6034336090088,
-6.48240756988525,22.7895298004150,
-3.40342259407043,-10.4831180572510,
26.3212833404541,-51.9464263916016,
42.4842987060547,-46.7466430664063,
23.4571094512939,4.06915616989136,
-6.64709663391113,34.2591247558594,
-17.5239353179932,7.68549728393555,
-6.46535539627075,-35.0660858154297,
9.90927219390869,-30.9036960601807,
15.3244590759277,17.1490859985352,
3.31332015991211,46.7031288146973,
-23.7361621856689,25.8768501281738,
-46.6052398681641,-3.92712879180908,
-40.2733879089356,1.22286486625671,
-9.70235347747803,27.3774719238281,
8.49352836608887,34.4740142822266,
-6.60952568054199,16.8788013458252,
-30.4057197570801,7.14389276504517,
-21.3605308532715,12.4803743362427,
19.5907859802246,4.07065820693970,
50.0823097229004,-29.0252723693848,
40.0428962707520,-50.9574394226074,
9.86698722839356,-33.4923973083496,
-8.14079666137695,6.38433361053467,
-11.9630737304688,29.4485816955566,
-17.2898101806641,25.3097419738770,
-26.2093391418457,20.4018707275391,
-25.0822315216064,30.5183601379395,
-11.1069335937500,39.7423019409180,
4.93765735626221,33.0964202880859,
13.0507316589355,17.9897212982178,
17.6369152069092,3.44288635253906,
20.9862461090088,-10.5645418167114,
22.2925968170166,-21.5213489532471,
23.5658683776855,-16.5189800262451,
28.6427688598633,-1.42387962341309,
32.3778839111328,-1.31867265701294,
21.7620048522949,-24.8522377014160,
-5.01964855194092,-42.7406044006348,
-25.1423168182373,-20.2458477020264,
-21.1363105773926,31.1540775299072,
-7.36196279525757,54.5308456420898,
-14.4434251785278,25.2626190185547,
-47.3892478942871,-19.9391422271729,
-76.6520767211914,-36.5137023925781,
-70.0798797607422,-20.3836212158203,
-28.2209529876709,-2.54403877258301,
12.1773433685303,0.280612915754318,
19.4779090881348,-9.86233806610107,
-4.29435396194458,-24.0555915832520,
-27.1404685974121,-37.4780349731445,
-21.7665557861328,-35.1060829162598,
9.14412307739258,-4.33282470703125,
31.2428665161133,35.1147537231445,
17.1237602233887,43.0403594970703,
-19.4864215850830,1.79385876655579,
-33.3070678710938,-48.4553871154785,
-5.40174579620361,-53.8664093017578,
33.1779708862305,-11.8472862243652,
42.9509963989258,32.1820297241211,
24.5913639068604,41.7937431335449,
16.2800102233887,19.8611373901367,
35.5837097167969,-9.55204296112061,
53.5278053283691,-27.0476989746094,
36.3792381286621,-31.2164173126221,
8.62151527404785,-28.2334880828857,
13.1474819183350,-23.5528488159180,
48.2968482971191,-17.4358501434326,
62.2629508972168,-4.70427322387695,
29.4654312133789,24.5309658050537,
-7.27938127517700,57.2647972106934,
0.332311511039734,63.3530502319336,
31.8332176208496,34.0971260070801,
32.2493057250977,1.33551347255707,
-6.20516061782837,-9.54766368865967,
-28.3646793365479,-10.7007379531860,
-2.12426400184631,-25.8771438598633,
34.0702590942383,-44.3795394897461,
28.0030193328857,-34.9824981689453,
-6.62138223648071,-3.48983502388001,
-14.6432094573975,1.76812076568604,
25.0822391510010,-33.8723945617676,
68.4776382446289,-54.2353401184082,
72.4255752563477,-9.64569091796875,
35.1245498657227,61.9940071105957,
-11.1444482803345,71.5853347778320,
-36.9606895446777,7.49271392822266,
-29.5556526184082,-48.0156593322754,
4.70737266540527,-27.2014789581299,
49.4706764221191,40.1660537719727,
72.3535461425781,75.8730010986328,
53.7683029174805,55.9307060241699,
10.9872369766235,19.1979713439941,
-16.7998142242432,-0.0870138406753540,
-9.18402290344238,-10.7059717178345,
23.5990810394287,-17.6222972869873,
51.7989196777344,-7.70913314819336,
46.4498023986816,25.0051002502441,
7.22590446472168,52.0269279479981,
-30.9977684020996,48.3649559020996,
-33.1132431030273,30.4102573394775,
0.591607093811035,31.4621925354004,
30.4604148864746,42.9975395202637,
12.6599607467651,31.6051445007324,
-36.8518257141113,-9.86185359954834,
-62.9681282043457,-47.8617591857910,
-41.5740432739258,-49.2734336853027,
-11.6654014587402,-26.8346729278564,
-17.4528198242188,-22.7928066253662,
-38.0794754028320,-48.9316596984863,
-27.9632263183594,-73.4362792968750,
11.7438077926636,-59.9614944458008,
27.6178760528564,-17.0849494934082,
-7.12275028228760,10.6154098510742,
-43.7875900268555,-3.68139481544495,
-22.8743858337402,-39.8072738647461,
30.7274055480957,-47.4988212585449,
45.6218070983887,-6.71879005432129,
3.76170730590820,41.7406768798828,
-41.3835830688477,53.7302589416504,
-44.1052970886231,30.0980606079102,
-28.4323616027832,9.62118434906006,
-32.7586288452148,10.0148811340332,
-38.5418777465820,9.80462932586670,
-8.83449172973633,-11.6837234497070,
37.8763923645020,-30.3101844787598,
42.3495788574219,-12.8325281143188,
-4.36688852310181,22.2107257843018,
-39.9999923706055,18.3072719573975,
-13.7713003158569,-32.6335372924805,
41.1727638244629,-69.1772689819336,
55.6439056396484,-41.0078506469727,
19.2863445281982,17.2873954772949,
-11.6660585403442,28.6528244018555,
1.47783648967743,-21.0221405029297,
33.8025245666504,-58.4804801940918,
43.8369560241699,-28.2715759277344,
19.6332836151123,29.0934524536133,
-11.7251987457275,37.6111335754395,
-27.4430599212647,-9.07506179809570,
-31.9981784820557,-46.0046958923340,
-37.1952095031738,-33.1949005126953,
-39.0260238647461,-2.36745524406433,
-23.1091461181641,5.07086801528931,
4.07417917251587,5.13966560363770,
18.1742973327637,27.9732303619385,
3.57729005813599,54.8989868164063,
-24.1701965332031,42.3559188842773,
-25.3939285278320,-6.04299020767212,
10.5279283523560,-35.1566429138184,
41.8721351623535,-14.8831977844238,
26.3874816894531,14.1550369262695,
-24.1831417083740,7.09570264816284,
-57.0350914001465,-17.1633872985840,
-48.7358512878418,-12.1712455749512,
-26.5558071136475,23.3364353179932,
-24.8379974365234,46.4052124023438,
-32.9438133239746,34.0211486816406,
-16.4717445373535,2.40184450149536,
19.7185459136963,-22.9352149963379,
30.8137035369873,-32.4589271545410,
-0.461276531219482,-23.7815856933594,
-37.9275932312012,5.15462732315064,
-41.5429992675781,38.2799911499023,
-19.8218898773193,41.7550239562988,
-8.48380661010742,8.07147884368897,
-11.4693136215210,-22.0451774597168,
-0.528676867485046,-13.2973279953003,
29.2361106872559,11.4837789535522,
40.7114486694336,8.59115600585938,
15.3185596466064,-27.8403549194336,
-13.6040811538696,-60.7894668579102,
-3.43142533302307,-61.0864524841309,
35.1395835876465,-35.5496597290039,
41.7041969299316,-9.94911479949951,
-4.62507200241089,3.83874869346619,
-56.0991516113281,3.41563534736633,
-62.0638046264648,-13.8134317398071,
-28.1315441131592,-37.7476806640625,
3.19863986968994,-44.9260559082031,
10.9101514816284,-26.3240013122559,
7.97016668319702,-8.67456150054932,
12.9019498825073,-19.2240638732910,
21.2615051269531,-40.3017234802246,
27.6225299835205,-37.1269912719727,
36.9997787475586,-8.40791702270508,
47.3921508789063,19.4974288940430,
47.9735679626465,29.4785614013672,
40.8789329528809,32.4534683227539,
42.6117744445801,40.8172035217285,
46.1593437194824,46.1892242431641,
21.3580265045166,36.2097358703613,
-33.9789237976074,25.6231212615967,
-70.2314376831055,25.2669506072998,
-47.1499137878418,17.0727310180664,
2.95984172821045,-10.8937911987305,
13.8295936584473,-31.6352462768555,
-26.3611869812012,-11.2871398925781,
-50.1990814208984,27.1472187042236,
-17.4246997833252,23.7006549835205,
27.5059013366699,-30.2367229461670,
25.7411174774170,-67.6932678222656,
-9.53379917144775,-39.1602706909180,
-22.1672439575195,19.8860492706299,
-0.687050580978394,34.2070198059082,
11.0079460144043,-4.93949937820435,
-6.64522552490234,-31.9656391143799,
-21.3177928924561,-13.4330987930298,
-6.94251823425293,9.78054428100586,
14.3487167358398,-5.43550634384155,
13.8380479812622,-39.4964179992676,
6.87081003189087,-48.4329071044922,
26.7287864685059,-24.5721092224121,
59.6052589416504,3.10369253158569,
58.2341728210449,16.8948173522949,
14.5825500488281,19.0355968475342,
-27.6339282989502,7.13689708709717,
-32.7703819274902,-21.4460659027100,
-13.1859788894653,-41.7582550048828,
-2.51449441909790,-19.9789409637451,
-12.5126447677612,31.1910858154297,
-29.7999973297119,51.0915565490723,
-34.6716003417969,17.6318988800049,
-16.1282310485840,-16.8247051239014,
21.3726863861084,0.920361757278442,
57.1084785461426,44.6808700561523,
58.0747451782227,49.4660148620606,
11.8395023345947,6.93417930603027,
-46.9147605895996,-22.8202228546143,
-68.5613250732422,-1.24948227405548,
-43.5342254638672,35.6335487365723,
-3.21678018569946,30.4133739471436,
23.0166511535645,-8.30047130584717,
24.6808719635010,-28.4339199066162,
6.30706119537354,-7.46269273757935,
-20.1472625732422,18.8848590850830,
-38.1864891052246,14.8944797515869,
-22.9734458923340,-14.2115421295166,
21.9447898864746,-39.0047645568848,
58.7104835510254,-39.9981613159180,
54.5601005554199,-14.9761714935303,
25.4319152832031,17.7000122070313,
10.5358428955078,36.9931564331055,
20.9519824981689,30.6679592132568,
24.0836486816406,9.37928771972656,
-3.03743839263916,-2.26431083679199,
-31.3234844207764,8.48157691955566,
-22.5910701751709,25.6672115325928,
15.2321596145630,27.9338035583496,
36.0649452209473,25.1702213287354,
5.33242511749268,35.3831977844238,
-49.8223381042481,49.0978965759277,
-77.3900985717773,41.4715042114258,
-54.1632957458496,16.8283405303955,
-8.79595851898193,9.62347316741943,
12.4061412811279,35.9526138305664,
-6.15038108825684,60.4581375122070,
-39.1194000244141,36.1544837951660,
-46.9722023010254,-29.4532604217529,
-16.8306560516357,-80.0205612182617,
20.1789817810059,-78.8240966796875,
25.2575569152832,-37.9333686828613,
-2.97576689720154,4.52007007598877,
-25.5899276733398,32.8463745117188,
-12.1619901657105,48.1037445068359,
24.3030300140381,49.1975021362305,
46.2165489196777,36.0655174255371,
40.1173477172852,22.0279712677002,
28.0297355651855,21.0889244079590,
30.5569438934326,23.9239368438721,
31.2287158966064,14.1749572753906,
12.4169435501099,-5.21894931793213,
-21.6712093353272,-7.32847166061401,
-44.5517387390137,20.1570167541504,
-44.6913032531738,52.1538124084473,
-35.8633651733398,46.4408645629883,
-31.4065036773682,1.69229006767273,
-25.1123981475830,-43.0533905029297,
-9.86026477813721,-52.2388839721680,
4.43360805511475,-26.5324249267578,
4.05951499938965,-1.60446751117706,
-9.42271709442139,1.16736757755280,
-18.9877319335938,-5.10172176361084,
-22.8418254852295,0.943202853202820,
-32.3421478271484,21.3650703430176,
-49.5370254516602,28.3652667999268,
-57.5250701904297,9.38128757476807,
-42.8687438964844,-14.6467752456665,
-19.3346633911133,-13.0381660461426,
-4.52038955688477,16.0809097290039,
1.39295864105225,40.2166023254395,
10.8685884475708,34.6450233459473,
27.0001316070557,13.7026634216309,
31.7599964141846,13.7176628112793,
22.0651092529297,39.5985908508301,
9.73092555999756,61.2792015075684,
3.78646469116211,56.1224174499512,
-10.2876319885254,26.2658157348633,
-39.2200698852539,-5.57158517837524,
-61.6913108825684,-29.2156066894531,
-51.2108001708984,-46.9202003479004,
-10.0803060531616,-51.7656631469727,
31.2268562316895,-33.6793594360352,
47.8602752685547,-0.861307740211487,
41.1941413879395,17.1773319244385,
23.9251441955566,10.5586118698120,
-1.64644777774811,2.61085700988770,
-30.4353771209717,15.6703758239746,
-49.9796638488770,28.6843185424805,
-51.0806694030762,4.63219738006592,
-39.0693969726563,-48.9239501953125,
-21.4907684326172,-75.9634552001953,
5.83893871307373,-41.9228630065918,
35.5674400329590,11.8576011657715,
42.9640998840332,26.7628574371338,
16.2970466613770,-3.68497967720032,
-21.4553146362305,-29.8682594299316,
-28.4510402679443,-25.6471176147461,
-1.82154107093811,-19.6830196380615,
23.6493949890137,-34.8795776367188,
18.9542808532715,-53.4409523010254,
-1.92519819736481,-41.1532325744629,
-14.4009704589844,-12.5428438186646,
-18.4918251037598,-9.22094917297363,
-23.9341220855713,-39.4120903015137,
-19.2888183593750,-58.6184043884277,
8.12945365905762,-29.8787441253662,
31.7724895477295,29.3324279785156,
16.9716854095459,64.8465881347656,
-31.0032958984375,46.8607177734375,
-57.0421485900879,-0.229543924331665,
-25.9180278778076,-37.2219734191895,
28.5191650390625,-39.5153884887695,
51.0640296936035,-7.80673456192017,
32.2430343627930,34.0014419555664,
9.06791591644287,61.2308197021484,
4.68977117538452,64.6267318725586,
6.08504915237427,48.6026649475098,
1.64286983013153,24.9970436096191,
5.19822883605957,7.94588994979858,
17.0617389678955,6.64195537567139,
14.3775310516357,20.0244789123535,
-17.3007678985596,32.8176155090332,
-50.9156303405762,24.1219406127930,
-45.6433486938477,-12.6007499694824,
-3.87241888046265,-42.3560600280762,
33.5508956909180,-28.7744884490967,
36.3543777465820,10.3210048675537,
18.0561542510986,24.6438789367676,
7.05282783508301,-5.49115705490112,
7.76456308364868,-38.0826568603516,
7.93073987960815,-26.4418449401855,
2.28700852394104,10.0577840805054,
-11.0153188705444,10.2841243743896,
-30.6117839813232,-31.4244403839111,
-49.9513626098633,-53.6182594299316,
-50.9988479614258,-15.6212444305420,
-25.7364120483398,32.6029434204102,
12.8981046676636,19.1687831878662,
38.8255653381348,-40.8800582885742,
39.7636528015137,-63.9577598571777,
26.0393123626709,-15.5700473785400,
18.0169105529785,38.2960662841797,
20.0925903320313,32.2731590270996,
25.7340526580811,-9.41837692260742,
22.1542987823486,-15.9514980316162,
1.56933760643005,23.9441986083984,
-25.0299644470215,48.0379142761231,
-36.5701675415039,16.6133861541748,
-22.6509838104248,-31.7578582763672,
-2.74860119819641,-41.8590011596680,
-5.86057853698731,-10.8513879776001,
-30.9771556854248,21.8202705383301,
-49.7549476623535,33.5623474121094,
-41.0198860168457,29.8986988067627,
-17.3820838928223,17.2721347808838,
-4.62400484085083,8.01051712036133,
-10.6220407485962,16.7795143127441,
-22.4054317474365,41.7439727783203,
-30.8864421844482,57.1172447204590,
-31.4473896026611,32.3603973388672,
-19.9107742309570,-16.8332443237305,
7.80453014373779,-31.8057575225830,
37.0692367553711,4.70088052749634,
43.2745018005371,41.5698471069336,
25.0041122436523,28.4953041076660,
9.36403083801270,-19.3418083190918,
16.5866394042969,-54.1105155944824,
34.0687026977539,-53.0292472839356,
32.2760658264160,-26.6930046081543,
7.27545261383057,7.57357406616211,
-16.3600730895996,35.6127548217773,
-21.0337486267090,35.3628120422363,
-12.6761713027954,-7.48010063171387,
-2.34736299514771,-55.9664878845215,
12.2894096374512,-45.9739761352539,
28.5654659271240,19.0350532531738,
25.5247955322266,64.5865020751953,
-6.89622259140015,39.8878440856934,
-41.3166961669922,-7.18923425674439,
-35.3746643066406,-9.78101253509522,
7.45572614669800,18.4138069152832,
34.3378829956055,14.7697257995605,
9.81463623046875,-22.3110923767090,
-40.4006271362305,-32.7600746154785,
-57.9553718566895,5.43330860137939,
-31.6496639251709,30.3233318328857,
1.44005370140076,-9.83443546295166,
10.8801622390747,-64.6319961547852,
8.38112640380859,-51.5368194580078,
12.7997503280640,21.6532554626465,
19.1053676605225,70.9815521240234,
15.0919113159180,54.0759201049805,
4.57051944732666,15.6592388153076,
-0.272208333015442,7.19779396057129,
-2.29449582099915,21.9648113250732,
-12.8348894119263,30.6163520812988,
-21.2220573425293,28.5694751739502,
-10.6574802398682,28.0167026519775,
9.35739612579346,26.7356033325195,
3.56368136405945,12.5054750442505,
-31.2389965057373,-4.70747756958008,
-53.6451606750488,-4.55518102645874,
-35.6814193725586,4.37647008895874,
-4.26144075393677,-5.11078929901123,
2.52066850662231,-29.4982852935791,
-9.48361110687256,-33.0348434448242,
-2.83644962310791,-2.78190302848816,
24.0641422271729,28.0060997009277,
25.3654174804688,31.8908386230469,
-18.6447830200195,16.1440639495850,
-62.8306961059570,3.18286943435669,
-58.4258880615234,-8.00249195098877,
-22.4326000213623,-28.4272651672363,
-10.4575834274292,-47.2977485656738,
-35.1258430480957,-38.9766921997070,
-48.5456466674805,-7.76640796661377,
-18.5386657714844,9.56934547424316,
25.5438747406006,-11.8244724273682,
39.3247108459473,-48.0563430786133,
21.1259841918945,-58.3442802429199,
4.49337959289551,-31.4239311218262,
5.48008489608765,4.17660760879517,
2.35307836532593,18.2379570007324,
-17.1849613189697,4.53441619873047,
-34.0886993408203,-17.7434711456299,
-26.0939884185791,-24.4170074462891,
0.572412490844727,-11.9795494079590,
15.0486049652100,4.40365314483643,
1.70236575603485,6.49320745468140,
-23.5008850097656,-4.33331966400147,
-28.8387584686279,-11.5300064086914,
-4.41817760467529,-5.58382081985474,
27.7033042907715,7.31280708312988,
32.1919937133789,5.97284269332886,
-2.79545164108276,-12.9406518936157,
-51.2218170166016,-34.7032318115234,
-70.4096069335938,-49.6928062438965,
-39.0938987731934,-55.9295692443848,
16.2795944213867,-51.5754699707031,
43.6027717590332,-35.2556114196777,
20.6249198913574,-10.1874380111694,
-27.4139785766602,8.92145633697510,
-55.6165428161621,12.1048450469971,
-40.4292297363281,10.8523015975952,
1.96676838397980,21.2064609527588,
29.8661289215088,30.9156188964844,
22.0365314483643,7.75531291961670,
-1.05109786987305,-44.9531059265137,
-3.85012531280518,-70.5662841796875,
23.8466415405273,-30.6577835083008,
45.8859481811523,32.8628692626953,
21.4841747283936,44.7489662170410,
-35.7938575744629,-6.27628755569458,
-57.7443656921387,-52.6697463989258,
-5.80189132690430,-41.1537437438965,
70.9585418701172,-0.460423231124878,
82.2029037475586,9.65746688842773,
17.1850643157959,-4.25113773345947,
-38.5162849426270,0.296088576316834,
-18.2393798828125,22.6194438934326,
41.9063301086426,18.5553340911865,
53.6252746582031,-11.5301189422607,
1.80525445938110,-16.8331489562988,
-41.2932281494141,20.6120853424072,
-30.1464080810547,41.5499572753906,
-2.93845486640930,3.34151625633240,
-13.5521039962769,-44.6552276611328,
-45.5469360351563,-31.1663379669189,
-51.9686050415039,28.1647148132324,
-30.1360168457031,49.0947341918945,
-22.4094276428223,5.65407562255859,
-37.7452507019043,-31.6524257659912,
-38.0387649536133,-12.0115165710449,
-9.67703533172607,23.2431240081787,
9.19138240814209,20.0095367431641,
-12.0123815536499,-3.37717247009277,
-48.5574493408203,6.19011068344116,
-53.2360458374023,45.9337387084961,
-23.4656600952148,63.9813003540039,
1.34906268119812,42.2117004394531,
9.44123554229736,18.3207378387451,
20.3912010192871,19.8402576446533,
40.7086143493652,26.8660392761230,
52.2512702941895,11.5448942184448,
42.1663513183594,-6.74298429489136,
23.5132350921631,3.91711950302124,
9.16674137115479,33.7565650939941,
-2.30459737777710,45.0161666870117,
-17.0678215026855,28.0145759582520,
-20.7230854034424,6.90005397796631,
-3.21784830093384,0.427055805921555,
18.9859046936035,5.64428234100342,
21.0495338439941,9.48525142669678,
10.0395765304565,7.65856695175171,
15.5960159301758,7.25179147720337,
38.2380371093750,13.4775438308716,
45.2932014465332,22.9947910308838,
21.1955261230469,33.0980796813965,
-8.22318553924561,39.3002471923828,
-11.4935741424561,37.2101058959961,
1.72066104412079,30.1245841979980,
-0.307138293981552,27.0077247619629,
-21.7534980773926,22.5892543792725,
-32.8399162292481,1.27826619148254,
-20.4616661071777,-34.8088798522949,
-7.41707944869995,-62.5727310180664,
-20.8069820404053,-64.1334838867188,
-48.4837608337402,-48.1976890563965,
-56.5933341979981,-40.4335136413574,
-38.2908706665039,-39.5469512939453,
-22.1256351470947,-23.2869606018066,
-27.0578136444092,17.1062526702881,
-36.9981994628906,55.9442138671875,
-26.0290374755859,60.2140998840332,
1.85810291767120,33.6182746887207,
14.3841896057129,10.5738792419434,
-7.78446292877197,12.1940536499023,
-37.8012504577637,18.1256828308105,
-36.6525764465332,-0.464617013931274,
0.524438381195068,-40.0201530456543,
37.0215110778809,-60.5926628112793,
41.7916069030762,-33.2741317749023,
18.7382907867432,22.0193424224854,
-3.94243955612183,51.7798309326172,
-14.9605302810669,26.5663757324219,
-24.1902198791504,-23.4713478088379,
-35.3542137145996,-46.4762878417969,
-29.1859207153320,-21.9168090820313,
0.877126574516296,19.0554904937744,
31.1445808410645,36.4588928222656,
29.7793502807617,21.8337154388428,
-2.76177930831909,3.91164183616638,
-31.7141265869141,4.00821971893311,
-32.9482460021973,10.1177577972412,
-18.3526325225830,4.35487556457520,
-16.3991832733154,-11.8156948089600,
-27.5996036529541,-17.7514305114746,
-29.7279834747314,0.409777134656906,
-11.9911670684814,27.7596073150635,
7.96855497360230,38.8002738952637,
4.86504602432251,31.7654323577881,
-19.9868659973145,20.1507530212402,
-41.8402900695801,7.46121549606323,
-43.9570541381836,-10.4387245178223,
-31.9629001617432,-25.5954170227051,
-23.3659458160400,-12.6260490417480,
-24.0744190216064,32.0909080505371,
-31.6728591918945,65.4671859741211,
-41.7758102416992,40.3530158996582,
-51.7179489135742,-26.6347236633301,
-52.0020446777344,-65.6768951416016,
-34.8975105285645,-32.5930786132813,
-6.79025268554688,31.6997985839844,
12.5693273544312,55.8630905151367,
9.20018196105957,26.5724296569824,
-8.82538414001465,-11.0014963150024,
-25.5059814453125,-19.8006019592285,
-25.7471160888672,-7.21567964553833,
-8.19264793395996,2.39796209335327,
20.1397819519043,-3.59830379486084,
42.9980964660645,-21.7902889251709,
45.1360054016113,-44.7478370666504,
22.5709571838379,-57.3915176391602,
3.51556015014648,-38.9113502502441,
12.7398242950439,-2.35643863677979,
42.0777854919434,10.3481245040894,
56.6288566589356,-19.9431648254395,
42.0082054138184,-52.1331291198731,
17.8517456054688,-31.3855686187744,
5.93538093566895,25.6813354492188,
-3.11511540412903,49.7713890075684,
-27.9381217956543,14.3765792846680,
-54.5317382812500,-28.8350296020508,
-52.4227066040039,-22.1990985870361,
-26.1286087036133,15.9638681411743,
-19.8852615356445,21.5876235961914,
-50.1981849670410,-24.0271072387695,
-73.8881225585938,-70.3771743774414,
-48.1209564208984,-64.3571090698242,
8.48327159881592,-15.2757930755615,
34.5086669921875,29.8594551086426,
13.6286315917969,41.2500267028809,
-12.1789455413818,28.2243423461914,
-2.71947789192200,13.9654541015625,
22.4847431182861,9.92184925079346,
25.9639186859131,10.6369190216064,
3.00522756576538,6.07126045227051,
-15.5883617401123,-6.35552406311035,
-20.5145759582520,-9.62901973724365,
-21.8135814666748,4.54939222335815,
-18.9732532501221,23.5599822998047,
0.993822097778320,21.2767181396484,
32.3583717346191,-7.43809795379639,
49.5312805175781,-35.4643096923828,
44.2184638977051,-33.3918762207031,
38.8361511230469,-7.73226165771484,
43.8851852416992,6.33435249328613,
37.9392929077148,-6.98941278457642,
-1.63970243930817,-29.9181003570557,
-48.3903846740723,-36.6863822937012,
-56.4436683654785,-20.1466102600098,
-34.3444747924805,3.66122627258301,
-28.5852699279785,20.4751033782959,
-51.4234428405762,24.8780364990234,
-58.6237449645996,22.4073390960693,
-17.1150093078613,21.2856101989746,
41.3025016784668,27.2922039031982,
61.8747863769531,32.8080825805664,
40.9604606628418,23.0257873535156,
19.9965229034424,1.09881150722504,
18.8838958740234,-10.8226737976074,
22.3814449310303,8.35495948791504,
18.1292266845703,46.4989166259766,
23.1503009796143,63.6926116943359,
40.7754821777344,39.8434028625488,
40.7680320739746,-1.85115957260132,
-1.83753967285156,-25.7904396057129,
-55.7194938659668,-21.1448364257813,
-64.5638427734375,-6.99096488952637,
-20.7812232971191,-6.44263076782227,
27.2613925933838,-19.7929286956787,
34.3286743164063,-29.2386493682861,
8.92249584197998,-22.8613071441650,
-4.04479312896729,0.590409159660339,
17.1681041717529,30.7846813201904,
43.4589157104492,46.5357818603516,
43.8611984252930,33.4734153747559,
16.7162551879883,4.88733100891113,
-7.77927684783936,-5.86752033233643,
-11.6432552337646,14.0468225479126,
-7.29307317733765,37.3660469055176,
-15.1001482009888,23.6196193695068,
-28.7716159820557,-20.1392688751221,
-26.2226371765137,-44.8220977783203,
-1.05720341205597,-22.2167606353760,
13.8321971893311,9.14379501342773,
-7.61345911026001,-1.88467383384705,
-47.5708084106445,-41.0351943969727,
-62.8041000366211,-46.4908256530762,
-34.6220741271973,-3.09029722213745,
12.9954566955566,29.5067043304443,
44.7334938049316,2.34246540069580,
48.3223609924316,-44.7092781066895,
33.3665504455566,-34.9539642333984,
10.1533813476563,28.0895767211914,
-8.36423778533936,65.8882522583008,
-11.3755655288696,35.8046951293945,
4.66890144348145,-10.0022106170654,
19.0991821289063,-3.57119727134705,
8.07132053375244,41.7128829956055,
-23.2950801849365,54.9517211914063,
-47.8637504577637,14.7090053558350,
-50.4313163757324,-27.3612117767334,
-42.4178886413574,-29.1532993316650,
-37.8902664184570,-8.01379299163818,
-28.5011329650879,-4.18757104873657,
-4.98093223571777,-19.2437477111816,
17.5050601959229,-21.9938507080078,
17.6112594604492,-0.126964807510376,
-0.332336425781250,21.1805610656738,
0.239110589027405,17.7561359405518,
31.3752079010010,-2.82806563377380,
63.2121047973633,-16.8775959014893,
55.7731704711914,-13.7717590332031,
13.3044862747192,1.37064540386200,
-15.7355365753174,10.8573760986328,
-2.07704234123230,4.16584444046021,
29.5587406158447,-9.58634471893311,
36.6452140808106,-13.4436922073364,
8.10230541229248,-3.44966983795166,
-23.4998512268066,9.46280574798584,
-30.2438030242920,9.51392364501953,
-20.2202053070068,-4.83145570755005,
-12.2519826889038,-16.2206993103027,
-6.51836013793945,-14.5489673614502,
9.40831375122070,-5.09104537963867,
34.7304000854492,5.25747203826904,
46.3982849121094,16.7173500061035,
25.6429347991943,29.0970973968506,
-13.3898639678955,31.2613925933838,
-39.6590156555176,9.31353759765625,
-31.7417945861816,-27.7484817504883,
6.14951896667481,-45.6653404235840,
47.8644180297852,-20.2727699279785,
58.0382614135742,31.2978153228760,
19.0336818695068,66.4717407226563,
-38.7325096130371,58.9198913574219,
-59.5659751892090,26.6166191101074,
-29.8778591156006,10.5203714370728,
1.63702821731567,23.0373172760010,
-15.0259590148926,30.1895847320557,
-60.3892211914063,2.89880967140198,
-62.0602951049805,-38.5190925598145,
-1.59362125396729,-49.1879081726074,
52.0825614929199,-13.2113380432129,
34.8000411987305,25.0068340301514,
-24.5007915496826,20.8694915771484,
-53.0198936462402,-8.21066665649414,
-33.4904365539551,-11.5523605346680,
-13.0773925781250,17.8092041015625,
-21.0462112426758,34.9469490051270,
-30.9205398559570,15.5562171936035,
-17.6613273620605,-7.68922853469849,
-7.22119188308716,5.28727149963379,
-23.0593547821045,36.4134750366211,
-39.4871292114258,25.6560516357422,
-17.0890235900879,-27.9366741180420,
30.1054763793945,-51.7523612976074,
43.6637344360352,3.00442242622376,
9.25452232360840,84.0356063842773,
-24.0517635345459,94.4726333618164,
-14.5612182617188,20.0997085571289,
17.0519065856934,-54.2000999450684,
33.8862876892090,-50.1347885131836,
27.2021141052246,2.84964299201965,
14.8829584121704,23.6840324401855,
10.4786291122437,-5.78307771682739,
10.8098402023315,-23.2808895111084,
15.7435455322266,7.54619073867798,
24.1365661621094,41.5737228393555,
24.1418399810791,23.8426475524902,
6.19863557815552,-24.4548435211182,
-12.8114604949951,-35.1118011474609,
-6.39098978042603,5.53164243698120,
16.8434181213379,42.7700920104981,
20.2566890716553,40.4385375976563,
-1.53772854804993,27.3913745880127,
-15.9985446929932,37.5428733825684,
-1.87189567089081,52.9128456115723,
18.2379856109619,39.9825553894043,
14.1727905273438,14.0485115051270,
-5.80802726745606,17.4011306762695,
-12.4935321807861,43.2919044494629,
-2.39812564849854,43.1606712341309,
3.95168876647949,1.37335836887360,
2.51087117195129,-40.1728591918945,
14.8651094436646,-44.3045501708984,
45.4300613403320,-30.4361667633057,
62.0415954589844,-31.3021392822266,
42.9509849548340,-41.5026016235352,
13.6517696380615,-36.1802902221680,
10.6252021789551,-19.3506622314453,
33.0462265014648,-17.5573444366455,
50.5636825561523,-26.9490909576416,
43.2943496704102,-7.11252880096436,
18.8018665313721,43.0472221374512,
-9.09687900543213,73.7799377441406,
-31.3574085235596,45.2161865234375,
-35.4536666870117,-12.3864507675171,
-13.6860704421997,-38.7709770202637,
13.5262422561646,-9.74828338623047,
8.36786556243897,38.9271125793457,
-29.4082050323486,53.4427757263184,
-54.0644454956055,21.5719223022461,
-32.0466117858887,-22.2635803222656,
4.48008441925049,-39.7236709594727,
2.24027681350708,-16.4877109527588,
-34.2221946716309,17.3830547332764,
-49.5270195007324,17.1626167297363,
-12.4479875564575,-30.9341068267822,
36.4213409423828,-76.4094619750977,
43.8619461059570,-66.6812896728516,
10.6464004516602,-17.7456302642822,
-16.3609924316406,4.97510290145874,
-11.7658538818359,-23.8717422485352,
3.00989174842834,-53.9879302978516,
-3.06311035156250,-32.0333290100098,
-24.4230918884277,20.9673614501953,
-37.8367500305176,32.5499534606934,
-39.0549392700195,-11.6620988845825,
-38.3504066467285,-49.9539756774902,
-37.4524803161621,-40.1131477355957,
-24.4285659790039,-11.3512134552002,
13.7897558212280,-0.523253321647644,
55.8229751586914,7.56113338470459,
60.4979782104492,40.5085563659668,
17.0909881591797,66.1732406616211,
-27.9626140594482,35.2202377319336,
-24.3696174621582,-30.8773021697998,
22.6502513885498,-51.0516586303711,
50.6599655151367,-4.54693412780762,
18.1696434020996,34.1718978881836,
-34.4710578918457,4.16767024993897,
-35.4978942871094,-48.7810440063477,
19.5261669158936,-47.3347396850586,
56.8692588806152,-4.44165706634522,
25.0042934417725,7.25893020629883,
-38.0359230041504,-25.1723880767822,
-59.5533599853516,-43.4965400695801,
-29.4527435302734,-21.4529094696045,
1.62891519069672,-6.43268632888794,
-2.65477490425110,-31.5731201171875,
-16.6504325866699,-55.3576889038086,
-3.31439614295959,-28.2984714508057,
24.0170269012451,15.5311155319214,
31.5938911437988,10.5572490692139,
17.8677444458008,-38.4355392456055,
8.63946342468262,-56.9784088134766,
12.1517410278320,-17.4444980621338,
6.90695858001709,19.1392650604248,
-15.1936368942261,-0.548951625823975,
-23.6794681549072,-41.0333404541016,
3.26527857780457,-44.2377700805664,
36.9836769104004,-1.83667159080505,
32.9265098571777,41.4488449096680,
-7.52586412429810,54.5516662597656,
-37.0898780822754,48.8442382812500,
-22.8415431976318,47.0243492126465,
7.86418008804321,42.8593101501465,
13.4855384826660,25.7420330047607,
-4.28626680374146,0.127480924129486,
-9.95445823669434,-17.9915390014648,
9.87365341186523,-21.8232498168945,
26.6718330383301,-10.5438861846924,
19.8007793426514,6.20703315734863,
0.0988909006118774,3.76594877243042,
-3.11065673828125,-31.3539142608643,
9.62059307098389,-73.5425109863281,
13.5558938980103,-76.0326080322266,
-2.46874427795410,-29.8610534667969,
-21.4215068817139,17.6605415344238,
-22.7523803710938,14.9167890548706,
-13.0416584014893,-28.5793743133545,
-6.06705999374390,-55.9444465637207,
-7.10106134414673,-41.4952888488770,
-4.12062501907349,-12.0698051452637,
13.5912876129150,-2.63567399978638,
40.0244522094727,-3.32335233688355,
51.5759963989258,10.9143314361572,
31.7167778015137,35.3637123107910,
-14.7679738998413,35.9980812072754,
-58.2182235717773,1.49861049652100,
-67.6894912719727,-39.1655006408691,
-38.8294219970703,-50.5805282592773,
-2.86711430549622,-33.6379241943359,
9.18447589874268,-14.0683765411377,
6.87534570693970,-7.85515594482422,
19.0411891937256,-9.63606929779053,
47.0696487426758,-3.83968830108643,
64.1728973388672,8.21722984313965,
52.7510375976563,13.4343767166138,
32.9942321777344,9.83347606658936,
35.5524368286133,2.85312795639038,
50.4894027709961,7.67247438430786,
43.9979248046875,26.0219993591309,
7.71452140808106,41.4833984375000,
-26.7490482330322,35.5954895019531,
-38.2738838195801,8.79404830932617,
-34.1475944519043,-21.3754062652588,
-23.8351745605469,-38.5806694030762,
0.214086920022964,-40.2568969726563,
38.7797622680664,-27.3744201660156,
54.3508605957031,-4.74450683593750,
20.2377376556397,21.4045333862305,
-33.4984512329102,28.5032653808594,
-43.1011314392090,-1.04962790012360,
5.57369899749756,-51.0036163330078,
58.6252059936523,-76.7048797607422,
63.5691528320313,-53.9194602966309,
39.4802398681641,-8.25713443756104,
28.1315155029297,15.9566612243652,
31.8968811035156,4.66527271270752,
18.5687122344971,-21.1782417297363,
-13.1195011138916,-36.3711509704590,
-30.2222232818604,-36.3502731323242,
-19.0797309875488,-22.2327251434326,
1.35399258136749,9.78427219390869,
9.34541988372803,51.1359100341797,
14.4912738800049,69.8139801025391,
27.0737342834473,45.4541969299316,
31.9472332000732,2.71726799011230,
13.8758668899536,-13.7518720626831,
-6.80199337005615,3.54695868492126,
0.663028597831726,14.4373083114624,
26.5074939727783,-7.56599092483521,
36.6259994506836,-30.0738162994385,
25.0647144317627,-16.4825801849365,
8.58858585357666,20.1337242126465,
-7.07585048675537,27.2662200927734,
-32.5106086730957,-10.0796251296997,
-58.7139244079590,-43.3362503051758,
-55.3592681884766,-25.5293197631836,
-17.6501979827881,19.4756603240967,
13.2839412689209,30.4287185668945,
3.60153007507324,-10.8143081665039,
-16.4259490966797,-58.8935661315918,
-0.0623939037322998,-60.6781234741211,
40.9301528930664,-16.9670906066895,
50.0143928527832,26.8440761566162,
16.8160076141357,29.0120525360107,
-9.01278972625732,-5.82955121994019,
1.45877742767334,-36.2507247924805,
15.2203540802002,-32.4438362121582,
-5.60610103607178,-3.20415067672730,
-38.8162422180176,12.9840106964111,
-38.5315055847168,-8.22912597656250,
-6.93360090255737,-36.1599769592285,
6.67390680313110,-22.4104328155518,
-11.6587686538696,33.2421188354492,
-25.8823394775391,71.1623001098633,
-5.93200254440308,53.9053077697754,
25.7615814208984,11.6016855239868,
36.8718376159668,-2.30304455757141,
35.9182472229004,17.2796974182129,
45.4756011962891,27.9101562500000,
54.6744461059570,7.84352636337280,
39.2837028503418,-2.08630824089050,
1.49519371986389,26.9191627502441,
-30.5923423767090,54.5850639343262,
-39.4750061035156,30.1238803863525,
-39.0187568664551,-28.0685729980469,
-48.4092941284180,-57.6933746337891,
-59.1927375793457,-46.0555343627930,
-53.6339836120606,-37.7864379882813,
-28.7790870666504,-54.7207984924316,
7.02154350280762,-56.2882461547852,
41.0845375061035,-12.6907482147217,
57.3190536499023,37.1042060852051,
42.9392547607422,43.0225601196289,
15.5990009307861,22.2726631164551,
11.8603734970093,33.0811882019043,
39.1238479614258,63.0220489501953,
61.3964805603027,49.3022460937500,
40.8679580688477,-11.4754657745361,
-2.86111307144165,-40.7611198425293,
-18.8221092224121,2.50187611579895,
12.0492277145386,49.0841217041016,
51.3231658935547,25.9319496154785,
56.4542961120606,-35.6067733764648,
32.0949707031250,-46.0915145874023,
8.89346885681152,0.500574111938477,
-9.59152603149414,23.3273239135742,
-26.3374958038330,-9.09674835205078,
-31.8494262695313,-33.2896690368652,
-16.0834999084473,4.55010128021240,
7.64951753616333,52.6583938598633,
12.2831954956055,31.1637401580811,
-2.28271317481995,-40.3439254760742,
-12.8989086151123,-73.5753860473633,
-9.65261268615723,-33.8541755676270,
-13.3031816482544,22.2032699584961,
-22.3376159667969,38.1674041748047,
-5.68280410766602,22.5772647857666,
47.8739204406738,24.1239681243897,
80.2704086303711,52.4831619262695,
33.6583061218262,71.1790924072266,
-51.7127990722656,50.6687316894531,
-77.1886672973633,8.49927711486816,
-15.2765560150146,-21.0928115844727,
48.1026535034180,-13.8183422088623,
29.5515670776367,21.1767826080322,
-36.4065666198731,45.9114875793457,
-48.4932746887207,32.6143493652344,
13.0552024841309,-1.93377661705017,
64.4603271484375,-14.1420774459839,
39.7376251220703,5.48771524429321,
-24.3678569793701,20.4661788940430,
-56.3547325134277,-0.720452129840851,
-45.9991035461426,-42.2101211547852,
-30.2481594085693,-56.7298126220703,
-24.0320301055908,-35.5261497497559,
-11.4927110671997,-19.7594108581543,
2.18667411804199,-39.1672096252441,
-3.52250576019287,-66.6196975708008,
-24.8405838012695,-58.3422012329102,
-24.0579986572266,-15.6805114746094,
19.0076503753662,20.8454151153564,
64.4799804687500,27.2180538177490,
66.2849960327148,17.1932888031006,
36.0640220642090,12.2347860336304,
11.3121528625488,13.8368949890137,
1.84979367256165,14.9682950973511,
-4.12543916702271,13.1744651794434,
-6.15893650054932,11.5740928649902,
0.150339603424072,9.31354999542236,
9.32575416564941,8.53579044342041,
8.73652362823486,17.5880298614502,
5.37246894836426,30.9557151794434,
21.2592468261719,22.6377296447754,
42.4030380249023,-18.0008964538574,
30.7881107330322,-56.6085815429688,
-16.3800849914551,-46.3921546936035,
-41.4447517395020,4.49898242950439,
-6.62232112884522,35.9687995910645,
44.7744979858398,14.3428859710693,
51.0583457946777,-23.3146648406982,
18.5454635620117,-21.0826187133789,
0.588660299777985,19.8497295379639,
12.4201984405518,44.2092514038086,
9.21033573150635,24.7096691131592,
-33.0578536987305,-3.99592661857605,
-69.3201065063477,-1.10419344902039,
-50.4308357238770,21.1589527130127,
0.684423446655273,19.2790412902832,
27.1782474517822,-17.8201961517334,
19.9556732177734,-57.8123092651367,
22.3055667877197,-58.7793045043945,
46.4115638732910,-17.8478450775147,
51.4982070922852,32.5149307250977,
9.87314510345459,51.2772979736328,
-41.8582763671875,26.0050964355469,
-54.7704124450684,-23.0222625732422,
-28.9749069213867,-58.7745056152344,
-5.60598659515381,-56.7439041137695,
-11.6836910247803,-31.9235439300537,
-28.5929145812988,-14.9305076599121,
-34.5011711120606,-10.9688367843628,
-31.1174736022949,2.05583310127258,
-32.1174163818359,25.1127452850342,
-38.0925025939941,26.7752475738525,
-39.1154251098633,-12.8792171478271,
-37.8032798767090,-59.9423294067383,
-33.3671188354492,-61.6577110290527,
-23.9756374359131,-15.4406147003174,
-15.8704948425293,20.1234226226807,
-18.5431461334229,4.47907304763794,
-28.3448429107666,-28.9316120147705,
-26.9836273193359,-26.1023445129395,
-7.34962415695190,15.1608581542969,
19.5131950378418,45.7149162292481,
33.5591354370117,36.3164062500000,
35.4011688232422,12.3930473327637,
35.2835464477539,3.15627527236938,
22.8754844665527,10.3172721862793,
-15.5660448074341,20.4786357879639,
-56.7248306274414,31.0690670013428,
-59.5670547485352,43.6844787597656,
-19.1737194061279,42.0946998596191,
15.4607887268066,12.3042945861816,
10.6432590484619,-28.7121391296387,
-9.24669742584229,-44.3829689025879,
-0.0631251931190491,-26.2599887847900,
26.5304660797119,-2.53410601615906,
21.3778915405273,3.91621351242065,
-23.7178268432617,0.390692591667175,
-49.7513580322266,-5.22488021850586,
-13.3623542785645,-15.2057428359985,
47.0811195373535,-23.2927665710449,
61.0686187744141,-13.4390716552734,
17.5137462615967,21.0781898498535,
-26.7414970397949,51.2087745666504,
-23.8194026947022,41.3645706176758,
9.71505451202393,0.0509522147476673,
32.4597473144531,-27.0110969543457,
32.4346847534180,-24.0184230804443,
22.3553581237793,-16.0043106079102,
15.3677635192871,-24.3946437835693,
9.02899074554443,-35.5824928283691,
2.52889466285706,-36.8350639343262,
6.98975753784180,-36.7988128662109,
25.9381561279297,-41.4976692199707,
38.5388526916504,-29.0755062103272,
25.3715686798096,17.2041435241699,
-11.0675086975098,59.7250938415527,
-43.2096939086914,44.4735984802246,
-42.2439880371094,-14.6092376708984,
-9.08528614044190,-42.0279502868652,
20.9693908691406,1.06361627578735,
17.6051349639893,55.1205329895020,
-10.3636322021484,44.5229339599609,
-27.3829135894775,-12.8039398193359,
-14.3245468139648,-44.5903015136719,
6.57104730606079,-27.8371200561523,
3.70191812515259,-11.6575622558594,
-18.1895465850830,-34.5298652648926,
-22.6730613708496,-65.2197341918945,
10.7166042327881,-54.7769012451172,
55.5598411560059,-9.79201412200928,
69.8914489746094,22.9274196624756,
47.5707893371582,23.1577167510986,
13.3167934417725,4.09878206253052,
-10.9722118377686,-18.8975334167480,
-20.4831695556641,-40.6944427490234,
-20.2912788391113,-41.5343742370606,
-9.86584663391113,-5.87200403213501,
0.585101842880249,39.2965850830078,
-5.35027456283569,53.9495315551758,
-29.9621009826660,35.9278717041016,
-47.5381393432617,24.0857429504395,
-36.7719879150391,36.3412284851074,
-10.8045835494995,42.2251701354981,
-1.91288042068481,9.14050292968750,
-10.7481842041016,-36.8345489501953,
-5.20903873443604,-44.5752716064453,
27.5134792327881,-16.3727741241455,
54.3379859924316,1.52435982227325,
38.2687225341797,-2.88147115707397,
-5.15049600601196,-3.20949292182922,
-29.9796161651611,8.06466293334961,
-24.6206684112549,3.30672264099121,
-20.0853519439697,-29.6494235992432,
-37.1391448974609,-59.1438484191895,
-51.7017326354981,-56.4446372985840,
-38.8724822998047,-44.5986976623535,
-13.9917755126953,-51.0334930419922,
-7.72323656082153,-54.9066276550293,
-14.0556688308716,-15.9429330825806,
-1.34572625160217,41.5359764099121,
29.1234703063965,48.6498031616211,
38.0121231079102,-6.64800643920898,
6.45429182052612,-50.4296951293945,
-35.1893920898438,-26.3534545898438,
-41.0726470947266,22.1503009796143,
-10.8116264343262,21.4724407196045,
19.9041748046875,-21.2139148712158,
32.4506187438965,-32.6274948120117,
38.6155700683594,18.5979156494141,
42.6390609741211,78.9451980590820,
39.8897590637207,82.0638427734375,
28.3684120178223,36.7705345153809,
20.9848594665527,1.77844452857971,
20.9674339294434,-0.947356283664703,
24.1247005462647,3.87726116180420,
28.3070011138916,-11.5979795455933,
36.2144889831543,-32.0128974914551,
36.7468681335449,-29.7108764648438,
5.08077669143677,-1.97254312038422,
-53.1886634826660,23.6762466430664,
-83.5394897460938,15.5255165100098,
-40.8775825500488,-24.2424297332764,
33.0335617065430,-55.6988334655762,
54.0822296142578,-43.9906082153320,
3.85134744644165,5.02214336395264,
-54.2575836181641,50.0378265380859,
-58.4156417846680,56.8701057434082,
-29.4541950225830,27.7042007446289,
-18.5464591979980,-4.95071792602539,
-27.3464107513428,-26.9740638732910,
-13.3976001739502,-37.8726577758789,
26.7404937744141,-36.8032493591309,
49.6855125427246,-15.7068109512329,
31.9451675415039,21.9473495483398,
11.0213003158569,50.8752365112305,
15.8135566711426,50.0314140319824,
19.5976543426514,27.0049514770508,
-13.0898303985596,3.38490867614746,
-55.9470939636231,-4.36689090728760,
-49.9118957519531,-0.186471343040466,
8.20227336883545,7.88152599334717,
57.9597091674805,19.7931137084961,
55.7128295898438,30.6737403869629,
19.6799468994141,38.2766799926758,
-1.25751066207886,41.6146507263184,
2.43362522125244,41.9973106384277,
14.3121623992920,31.5217342376709,
27.7114238739014,2.87963700294495,
42.3924560546875,-27.8100490570068,
44.7461013793945,-25.8478546142578,
21.4067153930664,24.2444534301758,
-9.66509342193604,79.6433639526367,
-18.7933921813965,81.1299667358398,
-4.82448053359985,19.4372100830078,
-1.45682728290558,-47.0695457458496,
-22.8081569671631,-51.2273483276367,
-46.8313636779785,2.14161133766174,
-48.0733299255371,52.3662643432617,
-35.8712654113770,54.8328247070313,
-37.6301574707031,22.7644481658936,
-50.5137596130371,-2.28674507141113,
-41.2486419677734,-4.71919393539429,
-1.61936950683594,4.09142255783081,
37.4212112426758,9.65864753723145,
41.5828323364258,7.78916120529175,
11.5403404235840,-9.08042335510254,
-18.5257205963135,-41.4097099304199,
-16.2611007690430,-67.3913116455078,
19.4477119445801,-56.5734786987305,
53.4794731140137,-8.63998985290527,
51.5995445251465,33.1743927001953,
13.5295162200928,25.7938289642334,
-26.7589874267578,-15.2527933120728,
-34.4070434570313,-40.8156585693359,
-14.8927698135376,-24.9963016510010,
-4.42007732391357,13.4906187057495,
-21.3379573822022,37.3116798400879,
-36.8611717224121,32.3190612792969,
-20.8303012847900,13.2611722946167,
12.8419561386108,-0.168586328625679,
17.1628932952881,3.09311866760254,
-13.3459739685059,20.4867515563965,
-38.6590385437012,29.6010475158691,
-23.1995792388916,6.67029237747192,
14.5717220306396,-34.3207435607910,
27.6193828582764,-45.9055747985840,
4.00215435028076,-9.58871650695801,
-22.8282318115234,24.7144298553467,
-27.5476760864258,4.58720922470093,
-15.8655843734741,-48.8586273193359,
-7.29461765289307,-67.5726318359375,
-5.25742292404175,-23.5429420471191,
-5.40514802932739,29.0215110778809,
-7.68814706802368,34.8219604492188,
-3.66630411148071,15.7427768707275,
19.6775112152100,18.5014877319336,
54.8075561523438,29.2067356109619,
64.0188598632813,8.23996353149414,
28.5670509338379,-26.6645336151123,
-21.7825660705566,-20.3658676147461,
-34.1233749389648,27.1519241333008,
2.06542181968689,49.7564086914063,
36.5540237426758,17.5546436309814,
30.1611003875732,-9.28896427154541,
-0.253742098808289,19.5389995574951,
-22.7624053955078,61.4639968872070,
-34.7029304504395,42.4359741210938,
-42.3931350708008,-18.8240947723389,
-37.0714225769043,-36.9432182312012,
-11.7412538528442,4.65538692474365,
13.2594881057739,28.1348419189453,
11.6667032241821,-8.31528186798096,
-2.51216030120850,-42.0877456665039,
11.7281179428101,-10.5750436782837,
47.0948867797852,46.8988189697266,
45.1231155395508,46.7710876464844,
-10.7722587585449,-9.30483245849609,
-56.3202514648438,-49.2675056457520,
-33.0315513610840,-35.5288467407227,
19.0681610107422,-13.9446229934692,
21.5084743499756,-28.5694770812988,
-23.2878227233887,-49.1403503417969,
-43.0156059265137,-27.2978744506836,
-12.1016969680786,22.9225330352783,
9.47117805480957,45.4737052917481,
-26.4344520568848,22.5558052062988,
-68.1065292358398,-10.4976119995117,
-41.2929878234863,-20.9431877136230,
29.9204597473145,-6.18692398071289,
56.9669990539551,9.68091773986816,
17.1841392517090,7.38476228713989,
-22.4824275970459,-15.0428905487061,
-14.0608549118042,-42.4781608581543,
8.66866970062256,-56.7085189819336,
2.09238386154175,-45.6329574584961,
-12.4618949890137,-19.0865364074707,
-0.816018581390381,-0.684135079383850,
16.0355300903320,0.583938360214233,
-6.40492486953735,-11.0144433975220,
-49.6009178161621,-25.5631179809570,
-46.8112258911133,-38.3481254577637,
13.9031276702881,-37.7419776916504,
56.0966987609863,-9.73775196075440,
21.1111412048340,33.8987770080566,
-47.2575759887695,63.3276290893555,
-60.1583251953125,57.6536941528320,
-8.14557552337647,28.6783866882324,
38.8358917236328,6.11078739166260,
25.6632099151611,5.94732904434204,
-22.1989898681641,19.8174858093262,
-43.8549652099609,29.7215843200684,
-22.1821517944336,22.1442337036133,
4.57921123504639,-3.07819223403931,
1.58126568794250,-35.6900634765625,
-20.5153350830078,-47.3095817565918,
-26.7406539916992,-20.3613834381104,
-8.69391632080078,30.7736167907715,
10.5472927093506,65.3768997192383,
5.95835304260254,53.6558074951172,
-23.2086143493652,7.98228645324707,
-49.7189483642578,-33.3408660888672,
-48.9135208129883,-48.0924224853516,
-25.7364044189453,-43.0735664367676,
3.38685250282288,-32.1331138610840,
28.9037570953369,-20.9616355895996,
43.2443389892578,-1.29251480102539,
37.2577857971191,20.1784515380859,
12.5447540283203,22.1472148895264,
-13.1484632492065,-7.21298456192017,
-11.0881252288818,-48.2742500305176,
23.2825260162354,-67.4132766723633,
54.3120117187500,-43.3704795837402,
43.2127532958984,7.69583034515381,
2.45329046249390,47.9567565917969,
-19.6789627075195,52.4214859008789,
-0.190777182579041,27.6491985321045,
26.3415241241455,1.02033460140228,
15.0064830780029,-8.41640853881836,
-25.6542434692383,-6.01573133468628,
-43.8289375305176,-11.9478683471680,
-22.0529575347900,-32.5716361999512,
-0.932512044906616,-41.1480484008789,
-16.9231319427490,-19.0579242706299,
-47.8208465576172,12.4570045471191,
-43.9754600524902,7.44284439086914,
-5.42407894134522,-37.0491409301758,
17.4890403747559,-66.7172393798828,
-8.23827934265137,-34.4154090881348,
-45.5793876647949,34.3601989746094,
-41.8432693481445,57.8585777282715,
-3.63851451873779,9.22001171112061,
21.3847293853760,-50.7864494323731,
8.21215057373047,-59.6894607543945,
-18.0724353790283,-21.4509277343750,
-18.7187194824219,15.1466636657715,
0.854665994644165,29.2536468505859,
0.653922796249390,38.6855735778809,
-30.5854816436768,45.6268539428711,
-57.4870300292969,33.2598152160645,
-44.2719383239746,7.26849937438965,
-0.816054105758667,7.03700733184814,
22.7597599029541,39.5925598144531,
-4.66890811920166,51.4142837524414,
-48.8775100708008,4.31547880172730,
-49.3029747009277,-57.8826942443848,
2.32575893402100,-55.7220230102539,
44.0299987792969,11.4527769088745,
20.6099681854248,62.1205139160156,
-45.7737236022949,40.0285568237305,
-74.3897628784180,-20.9663162231445,
-26.7070255279541,-59.0906448364258,
42.5632324218750,-55.4084625244141,
55.6440849304199,-36.2793464660645,
6.33733510971069,-16.4144134521484,
-37.8289146423340,11.1169824600220,
-32.0703048706055,33.1072654724121,
-6.75868320465088,23.3359127044678,
-10.1845388412476,-16.2351970672607,
-42.7893524169922,-44.5202407836914,
-59.3353118896484,-42.7541923522949,
-37.8915405273438,-32.1620903015137,
-7.39470577239990,-33.3696289062500,
0.560064077377319,-37.7761268615723,
-8.05218315124512,-40.6364364624023,
-14.0200386047363,-46.0492172241211,
-8.79918193817139,-51.7906913757324,
4.36268424987793,-42.2866210937500,
30.0588703155518,-6.45100164413452,
59.5937995910645,30.5781440734863,
56.6131439208984,38.0609588623047,
4.73651885986328,35.5997543334961,
-48.5543785095215,50.3549842834473,
-44.9449157714844,60.9358901977539,
5.76421594619751,21.6144065856934,
34.6969108581543,-46.1983108520508,
3.48378229141235,-63.4372825622559,
-37.9022560119629,-5.93016481399536,
-25.5756034851074,44.4381980895996,
24.5017490386963,14.5730304718018,
50.5813331604004,-49.6699104309082,
43.2859954833984,-47.2926406860352,
39.7872810363770,28.9979476928711,
53.7266387939453,75.5065002441406,
52.8383941650391,30.2798156738281,
23.5734252929688,-45.7992591857910,
2.31680750846863,-61.5674934387207,
13.3176784515381,-22.1082267761230,
20.1954059600830,-3.04059767723084,
-10.0842494964600,-26.0109939575195,
-47.8808250427246,-41.2994804382324,
-38.7673301696777,-7.60183763504028,
5.92791128158569,40.7854194641113,
11.6127243041992,54.4917259216309,
-41.2057991027832,28.3661594390869,
-79.2364883422852,-6.55292844772339,
-42.3042449951172,-26.3253860473633,
34.7275886535645,-37.9100341796875,
72.4395370483398,-48.9153633117676,
46.1534690856934,-46.1195449829102,
1.44829440116882,-19.6289024353027,
-19.8424453735352,12.9675855636597,
-14.2274951934814,31.5350608825684,
1.81106925010681,30.2809028625488,
21.6462802886963,26.3052177429199,
30.7457160949707,38.7785034179688,
7.74483489990234,57.5762481689453,
-34.4692001342773,50.0794486999512,
-49.1514625549316,8.07678031921387,
-18.2870540618897,-30.4906692504883,
11.5567808151245,-24.7593345642090,
-0.572913885116577,16.2871799468994,
-35.8718490600586,40.4666442871094,
-39.5553703308106,19.1251010894775,
-5.65658712387085,-12.9411983489990,
22.5023708343506,-4.65294027328491,
20.1580543518066,37.8579559326172,
12.5607500076294,62.9608078002930,
23.4010219573975,43.2238883972168,
28.3673553466797,9.73798370361328,
1.27462029457092,4.97115468978882,
-33.4116477966309,31.0649566650391,
-33.9736289978027,51.5437240600586,
-9.79490661621094,44.2364616394043,
-8.35894012451172,15.5646047592163,
-38.9793090820313,-14.9369955062866,
-50.7204170227051,-35.2352828979492,
-8.49693107604981,-38.4000091552734,
55.3519554138184,-21.2368164062500,
75.0397872924805,8.49509906768799,
33.1233825683594,33.2366828918457,
-22.4739723205566,39.4688034057617,
-41.4353561401367,22.8994483947754,
-21.6818199157715,-3.15224647521973,
8.86205101013184,-21.4753742218018,
26.5786075592041,-20.1127891540527,
25.5250549316406,4.09590339660645,
7.78603887557983,29.6256561279297,
-16.8131828308105,31.5985031127930,
-33.5117950439453,5.73623514175415,
-35.5620346069336,-26.4332675933838,
-29.0058879852295,-42.2490806579590,
-25.7826347351074,-38.2704315185547,
-31.2063102722168,-33.9295501708984,
-37.8257942199707,-40.8501510620117,
-35.6704216003418,-46.6395874023438,
-27.7494087219238,-42.0616645812988,
-21.9435997009277,-33.3822631835938,
-16.2872238159180,-35.5018463134766,
-6.99020862579346,-44.7263221740723,
8.62594795227051,-31.7887382507324,
26.4925727844238,12.5500240325928,
30.1500110626221,57.4982910156250,
10.3470439910889,55.7440452575684,
-17.9278450012207,8.13566875457764,
-24.2376003265381,-33.9475479125977,
4.29778051376343,-26.0867214202881,
42.0243835449219,13.8278617858887,
52.0199050903320,27.9952259063721,
25.7731933593750,-8.33427524566650,
-2.00026774406433,-56.2910728454590,
-2.97169589996338,-66.6275558471680,
8.16428661346436,-38.1766128540039,
-1.14869832992554,-13.1199064254761,
-21.1589603424072,-17.1245098114014,
-14.6063480377197,-37.9832992553711,
26.9655284881592,-44.7508354187012,
55.2488784790039,-34.1002540588379,
29.2002391815186,-24.8257560729980,
-25.9243640899658,-28.7930068969727,
-46.9239234924316,-38.6134567260742,
-21.1153697967529,-39.7659568786621,
3.87861323356628,-29.9357852935791,
-9.46132087707520,-15.9735574722290,
-33.0363807678223,-4.90171527862549,
-22.4571685791016,9.59002971649170,
12.1702690124512,29.7594261169434,
20.0515804290772,37.8488616943359,
-12.8499774932861,17.4833602905273,
-44.4482192993164,-19.0582160949707,
-37.0927963256836,-39.2615966796875,
-4.67558002471924,-16.3028030395508,
14.1368570327759,27.1618270874023,
8.34549999237061,38.3691482543945,
1.58471333980560,-2.99985384941101,
11.8961105346680,-52.8034248352051,
36.0637016296387,-60.0310707092285,
57.2734985351563,-33.0968208312988,
65.4279251098633,-21.5623073577881,
53.7322959899902,-42.3238372802734,
21.1011810302734,-50.1629066467285,
-14.2601623535156,-8.08897304534912,
-31.2528266906738,43.8577957153320,
-27.2088928222656,38.1779632568359,
-18.5554027557373,-21.5945816040039,
-15.0166568756104,-57.2401847839356,
-14.5392894744873,-25.1555404663086,
-10.2419185638428,27.1133213043213,
-7.19983148574829,34.8723144531250,
-16.6654624938965,5.18535614013672,
-34.2330360412598,-8.99365520477295,
-45.7070350646973,2.29708480834961,
-42.5487060546875,-5.74567461013794,
-24.9800987243652,-44.3982696533203,
7.51197052001953,-63.7465820312500,
44.7264289855957,-28.4234275817871,
62.9254989624023,30.3216342926025,
49.0578041076660,52.3892288208008,
21.9076404571533,32.4675865173340,
19.5700988769531,11.0231151580811,
47.2637252807617,6.51252794265747,
67.6799163818359,-3.28928494453430,
48.5320281982422,-20.7269420623779,
10.5320997238159,-20.1663150787354,
-0.962005496025085,5.12884521484375,
28.1264495849609,26.6480140686035,
57.8330345153809,13.0454607009888,
54.5098762512207,-24.9280300140381,
33.6981391906738,-44.1490516662598,
27.9509582519531,-27.7767333984375,
38.8448143005371,4.39949131011963,
42.0209770202637,30.1421127319336,
18.3989048004150,39.2549591064453,
-20.6073303222656,33.5339012145996,
-45.7893524169922,20.2601127624512,
-38.0805435180664,23.3377361297607,
-5.84689140319824,47.6039161682129,
22.7866973876953,64.1269989013672,
12.4967966079712,37.4854011535645,
-40.7480773925781,-18.6874122619629,
-87.0986633300781,-49.3822860717773,
-68.9764175415039,-27.9665107727051,
-3.02217674255371,6.26861143112183,
32.9066390991211,1.12246584892273,
0.363946914672852,-33.8963508605957,
-42.7727127075195,-43.6387481689453,
-28.2019290924072,-6.13499069213867,
24.4433593750000,36.2528152465820,
29.4339694976807,44.7300300598145,
-29.0005226135254,27.8132934570313,
-67.7783279418945,16.8861312866211,
-24.0892601013184,18.3921756744385,
44.8423995971680,18.6042861938477,
42.7889175415039,12.4657363891602,
-27.3953437805176,11.6943302154541,
-70.4543151855469,15.3564596176147,
-37.8987503051758,14.4899301528931,
16.2465591430664,3.33988404273987,
22.3370742797852,-10.4755945205688,
-4.31753110885620,-23.8583126068115,
-13.0401773452759,-42.9295043945313,
8.31671810150147,-58.6509628295898,
20.6851177215576,-50.7259140014648,
3.29320359230042,-17.0225086212158,
-17.9025535583496,9.30587673187256,
-16.4752788543701,10.8599348068237,
-1.49956846237183,5.95315885543823,
6.32527923583984,20.2327079772949,
6.28975248336792,50.5158805847168,
1.77186274528503,64.4342575073242,
-12.1533927917480,49.3284568786621,
-30.3121509552002,28.7033329010010,
-39.8689498901367,23.9766387939453,
-41.0283164978027,25.5508365631104,
-45.9122886657715,19.0004997253418,
-61.4676742553711,7.20344066619873,
-69.5047988891602,-7.53015899658203,
-45.7033843994141,-30.5368881225586,
-2.68559217453003,-55.1875724792481,
20.0989589691162,-52.8977241516113,
11.6970624923706,-4.15938901901245,
-5.50499820709229,50.3499603271484,
-13.2997322082520,49.8137207031250,
-18.6387634277344,-5.23759078979492,
-27.3026485443115,-46.7356986999512,
-29.2066535949707,-22.3600387573242,
-19.0743331909180,28.0018577575684,
-14.5931825637817,28.0638141632080,
-29.8220863342285,-27.8253974914551,
-40.5841484069824,-63.2440681457520,
-15.4794445037842,-27.3109760284424,
34.6543693542481,39.7367897033691,
52.8635520935059,62.5475616455078,
11.5574016571045,21.1130828857422,
-52.6699256896973,-33.8160095214844,
-74.3144607543945,-45.3400268554688,
-43.8784408569336,-14.1238136291504,
0.902838349342346,18.8458690643311,
25.3351478576660,16.3512153625488,
25.7315387725830,-19.9507598876953,
19.1419067382813,-57.4262237548828,
11.8540468215942,-60.8598861694336,
3.50613498687744,-25.5604190826416,
-6.06541347503662,11.1261072158813,
-14.2266426086426,14.0622053146362,
-21.2411670684814,-7.23351764678955,
-22.8149967193604,-12.0732288360596,
-16.5316066741943,4.50147533416748,
-11.0140399932861,12.1954154968262,
-23.4617862701416,-15.1092462539673,
-54.6429252624512,-49.6355590820313,
-67.6689605712891,-44.6473922729492,
-36.5969543457031,-4.42452001571655,
13.6736955642700,26.0233230590820,
36.8342666625977,24.6359920501709,
11.6039247512817,18.7519359588623,
-29.3588256835938,31.8770332336426,
-49.0039482116699,43.8194961547852,
-45.5780563354492,23.0818214416504,
-42.6486854553223,-19.7678127288818,
-47.6509323120117,-46.6049270629883,
-49.3408050537109,-46.0510940551758,
-41.0910873413086,-43.6747016906738,
-24.1183738708496,-57.4283103942871,
5.89647006988525,-73.1932601928711,
43.8816108703613,-66.0455245971680,
63.9476776123047,-34.8382339477539,
39.9208679199219,5.13951683044434,
-15.3673620223999,44.2780342102051,
-52.6814956665039,68.3064422607422,
-50.6207542419434,59.7563133239746,
-37.1862983703613,26.8942928314209,
-46.2335472106934,6.34816312789917,
-61.9063491821289,21.0129051208496,
-40.8570938110352,42.8082389831543,
10.4038887023926,22.6888465881348,
37.6865234375000,-31.5522384643555,
17.0858535766602,-65.0957260131836,
-8.11759662628174,-45.5743980407715,
7.89536762237549,-9.30220031738281,
46.4033813476563,-8.76181411743164,
58.2728271484375,-30.6567287445068,
29.7201271057129,-20.1979045867920,
-0.392773270606995,34.0537872314453,
-5.39069938659668,78.5051498413086,
1.30146765708923,59.0938072204590,
-3.54105210304260,-6.62902975082398,
-8.32221126556397,-50.5870742797852,
8.62258148193359,-35.4725837707520,
36.3908424377441,15.9518766403198,
51.4152526855469,45.9379615783691,
40.5157241821289,27.9912509918213,
11.2453632354736,-15.1175384521484,
-28.1836662292480,-40.1426086425781,
-60.7973442077637,-29.4611434936523,
-59.6526756286621,0.673692643642426,
-16.3053493499756,22.0000762939453,
33.9082183837891,20.8248882293701,
40.8379440307617,10.2478275299072,
6.21469497680664,3.77628040313721,
-12.8522272109985,-5.70951366424561,
14.4085140228271,-20.5076942443848,
49.8789482116699,-24.3313121795654,
37.0371475219727,-4.99300861358643,
-15.7888154983521,27.4609966278076,
-51.0317993164063,41.4295158386231,
-42.6439933776856,18.1742687225342,
-25.9814262390137,-20.3396434783936,
-33.6912307739258,-42.4358406066895,
-50.4514732360840,-42.6258926391602,
-36.7416915893555,-31.6285762786865,
3.70932435989380,-15.5305500030518,
27.6390018463135,5.76869201660156,
11.4777536392212,20.0063457489014,
-21.0627079010010,4.80356693267822,
-25.3200130462647,-36.4862098693848,
4.54431390762329,-62.5805015563965,
39.1659584045410,-41.4224472045898,
52.6880378723145,6.40193653106689,
39.9311485290527,26.4294853210449,
19.9611186981201,1.01953744888306,
15.6120500564575,-32.8785095214844,
25.4841403961182,-30.8466415405273,
34.4161872863770,3.28969812393188,
29.9185733795166,26.5306682586670,
9.82636070251465,19.8090400695801,
-13.6196260452271,1.94692933559418,
-31.4947471618652,-6.71548175811768,
-37.3404426574707,-5.48596906661987,
-26.2374763488770,-9.13863277435303,
6.86140823364258,-16.8194236755371,
46.7035865783691,-16.5593185424805,
55.4995574951172,-6.32371950149536,
14.7966432571411,2.15062165260315,
-41.3824882507324,-3.43871498107910,
-55.9560737609863,-21.3030834197998,
-10.1938610076904,-36.0744705200195,
48.2509880065918,-31.9061927795410,
60.4246482849121,-1.93359375000000,
23.3398704528809,32.6668739318848,
-17.8157463073730,37.4205017089844,
-27.4687767028809,6.11544084548950,
-14.0471305847168,-30.3738632202148,
-3.38877820968628,-31.6202449798584,
-0.0761609971523285,2.00452709197998,
3.97759866714478,28.1621589660645,
6.32585716247559,19.2136249542236,
-1.20809864997864,-6.93596076965332,
-12.9836568832397,-15.9877262115479,
-12.7416210174561,-6.24018192291260,
2.18953990936279,-2.12934374809265,
10.8721284866333,-7.74142408370972,
-1.01246643066406,-1.10572040081024,
-24.8552265167236,27.6927394866943,
-42.4293212890625,50.0964851379395,
-45.6057968139648,31.1724319458008,
-41.7051239013672,-19.8410758972168,
-32.9553375244141,-59.1709060668945,
-18.7150268554688,-57.0428276062012,
-0.224198579788208,-21.9559745788574,
15.4181585311890,17.2735176086426,
23.2934741973877,41.1521530151367,
24.4312648773193,50.4965209960938,
15.9277057647705,45.1524085998535,
-2.10535120964050,24.4626903533936,
-22.6803131103516,0.0281802415847778,
-31.5449981689453,-10.3563642501831,
-18.4126663208008,0.702982485294342,
6.55020236968994,20.9422950744629,
22.0335903167725,24.7034893035889,
18.1655788421631,5.37113094329834,
3.59927654266357,-18.8472900390625,
-7.46162700653076,-21.3695640563965,
2.19535017013550,-5.01259517669678,
27.3761787414551,6.68577003479004,
43.8912811279297,-6.10889244079590,
25.6137390136719,-34.5319366455078,
-24.0337524414063,-47.5010795593262,
-64.9627532958984,-34.4589843750000,
-56.0787849426270,-15.0916223526001,
-6.88846063613892,-14.4117612838745,
24.1314353942871,-29.2108879089355,
2.60375499725342,-29.5941276550293,
-41.2138023376465,-1.70377683639526,
-46.5857276916504,34.1944427490234,
-2.96191525459290,48.4166526794434,
29.5561752319336,34.8930244445801,
0.725875854492188,21.4460906982422,
-60.7967376708984,28.0379791259766,
-81.2503738403320,44.3963508605957,
-32.7230606079102,47.4959869384766,
32.4190063476563,29.0565109252930,
43.2732200622559,2.92527222633362,
-1.78954458236694,-18.1027297973633,
-41.3176765441895,-32.0534210205078,
-24.0075778961182,-40.6911544799805,
32.3271484375000,-34.3757591247559,
68.0995788574219,-12.4104766845703,
54.2845001220703,11.3361740112305,
13.5821075439453,23.3832054138184,
-6.56791353225708,25.8492717742920,
7.43040180206299,35.1118469238281,
24.2132148742676,55.5799179077148,
10.5526514053345,69.3247070312500,
-16.5051536560059,54.7459907531738,
-17.1582298278809,19.3459873199463,
17.3924598693848,-12.7629747390747,
49.1420898437500,-22.0699176788330,
38.0170440673828,-13.5909061431885,
3.32132244110107,-11.5676012039185,
-0.246729254722595,-26.9293689727783,
28.0323829650879,-39.2961692810059,
35.1268539428711,-22.2452430725098,
-7.14396047592163,26.3482379913330,
-54.9303817749023,69.0956954956055,
-51.5483474731445,68.5570831298828,
-6.26976108551025,28.8228607177734,
18.3534297943115,-10.0559072494507,
8.40960502624512,-17.3317222595215,
7.87463712692261,-10.4563159942627,
40.6396980285645,-20.7584934234619,
61.0896987915039,-43.0177650451660,
24.7595329284668,-42.2642364501953,
-32.4728736877441,-11.0575084686279,
-35.5739784240723,16.7730484008789,
21.9793319702148,5.29483127593994,
70.6102828979492,-30.8149719238281,
62.9381103515625,-52.5420989990234,
22.2740058898926,-40.2352867126465,
-0.574677348136902,-12.1544065475464,
4.51879692077637,14.9483718872070,
19.4283523559570,42.9767303466797,
35.3366546630859,65.9173431396484,
46.3639030456543,65.6913986206055,
38.8517112731934,40.5615005493164,
7.39189338684082,23.5403556823730,
-20.4028110504150,34.8474617004395,
-7.55356597900391,53.0393524169922,
24.5721530914307,44.2139511108398,
19.2808322906494,14.2090015411377,
-31.5465965270996,-4.92030334472656,
-66.9968109130859,-11.6034679412842,
-36.4130516052246,-32.0590972900391,
32.6494865417481,-66.1966018676758,
72.7921371459961,-65.5034255981445,
50.8195991516113,-5.67634820938110,
-1.31062674522400,53.6644363403320,
-38.8093376159668,45.9352340698242,
-39.8274078369141,-13.0026397705078,
-6.08988571166992,-43.2715911865234,
39.8292999267578,-8.85675525665283,
57.4721031188965,38.3358726501465,
19.4869441986084,41.9651451110840,
-46.1593284606934,6.84222221374512,
-68.5562057495117,-22.1519832611084,
-21.6252975463867,-27.1820507049561,
43.1672935485840,-20.7580928802490,
62.8041877746582,-7.16469383239746,
34.1334953308106,18.8205966949463,
2.34752130508423,36.7996025085449,
-2.67350006103516,18.4420375823975,
5.55244922637939,-24.8584537506104,
8.63279151916504,-46.5785064697266,
8.34243774414063,-30.8270587921143,
1.32518231868744,-8.75672054290772,
-24.6745109558105,-5.59415531158447,
-51.4352035522461,-9.93509769439697,
-41.9839591979981,-2.94764709472656,
8.57054328918457,4.78890180587769,
45.6356582641602,-11.6030063629150,
19.2074146270752,-36.9928550720215,
-35.9583091735840,-32.2693786621094,
-42.8055801391602,1.82427430152893,
6.77092885971069,22.5125408172607,
44.1643638610840,11.7447080612183,
14.2559852600098,-4.07532501220703,
-48.9907188415527,2.04799532890320,
-66.9786987304688,15.7561674118042,
-31.6588973999023,11.4278383255005,
-3.88271951675415,1.03696155548096,
-22.8473186492920,3.60679841041565,
-59.9900817871094,10.4098844528198,
-64.6709213256836,-6.03290557861328,
-29.2124252319336,-41.8699798583984,
8.18829154968262,-57.1600875854492,
16.8510189056397,-36.2969093322754,
0.499042391777039,-18.0119495391846,
-11.5958585739136,-34.4725112915039,
4.03684806823731,-59.5682868957520,
35.8182868957520,-47.9199409484863,
51.3386383056641,-0.0425820350646973,
25.3977737426758,38.3386077880859,
-29.9018611907959,33.1563873291016,
-64.8862838745117,-4.41981315612793,
-44.4431304931641,-41.1465873718262,
3.66777276992798,-54.5108108520508,
27.5098037719727,-36.3580932617188,
12.9625902175903,7.20285081863403,
-10.9808616638184,45.6741180419922,
-16.6842670440674,39.5043525695801,
-7.80739212036133,-8.23665142059326,
2.07875061035156,-43.5971565246582,
16.0083160400391,-21.9469890594482,
34.5356903076172,30.7934265136719,
35.3172836303711,51.6141433715820,
0.283967375755310,20.9819297790527,
-39.9062690734863,-13.9932346343994,
-36.2393836975098,-14.7116174697876,
4.53773736953735,8.82788085937500,
23.0490036010742,14.7837314605713,
-11.9797182083130,-1.74123334884644,
-55.1602249145508,-11.1111993789673,
-48.9330329895020,-0.448510706424713,
-2.63466882705688,9.23018360137940,
32.4224090576172,-4.19141006469727,
36.0791816711426,-30.3988380432129,
35.2399368286133,-34.6037216186523,
38.6455001831055,-7.02141952514648,
19.1454963684082,31.1997165679932,
-29.0594520568848,41.1765670776367,
-56.1897010803223,7.37390804290772,
-25.0722503662109,-48.0947036743164,
28.9545860290527,-82.0161972045898,
46.5559806823731,-71.3093566894531,
26.9828987121582,-25.9230041503906,
16.7572021484375,23.7044181823730,
28.8770523071289,47.6706123352051,
28.4718589782715,39.2774543762207,
-2.86753320693970,9.34770011901856,
-28.7071933746338,-20.4528160095215,
-13.5914592742920,-29.6118450164795,
23.8953189849854,-5.96666336059570,
39.1196899414063,33.8603591918945,
32.8218574523926,60.0124130249023,
33.6357307434082,58.6612243652344,
38.0352554321289,46.8727607727051,
16.9600753784180,44.4954414367676,
-25.9524593353272,45.2935714721680,
-47.2274475097656,22.6667480468750,
-23.8904113769531,-27.4082508087158,
14.4598913192749,-67.7225189208984,
28.7762222290039,-64.7993774414063,
18.0263862609863,-25.4008522033691,
10.2945709228516,9.31560897827148,
13.2015686035156,20.8834533691406,
13.5894298553467,28.2063598632813,
11.8911285400391,47.8221626281738,
18.5472850799561,64.6318206787109,
21.0120811462402,59.6260337829590,
-2.71055746078491,39.8521003723145,
-44.5917434692383,32.2823410034180,
-61.0521163940430,38.8633613586426,
-31.1574020385742,30.8523941040039,
12.6705379486084,-3.90773773193359,
32.8677368164063,-34.3064270019531,
27.3248291015625,-29.5009956359863,
20.3812732696533,0.0962589308619499,
19.8043251037598,14.9837217330933,
8.90530776977539,-0.605577230453491,
-12.7447566986084,-24.1045036315918,
-15.6717586517334,-33.6991004943848,
10.2860984802246,-22.2202529907227,
35.9783554077148,4.68909645080566,
26.7189292907715,43.9769706726074,
-14.1373558044434,76.4449234008789,
-54.4141311645508,66.9755935668945,
-64.8181991577148,10.1865806579590,
-40.7022171020508,-52.6055526733398,
4.06754589080811,-67.3588409423828,
41.0644874572754,-33.3614387512207,
47.8158950805664,1.21551156044006,
20.1844882965088,4.69300508499146,
-8.85331916809082,-4.75936079025269,
-0.999466896057129,-5.68347549438477,
35.8658714294434,1.33999109268188,
58.6987915039063,2.06041002273560,
44.7535552978516,3.79124283790588,
20.0848407745361,25.1131019592285,
15.5862255096436,61.3035697937012,
18.2116107940674,76.1106796264648,
1.34111142158508,48.6906127929688,
-25.8833332061768,0.0176427364349365,
-26.6509494781494,-35.1094474792481,
2.41482710838318,-36.9895782470703,
19.7781734466553,-10.8560867309570,
-7.44034242630005,16.2328910827637,
-50.6443672180176,9.04782390594482,
-58.6147918701172,-38.0879058837891,
-23.2058982849121,-85.5425567626953,
14.2948074340820,-84.2217407226563,
23.9929466247559,-36.8227691650391,
7.35105371475220,-5.24664258956909,
-18.6857128143311,-27.0076198577881,
-36.4499244689941,-57.8493957519531,
-31.3879833221436,-34.8857841491699,
-2.25441527366638,25.6266536712647,
31.5273265838623,42.2665443420410,
45.0159759521484,-6.90044784545898,
40.1180610656738,-42.0536918640137,
40.7243804931641,-2.08150529861450,
50.1788825988770,68.5030822753906,
34.2699661254883,72.5165023803711,
-19.2920265197754,1.53050041198730,
-59.4272766113281,-54.0600700378418,
-30.9884262084961,-34.1431617736816,
36.7745933532715,21.2021102905273,
61.1814613342285,44.1311073303223,
13.2103385925293,23.0287532806397,
-48.1471328735352,-2.89405369758606,
-57.9223785400391,-20.6542110443115,
-29.0505237579346,-42.1226844787598,
-17.3923015594482,-55.0074195861816,
-31.4743385314941,-27.9573001861572,
-36.1765785217285,25.3589305877686,
-18.4071159362793,47.7731857299805,
-11.6444301605225,6.36721801757813,
-32.8497619628906,-60.5065956115723,
-47.5251464843750,-85.6156387329102,
-30.9474601745605,-48.9627304077148,
-0.542348623275757,6.31067657470703,
10.8214864730835,27.9545707702637,
10.0611619949341,12.4084577560425,
19.7196083068848,-16.4358482360840,
31.7466602325439,-27.4010715484619,
22.0675277709961,-9.38227367401123,
-7.54333972930908,17.3219184875488,
-24.0580215454102,25.2667732238770,
-18.5007095336914,3.36357259750366,
-22.8627834320068,-27.1332283020020,
-44.5452651977539,-36.3558540344238,
-47.7894134521484,-19.3567199707031,
-6.92323493957520,3.53254652023315,
34.8891983032227,13.7428760528564,
23.3262329101563,11.9759359359741,
-32.7042388916016,6.70568943023682,
-65.6054611206055,-0.994703173637390,
-39.9231033325195,-20.2871093750000,
13.2290039062500,-41.5049133300781,
41.7701148986816,-47.0619087219238,
38.1785240173340,-26.2653865814209,
27.4165172576904,10.3355216979980,
20.4257717132568,38.0349006652832,
7.17447471618652,43.1942634582520,
-10.0843610763550,34.1769332885742,
-24.3319778442383,31.2794532775879,
-37.9182319641113,41.5821838378906,
-52.9190483093262,44.0283050537109,
-53.9114990234375,15.4523401260376,
-24.6141433715820,-29.3431262969971,
17.8762817382813,-48.9947929382324,
40.8888549804688,-18.8907604217529,
33.7352752685547,36.2523345947266,
22.0815048217773,62.9490585327148,
24.8454246520996,42.5305671691895,
23.7782096862793,9.60974502563477,
0.925805985927582,-0.367312818765640,
-18.1392230987549,8.32383155822754,
1.07469415664673,8.23234176635742,
41.0709495544434,-6.33795547485352,
55.1715698242188,-12.4854621887207,
33.7605705261231,2.89177989959717,
14.5089120864868,13.9816274642944,
19.5382041931152,-2.80512452125549,
23.3892726898193,-32.8756523132324,
0.468543410301209,-37.2264595031738,
-20.8786334991455,-18.0546035766602,
-3.07151579856873,-13.9200096130371,
37.3443412780762,-41.7329559326172,
45.6041641235352,-59.5979461669922,
7.02628898620606,-24.3730869293213,
-29.1419849395752,38.2602882385254,
-30.0979652404785,57.0172004699707,
-19.2751178741455,12.4374246597290,
-32.7415771484375,-39.9962654113770,
-54.6081390380859,-41.7145767211914,
-46.7265739440918,-5.78851890563965,
-11.3143224716187,18.4750633239746,
13.5498685836792,18.8285636901855,
5.45427703857422,20.6809215545654,
-12.2305889129639,32.7560348510742,
-9.61257457733154,40.0145492553711,
11.5905570983887,38.0037384033203,
27.3581829071045,44.7621498107910,
32.5485610961914,55.4558982849121,
32.9201393127441,43.7256622314453,
27.5609111785889,4.11370277404785,
11.1597204208374,-22.9208297729492,
-10.0627574920654,-7.70341777801514,
-28.6336765289307,19.8587894439697,
-37.7027816772461,10.7992925643921,
-31.2394294738770,-25.2571525573730,
-10.4590845108032,-31.8036251068115,
12.1993017196655,1.67837619781494,
12.7225313186646,24.7894401550293,
-14.1572818756104,3.61699438095093,
-32.4941596984863,-36.6679916381836,
-5.23375129699707,-51.2353782653809,
49.8381958007813,-41.4902153015137,
73.8306808471680,-36.4350280761719,
45.8889923095703,-39.9307746887207,
13.0598583221436,-31.2327556610107,
21.0861835479736,-16.0070686340332,
50.3285751342773,-18.2442855834961,
43.7423744201660,-39.5356864929199,
-3.46786355972290,-42.1761093139648,
-34.0880432128906,-12.2289419174194,
-9.67953014373779,12.5235967636108,
34.9720840454102,-2.18225193023682,
39.7820777893066,-31.4090671539307,
-0.353192329406738,-26.9180526733398,
-35.4167633056641,14.9350452423096,
-32.5256958007813,46.0663032531738,
-9.40703487396240,32.2556915283203,
1.15370297431946,-9.21376132965088,
-1.36079037189484,-30.3816623687744,
2.95109820365906,-17.5830421447754,
13.7665605545044,12.1548395156860,
17.1235294342041,36.5345611572266,
1.31732273101807,46.3203620910645,
-19.9827213287354,39.4387130737305,
-26.1287288665772,22.6478519439697,
-13.2247400283813,8.58301448822022,
0.588315606117249,2.66868448257446,
1.03727054595947,-2.10224676132202,
-12.6353225708008,-12.9634313583374,
-31.3763504028320,-24.3771781921387,
-39.1671943664551,-26.5496253967285,
-31.2749404907227,-27.9347858428955,
-20.1678848266602,-42.9912757873535,
-9.26661014556885,-67.6928482055664,
7.43584346771240,-71.6306610107422,
34.7220726013184,-37.0163078308106,
53.2033157348633,8.49615287780762,
39.2738914489746,26.4254016876221,
-0.207664489746094,11.8966293334961,
-25.8953456878662,2.09745860099793,
-9.36431884765625,25.1298599243164,
20.6593036651611,57.4024658203125,
20.6038246154785,59.0841026306152,
-3.13130187988281,19.9896354675293,
-3.43793678283691,-21.6521415710449,
33.1917839050293,-22.7718505859375,
56.6432037353516,13.7849197387695,
23.7879543304443,46.2875785827637,
-37.7331275939941,38.9448165893555,
-67.5323181152344,-0.0752789974212647,
-52.4845657348633,-36.2498245239258,
-34.1038894653320,-44.9600028991699,
-36.9117965698242,-37.5161972045898,
-29.7087478637695,-36.2264099121094,
11.3653297424316,-34.7266540527344,
57.2166023254395,-10.3040428161621,
63.3502731323242,30.2820510864258,
35.5835227966309,51.7520523071289,
13.4239091873169,32.4579010009766,
12.9104700088501,3.54474973678589,
18.4072399139404,11.1977500915527,
23.2237777709961,57.3663177490234,
32.7604141235352,84.1246795654297,
36.1721801757813,54.9067115783691,
6.71936702728272,7.06901264190674,
-46.5568084716797,1.88056063652039,
-69.5453491210938,33.8180503845215,
-31.0940189361572,43.9044227600098,
25.9152107238770,6.00862789154053,
35.2964935302734,-30.2090644836426,
-2.77432489395142,-13.7031688690186,
-26.1233367919922,35.2674598693848,
-2.98075819015503,50.9775810241699,
30.4544811248779,24.0969409942627,
33.0493011474609,6.58598804473877,
12.6548824310303,24.8666477203369,
6.86096763610840,44.0610694885254,
20.8107509613037,25.2707328796387,
22.5940303802490,-7.63178157806397,
0.512819766998291,-16.6007061004639,
-16.2410736083984,-12.7284908294678,
0.146882057189941,-29.6234741210938,
35.9678726196289,-54.0740089416504,
47.7301177978516,-42.5799980163574,
17.0496883392334,5.44295692443848,
-24.7902755737305,28.4110698699951,
-40.6458015441895,-4.24461936950684,
-20.9135837554932,-48.1390419006348,
7.02567100524902,-45.7753219604492,
14.6408243179321,-8.22376823425293,
1.00027775764465,17.1746177673340,
-18.2239227294922,23.6731777191162,
-39.2130432128906,35.3086929321289,
-57.5940284729004,45.5397720336914,
-58.6409416198731,16.9686431884766,
-25.9067344665527,-40.9914321899414,
24.8293952941895,-66.7969284057617,
52.5014686584473,-28.7695770263672,
39.0531425476074,24.3104648590088,
13.4109001159668,20.0209331512451,
16.7638015747070,-34.0787086486816,
40.9493560791016,-68.6830902099609,
38.6843872070313,-47.2310371398926,
-0.642761707305908,-8.78326320648193,
-32.8884201049805,-0.569998860359192,
-16.7121791839600,-19.9460430145264,
31.3028869628906,-35.0434913635254,
57.1693458557129,-23.8424720764160,
43.2712097167969,7.19526386260986,
21.7341957092285,33.9303779602051,
19.9412803649902,36.1846923828125,
19.4289474487305,3.99862813949585,
-10.6446475982666,-40.7579574584961,
-51.5162124633789,-55.4902000427246,
-52.6422958374023,-20.6861572265625,
-4.92651796340942,30.6359100341797,
38.9187088012695,45.6149826049805,
26.7109146118164,16.9998416900635,
-21.4395446777344,-9.28514385223389,
-40.4153404235840,-1.69686222076416,
-7.15140533447266,18.1132564544678,
32.3519630432129,15.0976572036743,
34.3831214904785,-7.69693040847778,
13.7783927917480,-9.29036521911621,
8.75435638427734,24.5518779754639,
18.7692489624023,56.7927017211914,
18.5182151794434,46.5394287109375,
12.5781650543213,1.70136404037476,
22.6000633239746,-27.5232772827148,
39.2816810607910,-10.6551494598389,
23.8036708831787,24.8172149658203,
-23.5376434326172,30.3277263641357,
-45.5845832824707,0.285285234451294,
-11.0283355712891,-33.2354125976563,
33.8910255432129,-39.2263259887695,
30.2039031982422,-22.2758865356445,
-3.58525562286377,-10.8213596343994,
-0.216372251510620,-7.95424604415894,
40.7377700805664,7.03858661651611,
48.0622863769531,34.7310600280762,
-5.11126518249512,46.0696945190430,
-54.1444931030273,18.6296958923340,
-36.8684921264648,-24.7220172882080,
16.2934265136719,-39.3643531799316,
31.3376884460449,-13.1993598937988,
0.385361194610596,7.61734485626221,
-18.9746894836426,-16.8353214263916,
2.66055321693420,-60.0699234008789,
28.1267242431641,-62.9979934692383,
21.0327167510986,-15.0509233474731,
-1.06695652008057,24.0408916473389,
-7.07957410812378,6.53209304809570,
-6.57930898666382,-38.0584907531738,
-19.8549346923828,-40.8977088928223,
-33.7676010131836,9.91748619079590,
-21.3779182434082,53.2239799499512,
9.89770603179932,42.7204666137695,
26.6636657714844,10.7642660140991,
13.6616859436035,10.1299457550049,
-13.4293098449707,33.1516876220703,
-30.4519672393799,33.4401359558106,
-38.8989868164063,4.56939697265625,
-43.1068611145020,-16.4933242797852,
-35.8425674438477,-19.1837158203125,
-17.4409008026123,-30.3004665374756,
-7.11725568771362,-58.7122116088867,
-16.6788558959961,-65.4076919555664,
-30.6922550201416,-30.4759807586670,
-28.5485343933105,1.51777625083923,
-10.2673349380493,-18.4518451690674,
9.06020832061768,-54.4312133789063,
24.3244380950928,-40.6110763549805,
37.8056488037109,14.2001514434814,
41.9952964782715,28.3499240875244,
22.0270557403564,-16.6024723052979,
-18.1731815338135,-41.6372489929199,
-48.3038330078125,1.68006134033203,
-45.4226951599121,46.8158264160156,
-22.8494262695313,14.9209403991699,
-6.24656677246094,-58.0869979858398,
-2.49618291854858,-63.9728507995606,
-1.88991367816925,11.4402132034302,
-4.33550119400024,59.1808929443359,
-5.34094810485840,7.36719608306885,
10.3939647674561,-76.7071533203125,
47.6765899658203,-82.9569854736328,
75.9940643310547,-9.45122337341309,
59.7781448364258,57.1506500244141,
3.88736009597778,65.9454879760742,
-36.0960464477539,43.7065124511719,
-26.7704524993897,28.1755695343018,
0.778298974037170,22.6482620239258,
5.75518178939819,15.8645887374878,
-4.24151802062988,14.9027605056763,
7.19965171813965,24.7554512023926,
27.4738159179688,31.4906826019287,
15.6411218643188,20.1369762420654,
-27.1930046081543,1.50248336791992,
-46.0909004211426,-1.23293304443359,
-10.7015953063965,6.20551824569702,
27.2243156433105,10.3709354400635,
6.34611606597900,15.5756502151489,
-50.3549079895020,26.1266479492188,
-65.4419326782227,26.1261444091797,
-17.9944763183594,6.47367382049561,
34.7346305847168,-19.8192462921143,
36.0049171447754,-25.6590881347656,
4.53474426269531,-0.228121042251587,
-13.5836467742920,28.5268821716309,
-15.6473226547241,39.1129341125488,
-29.1595382690430,31.9411659240723,
-49.5261077880859,13.7359027862549,
-37.3299980163574,-18.5625267028809,
15.1856164932251,-54.4885253906250,
62.2878952026367,-60.6490592956543,
57.4019241333008,-23.8509044647217,
11.9816360473633,14.5703849792480,
-17.7751102447510,5.56777858734131,
-3.25732779502869,-38.3177604675293,
25.4613761901855,-50.3450012207031,
30.0355281829834,-1.22872543334961,
15.6051769256592,58.0995483398438,
9.01795578002930,59.7855987548828,
16.9082756042480,4.53667163848877,
14.0399751663208,-41.7908134460449,
-14.7804918289185,-38.0287857055664,
-37.5635375976563,-8.32968997955322,
-16.9883518218994,8.69233417510986,
28.0052757263184,4.63347291946411,
39.4948463439941,-4.12450504302979,
0.993684053421021,-9.78534412384033,
-35.1126098632813,-17.1302452087402,
-16.1628341674805,-22.8082771301270,
37.1640052795410,-25.3193492889404,
50.7765121459961,-30.9392433166504,
3.19248723983765,-42.7675170898438,
-46.9113349914551,-46.2131538391113,
-42.3022308349609,-24.4757690429688,
-1.60806763172150,9.27936649322510,
15.6004619598389,17.1478118896484,
-10.2255411148071,-11.3236141204834,
-34.2073974609375,-34.7130317687988,
-17.8388919830322,-14.1153469085693,
20.1365356445313,36.4482803344727,
29.7875671386719,69.2492523193359,
-3.49597716331482,56.7208061218262,
-41.9484901428223,18.5287704467773,
-43.9624099731445,-6.53772211074829,
-9.16150188446045,-8.16227531433106,
26.6088180541992,1.40639078617096,
31.9471836090088,7.99119758605957,
10.3854846954346,11.3948125839233,
-9.53137779235840,14.3832015991211,
-5.66864109039307,16.8840961456299,
17.4176902770996,16.8180713653564,
37.7166328430176,12.3233900070190,
31.6886940002441,4.59854507446289,
-1.20709908008575,1.65795063972473,
-35.5496330261231,13.0814533233643,
-42.9825057983398,32.0047111511231,
-20.4623165130615,35.2629241943359,
3.31994533538818,9.12551689147949,
-1.11538386344910,-32.2988739013672,
-24.6286487579346,-59.4192504882813,
-29.9077148437500,-54.9628944396973,
-5.10243177413940,-36.0717124938965,
17.5011081695557,-20.5657691955566,
5.55099010467529,-7.12696456909180,
-32.3570175170898,15.5041389465332,
-52.5359268188477,38.6981773376465,
-34.8834266662598,46.1717262268066,
-4.03800106048584,38.0549316406250,
12.5701799392700,26.3830070495605,
11.6150894165039,18.4789257049561,
0.574141383171082,8.38662815093994,
-17.0659313201904,-5.00644731521606,
-33.3536109924316,-7.59050750732422,
-29.8268585205078,3.68455481529236,
-2.27787399291992,6.87415742874146,
18.4052505493164,-9.72451686859131,
7.50447177886963,-29.0058727264404,
-18.1066608428955,-25.9973888397217,
-14.2189512252808,-10.3606309890747,
20.3011150360107,-18.2733058929443,
39.4471206665039,-50.6136016845703,
12.8413820266724,-61.5533752441406,
-31.7038669586182,-19.3308429718018,
-44.0517692565918,38.1032142639160,
-24.5350055694580,45.7824668884277,
-8.21820259094238,-7.03581666946411,
-11.7026176452637,-58.2253608703613,
-15.0977449417114,-51.9601745605469,
-0.665355086326599,-1.79166293144226,
18.4358921051025,29.0497989654541,
23.5751743316650,9.02692699432373,
22.5017185211182,-26.6860389709473,
34.6645851135254,-33.2234878540039,
58.4189300537109,-7.45876979827881,
68.1754760742188,14.6179885864258,
47.9658317565918,11.5778026580811,
7.94393253326416,1.08868145942688,
-27.8226070404053,8.33064460754395,
-46.3762016296387,21.4910411834717,
-44.9054908752441,12.7133197784424,
-29.1907386779785,-13.4496765136719,
-10.1587619781494,-20.7418384552002,
2.72073984146118,5.02521181106567,
5.60092878341675,32.2442512512207,
3.55707716941834,18.8654479980469,
-0.795868992805481,-28.9710922241211,
-7.62607908248901,-50.8429374694824,
-20.3274745941162,-13.0454921722412,
-32.4269943237305,45.5318717956543,
-27.9883060455322,61.1438598632813,
-4.84131908416748,22.6039104461670,
22.2472858428955,-17.6097335815430,
36.0323410034180,-10.5498437881470,
30.5360355377197,28.5660457611084,
13.4135293960571,47.3966140747070,
0.184419825673103,31.2027072906494,
3.00501728057861,15.6591463088989,
17.1486759185791,24.3696804046631,
20.5788726806641,30.2073745727539,
-1.78181576728821,3.69787526130676,
-38.1060523986816,-36.4540634155273,
-56.1337585449219,-43.5058021545410,
-42.8653602600098,-14.7375364303589,
-27.1759109497070,6.01239013671875,
-42.4316024780273,-7.58398008346558,
-69.5981292724609,-24.6228637695313,
-57.4927062988281,-14.7354087829590,
1.12401986122131,4.96761369705200,
53.4272079467773,1.20347833633423,
59.2138671875000,-19.2324619293213,
42.4528083801270,-18.5788784027100,
46.6997146606445,4.64562940597534,
63.5437927246094,12.0576753616333,
49.4453468322754,-12.6297369003296,
3.23346877098084,-36.0106124877930,
-20.0144634246826,-32.4675559997559,
1.28869283199310,-23.4852809906006,
18.7234325408936,-36.5218200683594,
-9.13897418975830,-59.0362739562988,
-44.7684974670410,-57.1659660339356,
-25.0973129272461,-29.4949932098389,
39.3544921875000,-11.3465166091919,
78.3956146240234,-16.7238368988037,
58.9575462341309,-20.2052288055420,
23.8207664489746,-5.07720184326172,
14.2713775634766,8.86649894714356,
18.8042678833008,0.141331732273102,
12.8266592025757,-17.8087291717529,
8.33778190612793,-22.2569217681885,
33.6240425109863,-14.2119026184082,
64.3173599243164,-7.15719270706177,
54.8472137451172,-1.61297965049744,
10.1847457885742,10.4227085113525,
-15.2469406127930,24.7305679321289,
6.70295286178589,20.5711059570313,
41.0938987731934,1.64979338645935,
47.5133895874023,-6.46006965637207,
26.6939735412598,7.44029235839844,
2.65574145317078,18.3583354949951,
-12.4900236129761,4.22773838043213,
-24.3693275451660,-23.7685718536377,
-33.0300865173340,-39.3591651916504,
-26.9795417785645,-39.7714996337891,
-19.7727050781250,-37.4522399902344,
-28.0507717132568,-31.0049133300781,
-43.7460937500000,-10.3430337905884,
-39.5312843322754,17.6400470733643,
-12.4513120651245,23.7103309631348,
10.0196056365967,-5.98809576034546,
17.5540904998779,-42.9702453613281,
29.2287712097168,-50.2652893066406,
45.8715095520020,-22.6702804565430,
41.0084228515625,12.0782299041748,
-0.157569766044617,30.9946460723877,
-40.1215209960938,27.2104282379150,
-27.0750579833984,6.70612335205078,
28.2779312133789,-11.1244258880615,
56.1384811401367,-1.76213598251343,
19.7134552001953,36.9724006652832,
-42.9120407104492,67.4673385620117,
-71.3568496704102,51.1471405029297,
-53.9426765441895,-4.70638561248779,
-13.0001382827759,-42.6794281005859,
28.5180320739746,-27.6586456298828,
53.1153793334961,11.2251424789429,
40.6057052612305,24.7277088165283,
-6.90131139755249,10.6120891571045,
-50.3441238403320,7.53778457641602,
-47.7708816528320,21.2800960540772,
-13.7110252380371,24.6584129333496,
-2.81524515151978,2.77674937248230,
-33.6251983642578,-19.0822811126709,
-58.5359039306641,-19.1155700683594,
-42.0426521301270,-14.0032453536987,
-15.8076286315918,-28.0582313537598,
-17.6145973205566,-51.0735473632813,
-25.5756931304932,-50.7539482116699,
-4.92454338073731,-27.6044158935547,
25.7080669403076,-10.4117116928101,
20.3677253723145,-11.7922735214233,
-22.2310562133789,-12.0776176452637,
-38.4806747436523,-6.42376232147217,
-4.47683238983154,-16.1192302703857,
22.5966129302979,-41.9804916381836,
2.35876893997192,-52.9577064514160,
-25.5138854980469,-34.4144821166992,
-3.04116296768188,-16.8726615905762,
40.2260437011719,-27.5959892272949,
35.2052459716797,-42.4993934631348,
-12.6367864608765,-15.5672645568848,
-26.1357288360596,40.4750747680664,
15.1266231536865,58.7601776123047,
42.6920890808106,20.6363468170166,
5.28940534591675,-19.9555263519287,
-43.0010986328125,-14.0065240859985,
-22.5822963714600,12.2242250442505,
47.1922111511231,10.8596105575562,
72.5447387695313,-11.8923511505127,
18.9977436065674,-12.7966365814209,
-44.6620407104492,9.60948085784912,
-53.2853660583496,15.4010887145996,
-24.8043804168701,-6.83788919448853,
-10.7976970672607,-14.9698228836060,
-16.8432865142822,19.8732528686523,
-19.6531276702881,53.8646354675293,
-12.6708202362061,30.7454528808594,
-9.91144084930420,-38.0982856750488,
-13.7517929077148,-78.5366058349609,
-7.34281063079834,-50.5064315795898,
14.7336988449097,7.29073143005371,
29.2322387695313,34.0922164916992,
20.1403827667236,11.7124137878418,
0.474465608596802,-25.6734523773193,
-11.5444135665894,-35.8161239624023,
-15.8676700592041,-12.8228626251221,
-17.5950622558594,18.8384742736816,
-15.7211284637451,29.7175045013428,
-16.0421714782715,10.5685577392578,
-26.0112705230713,-24.3070316314697,
-39.5909309387207,-52.9476509094238,
-37.0864601135254,-59.5808219909668,
-12.5977325439453,-48.1773872375488,
10.2571220397949,-29.6392650604248,
3.32698583602905,-10.7022628784180,
-28.6777877807617,4.45624971389771,
-48.9001693725586,10.2221651077271,
-35.1131057739258,4.77898216247559,
-7.45074796676636,-14.4470615386963,
4.46906280517578,-38.4500122070313,
-0.232222884893417,-50.7895812988281,
-8.99589729309082,-38.6583557128906,
-11.4950113296509,-8.09834861755371,
-7.10952425003052,16.4406433105469,
0.889460623264313,11.6271638870239,
4.80709981918335,-14.7157669067383,
-5.81341791152954,-36.7226600646973,
-30.5001678466797,-39.7512893676758,
-40.5129203796387,-31.4563846588135,
-8.14430236816406,-26.1909503936768,
42.0599555969238,-21.0939483642578,
53.5576438903809,-9.32108402252197,
8.42240810394287,0.982003569602966,
-35.9814338684082,-8.20924186706543,
-17.1281986236572,-30.1906070709229,
44.4301834106445,-38.4628906250000,
76.0295028686523,-21.2197113037109,
47.1060180664063,1.62545275688171,
6.35052394866943,3.76145935058594,
3.74101567268372,-8.25278949737549,
18.7302093505859,-0.423681646585465,
-0.749269723892212,32.6433601379395,
-50.1431884765625,56.6081886291504,
-72.3290023803711,35.2189979553223,
-36.6609535217285,-17.1551361083984,
19.2135715484619,-52.1921615600586,
41.0736999511719,-41.2030830383301,
24.8466529846191,-14.8711042404175,
6.08353233337402,-18.0050392150879,
-0.806093573570252,-46.8376235961914,
-4.29939413070679,-55.2110023498535,
-15.4642267227173,-15.2623243331909,
-24.6721611022949,42.8035812377930,
-16.7679271697998,63.8389472961426,
5.19778490066528,32.1679344177246,
20.5961837768555,-8.37135696411133,
22.9180107116699,-12.6199026107788,
22.0312690734863,15.3469343185425,
26.0686893463135,40.1494255065918,
32.4652900695801,42.6288757324219,
27.9391250610352,39.9259300231934,
1.52872550487518,47.2726097106934,
-31.6693801879883,53.5529785156250,
-31.2038764953613,32.4188385009766,
14.7639646530151,-11.5521497726440,
66.9049301147461,-36.8243446350098,
74.4660644531250,-20.5639362335205,
30.8828639984131,15.2748594284058,
-6.63346576690674,27.8233261108398,
1.44484424591064,2.48111891746521,
21.8808002471924,-22.1875476837158,
-3.32466340065002,-6.92026138305664,
-60.7847366333008,31.2186164855957,
-75.5498352050781,44.8690795898438,
-17.8366489410400,13.7436666488647,
43.7311325073242,-31.3697586059570,
35.9639244079590,-48.8408164978027,
-17.7809734344482,-34.3703422546387,
-31.4147224426270,-21.5504798889160,
15.7346544265747,-19.8539867401123,
48.5241889953613,-3.21283698081970,
5.37099266052246,39.9375762939453,
-72.7072067260742,67.1507644653320,
-102.519279479980,36.1003456115723,
-61.9150009155273,-31.7559452056885,
-9.80652999877930,-60.4389228820801,
6.17068719863892,-19.1806049346924,
-5.20919036865234,34.2807655334473,
-21.7227497100830,31.2676963806152,
-37.8651657104492,-12.2918357849121,
-48.1096115112305,-27.3211193084717,
-37.5772895812988,3.57748150825501,
-4.64929914474487,25.2637176513672,
33.6156387329102,-3.21606683731079,
53.5904312133789,-40.9650154113770,
49.5017776489258,-29.0168037414551,
33.6884040832520,18.5657634735107,
11.9780645370483,38.6639671325684,
-8.00456905364990,9.43517112731934,
-2.28773212432861,-27.5198917388916,
27.8298454284668,-34.8232536315918,
35.2182083129883,-23.6039676666260,
-9.91080474853516,-21.1948127746582,
-58.7135772705078,-26.9727878570557,
-41.6973991394043,-22.5689144134522,
27.4504451751709,-10.8622751235962,
55.9571762084961,-4.12931299209595,
3.80351781845093,4.57583141326904,
-52.9024543762207,18.4268741607666,
-31.6686096191406,21.0300102233887,
38.0453605651856,-3.92802071571350,
56.8282012939453,-37.6896171569824,
11.3860883712769,-48.4184989929199,
-12.1281747817993,-34.6836090087891,
27.3893127441406,-21.8019351959229,
66.5347290039063,-19.0129299163818,
42.9487838745117,-1.93532657623291,
-7.74932765960693,38.0966186523438,
-16.5063533782959,64.0520248413086,
14.9352121353149,39.9423675537109,
32.0324058532715,-6.61264419555664,
21.7031803131104,-17.6411628723145,
18.6532878875732,20.4134578704834,
31.2842121124268,62.5249099731445,
17.6548385620117,65.5738296508789,
-32.3630065917969,39.7742042541504,
-58.2763633728027,22.4435367584229,
-22.7455921173096,23.8303833007813,
25.1042633056641,27.3257637023926,
31.3276443481445,21.2830924987793,
15.3112325668335,12.8915548324585,
20.0556812286377,16.1940116882324,
34.3643035888672,23.6601448059082,
14.1455459594727,26.0250988006592,
-29.2092304229736,25.4898395538330,
-36.2146072387695,30.6855068206787,
1.31291675567627,38.6777610778809,
19.3824424743652,36.5404624938965,
-17.9826297760010,17.1524124145508,
-48.3456802368164,-9.75354290008545,
-14.5217800140381,-16.7183380126953,
41.1838989257813,6.52309417724609,
35.0868568420410,32.9986572265625,
-25.1558284759522,26.9888820648193,
-58.9296264648438,-18.8872699737549,
-35.7168426513672,-62.8071708679199,
-9.85489463806152,-58.4767684936523,
-26.7133274078369,-8.71475791931152,
-53.5102005004883,31.1836795806885,
-35.2105178833008,22.4976272583008,
14.9022016525269,-12.7390699386597,
44.5882720947266,-19.5070438385010,
41.9635848999023,13.3058729171753,
42.1316528320313,40.7600860595703,
54.9307518005371,23.9082088470459,
52.6937713623047,-20.2353000640869,
28.8395271301270,-41.6962318420410,
16.7934951782227,-22.6226329803467,
33.8732185363770,6.30901861190796,
51.9814300537109,11.7915372848511,
40.4330749511719,1.19766640663147,
11.9065504074097,-0.861852109432221,
4.71619749069214,16.3546199798584,
25.9253978729248,37.7118415832520,
39.2111396789551,42.0242958068848,
23.8477134704590,24.6573009490967,
-3.37515211105347,-5.68879604339600,
-14.7341756820679,-28.5413169860840,
-13.0399322509766,-22.2022895812988,
-17.4371471405029,11.7793560028076,
-30.3074188232422,41.7731208801270,
-36.8327827453613,37.5214691162109,
-25.9701213836670,5.70434427261353,
-6.66105365753174,-10.6769733428955,
4.33973789215088,13.9335203170776,
2.91982507705688,52.9237060546875,
1.25499975681305,61.0502586364746,
5.62814235687256,30.9778804779053,
2.77219176292419,0.346735954284668,
-17.1560516357422,-1.71208477020264,
-40.7569046020508,14.8239154815674,
-42.3028335571289,18.6561012268066,
-17.1247444152832,-0.203350663185120,
8.91099262237549,-20.3926410675049,
5.50863552093506,-22.1816635131836,
-17.6716632843018,-7.47312116622925,
-26.8940181732178,10.8118495941162,
-10.8817758560181,21.6474761962891,
3.96493816375732,26.7049236297607,
-9.50058078765869,28.4872074127197,
-39.2563247680664,27.3181438446045,
-49.4565582275391,22.8450870513916,
-28.9354171752930,5.51096248626709,
-4.73639488220215,-24.2771816253662,
-5.74209070205689,-47.8208770751953,
-24.9404773712158,-49.8082733154297,
-29.4097080230713,-31.1276779174805,
-4.61481332778931,-11.4511241912842,
25.6959800720215,-7.62132215499878,
31.6837692260742,-10.4763059616089,
9.75309085845947,-3.42939901351929,
-14.1303548812866,11.2173070907593,
-18.2539215087891,21.5544414520264,
-7.36597537994385,29.6686801910400,
0.846608877182007,42.1160545349121,
-3.23057389259338,42.9300384521484,
-15.7282686233521,9.69571304321289,
-26.9317111968994,-45.4721069335938,
-27.8373146057129,-67.6324691772461,
-15.5656719207764,-26.6480941772461,
3.12406492233276,32.1338996887207,
8.53290653228760,37.7689933776856,
-3.80157470703125,-13.8593502044678,
-15.6827917098999,-59.0123481750488,
-10.3482856750488,-48.4269905090332,
0.648303210735321,-13.6978559494019,
-9.60282707214356,-7.28074550628662,
-39.7055282592773,-28.3270988464355,
-55.7176055908203,-36.5704536437988,
-35.3943862915039,-20.6776027679443,
-6.75970268249512,-10.5026569366455,
-6.68387794494629,-24.8940181732178,
-23.1438350677490,-42.5641250610352,
-16.8950405120850,-36.2486038208008,
12.6986227035522,-13.4065246582031,
18.7678623199463,3.53399848937988,
-18.1941490173340,5.55360412597656,
-51.9882431030273,1.83027112483978,
-31.7890205383301,-8.22370243072510,
22.6931438446045,-29.1711883544922,
48.4805984497070,-40.7377433776856,
27.4533920288086,-22.2695426940918,
3.60509634017944,9.65112495422363,
11.4380779266357,20.6003284454346,
26.1656894683838,-2.89438295364380,
7.31867074966431,-37.6030540466309,
-33.5315132141113,-54.9429130554199,
-47.9984588623047,-44.7862663269043,
-20.1546802520752,-18.7928180694580,
17.2929286956787,11.0242309570313,
29.1209049224854,23.9084014892578,
15.4626255035400,-3.46123695373535,
-0.285625457763672,-56.9885520935059,
-1.70739567279816,-73.1010589599609,
4.91227245330811,-22.1770992279053,
4.12923288345337,42.0482215881348,
-5.52849960327148,44.8138008117676,
-15.4086608886719,-7.11313438415527,
-10.2283391952515,-34.4893302917481,
18.4111194610596,-4.48134708404541,
45.6375083923340,25.4026489257813,
40.7792549133301,0.570818662643433,
0.715303897857666,-39.7143058776856,
-40.8303871154785,-24.3476676940918,
-54.5403900146484,30.3478755950928,
-45.2662277221680,38.3262939453125,
-33.6461486816406,-17.2496528625488,
-23.4667339324951,-55.2236022949219,
-1.63820397853851,-13.6727371215820,
25.5874500274658,56.2309799194336,
26.4514980316162,65.4720153808594,
-8.54080677032471,15.0249862670898,
-43.4970626831055,-20.8109035491943,
-31.2869262695313,-6.73601341247559,
23.8160476684570,15.9383287429810,
68.2642211914063,4.34456825256348,
64.7970046997070,-22.2640438079834,
30.3839149475098,-19.9941577911377,
6.30658435821533,6.09814405441284,
6.13466072082520,16.1672325134277,
9.90682888031006,-1.52807092666626,
-4.31046915054321,-20.6801128387451,
-27.4358177185059,-19.1995334625244,
-35.3344345092773,-5.63275432586670,
-19.9772090911865,4.41698455810547,
2.49476289749146,1.24379801750183,
5.27962875366211,-12.8960094451904,
-16.1598873138428,-30.7586631774902,
-38.9736862182617,-46.2594299316406,
-36.5294609069824,-54.1940383911133,
-3.54137825965881,-48.7039031982422,
30.4582633972168,-37.0633964538574,
30.5804767608643,-27.2311458587647,
-2.28041338920593,-17.7639579772949,
-30.8726978302002,-7.79243230819702,
-18.0695056915283,4.53690481185913,
30.1319599151611,21.9137744903564,
65.9191207885742,41.8701477050781,
47.7083702087402,48.6836357116699,
-9.09412860870361,26.5945835113525,
-47.1045455932617,-14.5951786041260,
-29.1109199523926,-42.9018478393555,
16.3805236816406,-33.2275886535645,
28.4161682128906,-4.05120992660523,
-6.68053865432739,6.35298490524292,
-39.0345573425293,-14.1569032669067,
-19.8835601806641,-33.3263549804688,
31.2217960357666,-18.0744342803955,
47.9143257141113,25.0490226745605,
3.94440126419067,54.2430648803711,
-53.0556106567383,47.7660255432129,
-63.1013374328613,23.6866397857666,
-23.6342449188232,8.86727428436279,
21.5114154815674,5.31806993484497,
39.0499420166016,-3.47272706031799,
37.8740043640137,-25.1560287475586,
42.0533866882324,-39.9057731628418,
48.0852050781250,-27.9030094146729,
45.6930847167969,7.99507427215576,
35.8700218200684,41.9031982421875,
28.4872303009033,49.5646095275879,
24.1487789154053,31.9463500976563,
9.63884353637695,9.80842018127441,
-18.1855964660645,4.35553121566773,
-43.9401321411133,16.2960243225098,
-46.1424522399902,27.6534519195557,
-29.2093467712402,19.0978126525879,
-13.7868041992188,2.32084417343140,
-14.8925590515137,-0.368579089641571,
-25.1570301055908,20.5596733093262,
-16.2179622650147,39.0959701538086,
18.7511425018311,29.1108303070068,
55.3790473937988,-1.87201249599457,
60.5218467712402,-16.0447521209717,
23.3127155303955,7.35461282730103,
-27.0572204589844,42.5499496459961,
-49.3956451416016,50.6101074218750,
-26.8625259399414,20.5423851013184,
16.7115840911865,-14.8246164321899,
46.7188568115234,-18.0865859985352,
50.0964202880859,8.52678108215332,
39.6193466186523,36.5122108459473,
32.1625747680664,46.6998443603516,
23.9242534637451,43.4797019958496,
-1.92846608161926,41.8645095825195,
-38.0975074768066,42.5505790710449,
-54.7320060729981,36.3282775878906,
-33.1146697998047,25.2206153869629,
5.10203027725220,20.0532932281494,
16.5555953979492,13.2676048278809,
-8.26626205444336,-11.5593328475952,
-33.9819221496582,-47.0429306030273,
-21.8817653656006,-58.7899017333984,
16.8958950042725,-29.9038467407227,
42.3837623596191,8.03056049346924,
43.2882499694824,10.3447446823120,
42.9211769104004,-13.1887664794922,
52.5056877136231,-11.9548931121826,
45.7779083251953,26.7881031036377,
3.97613096237183,52.8872337341309,
-43.4463119506836,25.7520656585693,
-52.0418968200684,-22.0006103515625,
-13.9931182861328,-26.1267127990723,
29.8810291290283,12.1556873321533,
43.9220199584961,31.4142074584961,
32.3492012023926,3.76398515701294,
14.5650806427002,-29.6120586395264,
-3.18992543220520,-20.0295867919922,
-15.8935852050781,15.2539043426514,
-12.4328880310059,28.0259571075439,
1.05361139774323,9.99255943298340,
-0.917717814445496,-3.80781984329224,
-20.9764080047607,6.91590404510498,
-20.5388736724854,21.8371582031250,
19.5603218078613,16.2089633941650,
58.4839859008789,0.559278666973114,
37.6556243896484,-9.14733791351318,
-25.1929893493652,-15.4275169372559,
-47.8536911010742,-25.6434898376465,
6.82542610168457,-29.7998580932617,
67.5742797851563,-16.2309265136719,
56.9511146545410,10.2926979064941,
-4.61949110031128,30.2532711029053,
-33.1500205993652,35.0689392089844,
-1.94215893745422,34.8802909851074,
34.9047698974609,39.5533447265625,
29.1792392730713,42.3772392272949,
-4.71354103088379,36.2006072998047,
-29.7356605529785,19.3830947875977,
-39.5048065185547,-7.89070367813110,
-45.2367477416992,-43.3592987060547,
-35.7236785888672,-71.2996215820313,
-2.52876853942871,-68.8777465820313,
26.7582817077637,-30.6580505371094,
15.6771373748779,15.3381347656250,
-28.1021556854248,31.1029453277588,
-55.1799278259277,10.4668645858765,
-46.3578567504883,-17.2628402709961,
-39.1508026123047,-22.2553710937500,
-50.1243171691895,-6.31324386596680,
-52.1927909851074,0.0545630753040314,
-17.1235275268555,-18.3124961853027,
29.9705123901367,-42.4867477416992,
33.5521469116211,-45.1926155090332,
-11.8727664947510,-29.3828372955322,
-44.5378646850586,-21.8692512512207,
-19.9996299743652,-38.4437522888184,
34.7836265563965,-53.3191795349121,
58.9864997863770,-35.2306594848633,
29.3176689147949,4.65558958053589,
-17.8209304809570,24.2543277740479,
-33.9211730957031,-0.608369827270508,
-7.48651361465454,-35.8285293579102,
38.5419502258301,-33.2327194213867,
70.3060989379883,5.74748420715332,
64.8355255126953,36.6642150878906,
26.9367179870605,22.8919601440430,
-15.9539422988892,-17.5472850799561,
-34.4434204101563,-41.0506973266602,
-12.0598907470703,-25.5270061492920,
30.9562644958496,7.89172315597534,
51.8337364196777,29.8766651153564,
29.4542751312256,27.2469177246094,
-17.5916366577148,15.2061996459961,
-52.7102165222168,13.1429080963135,
-55.2232704162598,26.2073707580566,
-42.0837326049805,36.6086311340332,
-43.3401565551758,26.6730155944824,
-50.2096328735352,-6.63999986648560,
-32.1546630859375,-41.8574066162109,
17.9577789306641,-54.1235809326172,
61.2445030212402,-40.6614990234375,
50.1992721557617,-24.4909744262695,
-10.8297176361084,-21.5750293731689,
-56.0889434814453,-32.3319816589356,
-38.9908638000488,-45.3379402160645,
15.9008541107178,-47.3802337646484,
40.5412521362305,-35.7684440612793,
5.91931343078613,-15.3347549438477,
-38.1355056762695,2.54854536056519,
-30.0457763671875,-0.367597162723541,
28.6280460357666,-23.8872966766357,
73.3797302246094,-47.0806427001953,
56.3311767578125,-46.2569427490234,
2.39247608184814,-25.1399574279785,
-27.9594631195068,-3.98819518089294,
-12.5895576477051,6.90130853652954,
10.9881200790405,20.8031711578369,
2.33184719085693,43.5445938110352,
-34.5545463562012,51.7027702331543,
-57.4823837280273,22.9044551849365,
-36.5142707824707,-23.3797264099121,
13.2323036193848,-37.9356155395508,
51.5726890563965,-1.89998292922974,
48.7646942138672,46.9616928100586,
14.9505949020386,61.0274276733398,
-8.59724330902100,35.6569061279297,
1.86225640773773,9.59572505950928,
27.5276069641113,6.32217884063721,
31.8313903808594,7.53412628173828,
2.60814380645752,-9.42602825164795,
-31.1495265960693,-31.2399787902832,
-35.7600402832031,-30.6175270080566,
-18.1114234924316,-4.80896282196045,
-7.49930810928345,11.4588479995728,
-4.37043094635010,-7.95814418792725,
9.05684757232666,-39.6933937072754,
30.7633800506592,-40.0670967102051,
33.3128662109375,-0.623198032379150,
10.8036489486694,38.5837211608887,
-5.93050003051758,35.4656639099121,
8.86746215820313,-2.72638893127441,
30.9526157379150,-28.8992080688477,
18.8658943176270,-11.3976640701294,
-20.8176422119141,20.6943035125732,
-41.5805740356445,20.1555480957031,
-29.3854370117188,-12.0416908264160,
-21.4802227020264,-25.0817623138428,
-37.6262855529785,11.3154830932617,
-44.2241058349609,58.4457359313965,
-8.34071063995361,56.9764671325684,
38.2407035827637,0.110062599182129,
45.9707946777344,-43.0819396972656,
19.1112270355225,-21.9569396972656,
5.48964500427246,30.4365520477295,
18.6559696197510,52.4050407409668,
13.6574859619141,40.8782997131348,
-32.9657707214356,35.1317672729492,
-71.7580108642578,42.4218788146973,
-51.1763076782227,24.9996032714844,
3.45241546630859,-21.9855499267578,
18.5212821960449,-47.5036659240723,
-23.1724681854248,-19.8094139099121,
-65.9851989746094,10.6224222183228,
-60.7970809936523,-14.6364860534668,
-15.6908969879150,-61.2730102539063,
28.8567008972168,-46.9241714477539,
51.9041900634766,28.0553436279297,
47.5656509399414,70.5205612182617,
15.8827695846558,30.2088718414307,
-29.7638931274414,-24.2320995330811,
-54.9627342224121,-21.0966529846191,
-30.6536102294922,12.5925521850586,
20.9050655364990,7.56746101379395,
49.8095626831055,-25.6141929626465,
42.9260711669922,-15.4750595092773,
27.6390647888184,44.4780807495117,
19.6909980773926,76.4438552856445,
14.1702127456665,37.2818222045898,
2.09373807907105,-19.9444255828857,
-10.3575735092163,-27.5000286102295,
-17.0298557281494,-5.35797119140625,
-20.7657012939453,-4.96447801589966,
-27.8305130004883,-20.3431072235107,
-25.3528308868408,-6.63507080078125,
-11.2911243438721,24.6575298309326,
-10.3088331222534,17.1226558685303,
-32.9493980407715,-39.7474098205566,
-46.5933074951172,-83.7284851074219,
-13.2425994873047,-61.5597381591797,
46.4086837768555,-2.60143518447876,
61.0516777038574,24.3827819824219,
7.48897457122803,0.668257772922516,
-53.5919342041016,-33.3439598083496,
-56.2399559020996,-45.4994621276856,
-12.7949409484863,-45.7744522094727,
8.89155292510986,-45.6726799011231,
-19.2005443572998,-43.3828659057617,
-54.7710418701172,-35.5182838439941,
-48.5283203125000,-23.7228126525879,
-13.1928024291992,-11.1412181854248,
9.69187259674072,4.76792669296265,
4.37389230728149,23.3268985748291,
-2.88400053977966,36.4437179565430,
7.45086145401001,36.5854148864746,
28.8495521545410,24.0751056671143,
37.9655227661133,7.08056640625000,
26.3415470123291,-11.8485393524170,
-0.659428477287293,-25.6975536346436,
-23.4677085876465,-14.5984563827515,
-28.1455516815186,19.8153686523438,
-18.0544776916504,43.0814666748047,
-9.80790042877197,25.8435688018799,
-20.5022506713867,-17.0081233978272,
-45.8208427429199,-35.3923225402832,
-61.9032287597656,-16.3204212188721,
-56.5085487365723,8.20960617065430,
-46.5038719177246,6.57217979431152,
-48.7188644409180,-4.90760135650635,
-60.4588088989258,3.04881739616394,
-62.9360771179199,21.3932456970215,
-44.9320602416992,10.1207838058472,
-12.4905185699463,-34.4310646057129,
20.6141567230225,-62.9793205261231,
44.4963798522949,-41.5551757812500,
52.1245574951172,5.97309017181397,
39.4583206176758,33.8622817993164,
18.4092445373535,26.6245651245117,
12.2209596633911,-0.459830611944199,
24.8623828887939,-31.6676025390625,
32.2062339782715,-53.1904487609863,
16.1002655029297,-49.4407691955566,
-11.8553638458252,-19.7992210388184,
-20.5090065002441,5.30206394195557,
-5.19031620025635,-12.2674942016602,
10.6148376464844,-53.0816116333008,
10.6909685134888,-54.1578445434570,
12.3123130798340,0.357310175895691,
29.4483070373535,50.7538604736328,
46.9026603698731,48.9360046386719,
35.6798515319824,19.3626594543457,
5.11862277984619,13.0578422546387,
-4.19032526016235,22.7706317901611,
22.1606502532959,10.1035985946655,
45.9966354370117,-21.5233402252197,
24.0885467529297,-22.7970695495605,
-30.3616695404053,12.4087114334106,
-60.9593811035156,20.0099906921387,
-36.6732254028320,-27.3705501556397,
14.7740631103516,-67.4412307739258,
42.5808067321777,-38.4852714538574,
27.4120521545410,19.3930950164795,
-0.372425079345703,21.9567890167236,
-10.7809247970581,-27.9902667999268,
-1.18213796615601,-43.5031700134277,
7.18109989166260,10.5018386840820,
0.372767329216003,67.3549423217773,
-12.9710874557495,61.8598785400391,
-13.4563474655151,20.3034210205078,
7.93140554428101,11.8135986328125,
30.9026603698730,32.2996215820313,
32.7200584411621,24.8331661224365,
18.2534599304199,-21.3571681976318,
7.58165502548218,-47.0581054687500,
5.12635087966919,-15.1632146835327,
-5.77069711685181,31.2528457641602,
-38.2955818176270,38.3548851013184,
-70.8490142822266,13.8645763397217,
-71.2031860351563,-0.948237836360931,
-48.1733627319336,9.24217033386231,
-37.5178680419922,22.6901397705078,
-41.0282325744629,20.4191493988037,
-26.8946056365967,14.5255022048950,
15.8016490936279,21.1721897125244,
43.5581283569336,25.6406497955322,
21.2435855865479,8.33286094665527,
-17.6217422485352,-22.3850784301758,
-9.98563575744629,-42.4681282043457,
40.8813705444336,-34.9597434997559,
61.4231338500977,-2.87253618240356,
19.6593074798584,31.1455116271973,
-25.7227973937988,31.9331684112549,
-8.04961013793945,-4.30972051620483,
44.9907798767090,-34.9914207458496,
47.4821929931641,-17.8353652954102,
-19.0532913208008,35.8272552490234,
-80.4642715454102,61.4473037719727,
-81.5359268188477,18.4784355163574,
-43.8658561706543,-47.2216873168945,
-20.5874710083008,-56.8538246154785,
-19.0036354064941,-5.38282203674316,
-11.0279493331909,40.9916076660156,
8.11529254913330,43.7299957275391,
13.0697193145752,35.7428550720215,
-8.37953090667725,43.4886512756348,
-33.8352584838867,34.8649978637695,
-41.8112907409668,-18.2297935485840,
-30.8103733062744,-72.2642822265625,
-2.15281462669373,-55.9224586486816,
37.9898300170898,14.9312400817871,
58.5026664733887,44.9486351013184,
27.9799270629883,-1.74444007873535,
-27.9925289154053,-50.4949989318848,
-46.6814880371094,-31.5389003753662,
-6.05301761627197,19.9287204742432,
45.8390579223633,23.1759262084961,
44.5540733337402,-15.1584434509277,
7.16270399093628,-23.2296504974365,
-2.23556923866272,11.3099937438965,
31.7175731658936,33.0532341003418,
56.4046211242676,13.5792579650879,
39.0657844543457,-2.69086480140686,
10.2565469741821,24.0936908721924,
10.0881872177124,50.8705558776856,
24.9235553741455,23.4954910278320,
25.5283412933350,-32.4747314453125,
14.4580717086792,-44.4807167053223,
18.1908569335938,2.24232625961304,
26.3445529937744,46.3647918701172,
3.58867788314819,50.4440956115723,
-48.4926033020020,37.4802970886231,
-78.4180297851563,27.4637050628662,
-51.3263893127441,7.03112792968750,
-1.95269012451172,-31.9963703155518,
12.9330949783325,-59.0209236145020,
-9.17644882202148,-44.1464462280273,
-23.9033737182617,-5.31049013137817,
-6.39794921875000,8.95857810974121,
24.5285243988037,-10.6680269241333,
43.6899795532227,-26.3961219787598,
48.1972351074219,-16.8429737091064,
49.9014701843262,2.71615862846375,
47.3125190734863,14.2661352157593,
31.4016666412354,19.8867549896240,
4.90767288208008,15.2903089523315,
-12.4936122894287,-9.83297157287598,
-11.1500520706177,-38.9212303161621,
1.11650395393372,-39.0456848144531,
7.00723123550415,-6.76694583892822,
-0.877310156822205,12.0202121734619,
-18.5186920166016,-18.0486927032471,
-33.0518341064453,-61.9893264770508,
-33.8989257812500,-58.2250900268555,
-23.9701251983643,-3.08156585693359,
-12.5238656997681,38.8771171569824,
-5.88508272171021,25.4479541778564,
-3.23380351066589,-10.4717683792114,
-1.05429315567017,-20.8516731262207,
1.43781745433807,-8.18266487121582,
-1.46218442916870,-2.60492229461670,
-9.81790828704834,-8.12282848358154,
-22.3482913970947,-0.738293707370758,
-30.6474494934082,22.1197052001953,
-26.0935192108154,28.7642135620117,
-5.85538196563721,1.24771881103516,
20.6075973510742,-36.2488937377930,
40.8793067932129,-47.1893310546875,
45.4378356933594,-27.6796474456787,
37.1389694213867,1.06329345703125,
25.3131332397461,24.8142375946045,
15.7751884460449,41.2285537719727,
10.6925230026245,41.4195976257324,
16.2252635955811,22.5951557159424,
28.2789306640625,1.93272900581360,
30.4366111755371,-0.524560868740082,
10.2477169036865,13.8940925598145,
-19.1833610534668,20.8969020843506,
-27.5013370513916,8.52542781829834,
-0.890081882476807,-5.39847469329834,
28.0345230102539,-0.285632848739624,
17.5023975372314,15.0574836730957,
-30.7179718017578,16.8300304412842,
-64.3438796997070,3.81642460823059,
-40.8192520141602,-3.40236282348633,
17.0213851928711,4.12516975402832,
42.9155921936035,15.3368768692017,
10.8569192886353,13.6439495086670,
-33.2576255798340,5.33854341506958,
-30.3616371154785,5.62393474578857,
7.30924987792969,15.8542633056641,
16.9359130859375,27.1051807403564,
-26.9677467346191,28.6604385375977,
-69.4574584960938,21.2659244537354,
-47.4552764892578,9.04252243041992,
22.0671806335449,-6.82935714721680,
66.2981948852539,-18.6319942474365,
47.1016578674316,-17.9546775817871,
2.60697960853577,-2.92431974411011,
-15.5945329666138,12.8715610504150,
-8.02854347229004,11.8038396835327,
-7.58265876770020,-8.76726055145264,
-19.6713981628418,-36.2725830078125,
-18.4214515686035,-49.8600196838379,
8.18450832366943,-38.8072357177734,
35.4285507202148,-8.48566913604736,
38.8233070373535,21.3118991851807,
16.7237949371338,29.9871654510498,
-15.7957725524902,13.2125253677368,
-34.3159103393555,-12.8567104339600,
-19.7257366180420,-18.5927238464355,
21.4846668243408,5.90898990631104,
52.8893737792969,46.3159523010254,
40.6867523193359,68.7360229492188,
-4.45600080490112,53.8213729858398,
-24.9303112030029,15.5491056442261,
10.1586999893188,-17.6053009033203,
54.9087181091309,-28.8540229797363,
54.6531715393066,-25.5759506225586,
24.1336059570313,-22.2721004486084,
16.5687675476074,-23.6144561767578,
34.8967208862305,-23.3450889587402,
31.2765731811523,-13.4199466705322,
-9.86145782470703,4.17491006851196,
-37.3416862487793,29.4794120788574,
-10.8201017379761,54.0582008361816,
29.0620918273926,58.3971099853516,
22.2826213836670,28.7588863372803,
-15.8435544967651,-16.0989532470703,
-18.8520298004150,-36.3137893676758,
21.8262901306152,-13.2771596908569,
43.0845718383789,22.3947067260742,
12.4686613082886,27.0007495880127,
-19.9855327606201,3.28804063796997,
-6.67524909973145,-8.30993652343750,
23.4563293457031,12.9813184738159,
17.9445571899414,35.7665405273438,
-16.8427200317383,19.3536911010742,
-31.8224449157715,-28.3806819915772,
-15.5024223327637,-58.9510078430176,
-2.89363718032837,-52.3438186645508,
-8.47009277343750,-33.2368125915527,
-0.894273996353149,-29.4001407623291,
35.0816383361816,-34.5963439941406,
60.0508003234863,-19.2370052337647,
46.6575088500977,19.2688674926758,
26.2092437744141,54.0557975769043,
32.6424674987793,61.0218048095703,
45.4751129150391,42.5999565124512,
28.8267784118652,20.2481937408447,
-5.25609827041626,11.1375646591187,
-9.32975959777832,12.4493722915649,
20.1705760955811,11.2997703552246,
36.3629837036133,-2.92132091522217,
15.5667209625244,-29.1767482757568,
-8.23407649993897,-46.8903923034668,
-1.91741085052490,-34.9408035278320,
7.58480930328369,0.597443580627441,
-13.6634187698364,33.3293418884277,
-41.0336837768555,33.1094245910645,
-32.4195747375488,0.0314354896545410,
2.34095382690430,-36.5403518676758,
9.17470169067383,-48.4741859436035,
-21.5910205841064,-36.8265419006348,
-38.9740295410156,-25.5854511260986,
-2.38622093200684,-32.6754379272461,
55.1584663391113,-47.8433532714844,
77.0620040893555,-40.9663810729981,
51.1497573852539,-5.46344041824341,
14.7739562988281,31.8590507507324,
-11.0808019638062,36.3032989501953,
-32.0435638427734,4.53433895111084,
-44.1345367431641,-35.4497451782227,
-22.0438137054443,-50.5157432556152,
30.3022460937500,-32.4109954833984,
71.6712493896484,5.81808757781982,
65.8564376831055,41.5702590942383,
27.8017425537109,47.6489601135254,
-4.72381162643433,16.8430061340332,
-8.17292976379395,-26.5781764984131,
3.50018835067749,-42.0250167846680,
7.70644617080689,-16.7852382659912,
-0.404138445854187,13.9459838867188,
-15.3627634048462,16.1154708862305,
-31.0902481079102,-2.39164566993713,
-38.8015632629395,-10.7692728042603,
-32.4815483093262,-2.55011534690857,
-25.5454959869385,-1.90130114555359,
-28.6603546142578,-18.6946277618408,
-36.1943855285645,-25.2058467864990,
-32.7060432434082,-0.341241240501404,
-26.4782199859619,30.7186603546143,
-39.5718727111816,36.9676437377930,
-70.2228393554688,22.2303676605225,
-81.4267501831055,13.9879455566406,
-39.4335021972656,19.2722511291504,
25.7904262542725,14.8968200683594,
53.1293525695801,-4.42853927612305,
24.7775783538818,-15.7035684585571,
-14.4887609481812,-11.8608207702637,
-20.9087543487549,-18.4942626953125,
-4.21651649475098,-52.0007934570313,
0.730925977230072,-80.6760177612305,
-11.7743368148804,-57.5523185729981,
-18.5852069854736,7.74770116806030,
-13.2610359191895,49.7032470703125,
-14.4799499511719,30.6790103912354,
-30.3306980133057,-15.2207584381104,
-36.8455848693848,-31.4910774230957,
-15.6303920745850,-5.73636484146118,
19.6612663269043,25.4848537445068,
37.1301803588867,25.9218521118164,
28.1632556915283,2.25644516944885,
14.6773843765259,-15.1758060455322,
6.71079349517822,-6.99248886108398,
-0.481546044349670,13.8663024902344,
-8.34572219848633,17.7612743377686,
-13.2857770919800,-10.5282382965088,
-13.6197528839111,-52.4257888793945,
-13.9708700180054,-64.3304977416992,
-19.1372566223145,-26.2508602142334,
-23.1712894439697,28.8771686553955,
-19.9302730560303,43.1707763671875,
-9.61044502258301,3.69558691978455,
7.54902791976929,-44.4478187561035,
36.2112464904785,-52.8673553466797,
61.7872619628906,-20.5535736083984,
52.7134857177734,13.9165296554565,
3.97130298614502,23.6430816650391,
-38.8704185485840,19.1126937866211,
-35.1436157226563,11.8803167343140,
-0.120684623718262,0.298309683799744,
16.6733951568604,-16.5471153259277,
4.24534702301025,-27.0646133422852,
1.97280526161194,-19.4875106811523,
32.5885086059570,-5.87085914611816,
57.4945678710938,-7.65670967102051,
35.8183898925781,-25.3684864044189,
-5.97391891479492,-35.2753257751465,
-9.07309341430664,-25.6606044769287,
25.5873146057129,-6.82882499694824,
40.5073165893555,5.01709938049316,
15.9920444488525,11.1451396942139,
-5.11236286163330,24.3486843109131,
13.5066280364990,45.9749603271484,
38.2999076843262,55.9309158325195,
20.9386615753174,40.4200859069824,
-19.1723346710205,4.97343492507935,
-24.5199680328369,-30.4430961608887,
12.7891349792480,-47.1088562011719,
41.0121459960938,-36.2635231018066,
30.9294567108154,-8.23400497436523,
12.8065013885498,18.4524497985840,
18.7356700897217,32.3692436218262,
24.4560832977295,34.6209754943848,
-3.69898080825806,32.3520393371582,
-37.9327011108398,27.1934661865234,
-24.7133064270020,18.9314918518066,
31.3972854614258,16.4364833831787,
62.8126640319824,34.6637344360352,
24.6130523681641,62.6376495361328,
-44.8463211059570,63.5346603393555,
-68.4690628051758,22.8254718780518,
-25.1410846710205,-19.3658447265625,
28.2831974029541,-17.3973712921143,
33.6103515625000,27.1086959838867,
-10.2738895416260,61.0740585327148,
-57.2323493957520,48.5620040893555,
-68.2261199951172,10.6120471954346,
-45.9639549255371,-22.1529541015625,
-23.0260639190674,-46.2451705932617,
-19.5769195556641,-74.1309814453125,
-22.3392562866211,-88.2493438720703,
-9.87048053741455,-57.5613822937012,
15.0899648666382,0.905944824218750,
27.3264389038086,29.8600997924805,
12.5952959060669,6.01410579681397,
-9.94895839691162,-25.2888393402100,
-10.1988706588745,-15.1898651123047,
16.9395313262939,29.2974376678467,
38.4948806762695,60.3948516845703,
34.7934722900391,52.7405204772949,
15.2335319519043,21.6462421417236,
0.0756206512451172,-10.3991279602051,
-7.93522739410400,-40.5465736389160,
-19.9526824951172,-65.4748840332031,
-32.7980804443359,-69.0564422607422,
-19.5186252593994,-56.4598579406738,
22.4932479858398,-51.1661071777344,
58.4939765930176,-50.3120765686035,
48.7396697998047,-28.7409687042236,
1.42510819435120,18.7668838500977,
-36.6077117919922,41.5061645507813,
-31.8569374084473,5.30551147460938,
-7.02925252914429,-49.6979560852051,
-3.46036982536316,-52.3558158874512,
-26.1820087432861,-3.44377994537354,
-42.3393058776856,25.8757801055908,
-27.4134502410889,-8.97006797790527,
1.98900961875916,-53.6501274108887,
9.18240356445313,-39.0387954711914,
-11.5930490493774,16.1352958679199,
-32.2209129333496,35.5510711669922,
-26.2738838195801,-6.33408117294312,
-6.05841588973999,-54.7339057922363,
-3.18092679977417,-56.6103935241699,
-23.6953296661377,-18.0623035430908,
-39.5002326965332,16.4948787689209,
-19.8326301574707,24.8297290802002,
30.6898536682129,19.1050739288330,
65.5124435424805,15.9410228729248,
51.1652221679688,26.0994434356689,
5.99284219741821,51.3490219116211,
-28.6134185791016,73.1425552368164,
-28.1040115356445,59.1199226379395,
-7.77294206619263,2.72784662246704,
8.75671768188477,-46.1838378906250,
23.2600193023682,-36.5076179504395,
44.6997947692871,14.4835329055786,
59.8543319702148,43.4611320495606,
40.3037719726563,27.2009525299072,
-9.60964012145996,8.05986309051514,
-48.5183639526367,21.7034912109375,
-49.1585273742676,41.0708923339844,
-33.7549934387207,12.9232225418091,
-37.2778053283691,-47.3666076660156,
-51.6676101684570,-72.0124511718750,
-37.6530952453613,-31.8324127197266,
12.9133691787720,22.3655300140381,
58.0592994689941,33.7912864685059,
61.4627380371094,8.34099864959717,
30.4084453582764,-14.4003267288208,
-0.00258708000183105,-11.9847450256348,
-18.0784893035889,4.20918178558350,
-31.4100894927979,20.7469081878662,
-31.9837932586670,22.9293441772461,
-10.6498336791992,4.03633880615234,
17.8631439208984,-30.1387786865234,
25.5332584381104,-54.8418235778809,
13.7642621994019,-48.3804931640625,
15.4983549118042,-29.3551368713379,
45.0086784362793,-31.9718856811523,
75.4966812133789,-45.9300613403320,
74.8557434082031,-26.0268306732178,
53.5532989501953,22.7026100158691,
34.1019744873047,39.1022567749023,
18.2435379028320,-1.37152791023254,
-13.1000480651855,-44.6038284301758,
-45.2682838439941,-31.8122863769531,
-39.0652427673340,7.95527505874634,
7.42945241928101,4.53244686126709,
43.1229553222656,-41.6381530761719,
19.5003604888916,-51.2932701110840,
-38.7825164794922,-1.92272806167603,
-65.1480865478516,33.7164421081543,
-32.0455017089844,0.408576846122742,
17.7247505187988,-49.2921600341797,
27.7654018402100,-29.1016445159912,
-1.41963529586792,39.0049057006836,
-23.6439895629883,60.4415245056152,
-6.31864547729492,4.06078720092773,
30.1735992431641,-50.1431236267090,
55.2640914916992,-33.5316352844238,
60.4089202880859,23.1097126007080,
59.0248260498047,48.6394042968750,
52.1717185974121,34.0651016235352,
28.6539592742920,32.2688293457031,
-10.6408405303955,63.3279647827148,
-40.0977172851563,84.2861862182617,
-33.3618545532227,58.8646240234375,
-6.02091312408447,6.96388387680054,
8.13382816314697,-32.5101737976074,
2.23694157600403,-47.6159820556641,
-1.86998081207275,-45.6853065490723,
16.3929538726807,-38.5128021240234,
39.7823448181152,-31.9006900787354,
35.9236450195313,-23.4303207397461,
4.31719732284546,-9.54331016540527,
-17.2220401763916,9.58781909942627,
-2.95717287063599,25.5121059417725,
21.2186565399170,21.3751525878906,
15.7369813919067,-8.78914070129395,
-19.2816314697266,-33.6118431091309,
-33.0133171081543,-27.2927989959717,
2.19418048858643,-7.89942789077759,
53.7813148498535,-4.20329570770264,
61.8978118896484,-6.66720247268677,
18.3981742858887,15.6980180740356,
-24.6640052795410,57.2174186706543,
-29.0078182220459,66.3655853271484,
-18.6184082031250,19.3468341827393,
-25.0139026641846,-31.1893482208252,
-33.0034561157227,-31.0617179870605,
-8.47402858734131,4.23963165283203,
38.1880645751953,7.95030260086060,
58.0137863159180,-26.1827335357666,
35.7430686950684,-35.5666809082031,
7.23504066467285,12.0130195617676,
0.761706173419952,63.2296104431152,
-4.12931919097900,52.2737350463867,
-26.5614280700684,-0.361169457435608,
-37.7253379821777,-15.6785678863525,
-7.39270401000977,28.1382446289063,
30.4323024749756,75.0052032470703,
16.0051422119141,67.1607055664063,
-39.7784614562988,17.8983020782471,
-66.1782379150391,-25.1234340667725,
-33.5480346679688,-45.4880752563477,
4.18967390060425,-61.8018379211426,
-3.36059474945068,-72.9380111694336,
-26.7613735198975,-56.1748657226563,
-10.7412786483765,-10.0796813964844,
39.3333663940430,29.1649570465088,
65.2573471069336,29.7441787719727,
47.1539573669434,2.73021316528320,
27.8265285491943,-17.1499652862549,
31.2829532623291,-7.60230064392090,
27.6525211334229,21.9581298828125,
-3.94795608520508,45.4262390136719,
-32.8152618408203,51.3190650939941,
-19.2975730895996,40.7995452880859,
22.0407638549805,20.4396820068359,
45.7509384155273,-0.761961102485657,
40.2051086425781,-8.52270889282227,
26.4367008209229,1.20829892158508,
16.7345943450928,22.7634353637695,
-3.89275693893433,40.8029937744141,
-34.6568183898926,37.6092453002930,
-46.9769668579102,4.43766355514526,
-25.8750953674316,-33.8195571899414,
2.06291627883911,-45.5498962402344,
2.66530609130859,-25.7418937683105,
-10.4706029891968,-1.99254679679871,
-4.25838613510132,-3.38631367683411,
25.4768486022949,-20.7168178558350,
43.5917549133301,-19.9894695281982,
24.6127262115479,1.11521852016449,
-13.7977466583252,6.93540763854981,
-30.0841197967529,-20.1280269622803,
-13.5282306671143,-40.9529037475586,
8.63077163696289,-10.5735597610474,
6.88588476181030,44.3822021484375,
-16.2569637298584,55.3277511596680,
-28.0434150695801,1.30927324295044,
-5.15178537368774,-54.7521553039551,
38.8282051086426,-46.1749954223633,
66.7919616699219,5.41935253143311,
50.3012199401856,30.1066875457764,
4.46755504608154,8.73660850524902,
-27.0381870269775,-12.3971347808838,
-19.0885791778564,4.94204807281494,
12.3924932479858,39.5025520324707,
28.5976696014404,51.9126663208008,
6.45505285263062,46.8171043395996,
-38.7476310729981,47.8786048889160,
-68.4271011352539,47.3413162231445,
-60.8004646301270,17.2862129211426,
-26.5475749969482,-36.0177268981934,
6.80769777297974,-63.4158020019531,
14.8781938552856,-36.4172477722168,
-5.41039991378784,16.9404392242432,
-30.8407192230225,37.8319473266602,
-33.1527557373047,12.4491720199585,
-1.20560765266418,-16.9138469696045,
39.9112777709961,-12.2937126159668,
48.3035926818848,22.5493354797363,
16.8637580871582,51.9114990234375,
-23.0227241516113,41.4938583374023,
-35.2770881652832,-4.81756734848023,
-16.9982414245605,-48.3387298583984,
0.673878431320190,-52.3361015319824,
2.98030185699463,-20.5734081268311,
3.50451040267944,10.9007825851440,
11.0024518966675,15.3609504699707,
14.2466468811035,6.31134510040283,
3.00153160095215,13.3899660110474,
-18.4628028869629,36.1403236389160,
-34.5838584899902,36.3382301330566,
-39.0197944641113,0.209789395332336,
-30.9968223571777,-31.3208427429199,
-5.26788949966431,-17.4391269683838,
26.6630821228027,27.6712207794189,
33.7509117126465,50.3565444946289,
-3.26608872413635,25.6835155487061,
-50.5344276428223,-17.9715995788574,
-48.3153610229492,-40.2046623229981,
6.02110052108765,-36.1293640136719,
44.5189056396484,-18.4992256164551,
21.2004432678223,10.3567571640015,
-27.4173259735107,44.2609939575195,
-40.1279487609863,58.9888687133789,
-11.0763731002808,32.4307937622070,
10.8423662185669,-10.6470403671265,
0.491533637046814,-21.0695457458496,
-15.2673740386963,7.68723773956299,
-15.3465242385864,29.6364765167236,
-19.5628643035889,17.2773761749268,
-40.4346885681152,-3.20126962661743,
-48.6156539916992,1.04509294033051,
-24.2668685913086,20.2940464019775,
1.79745435714722,19.1099166870117,
-6.72523307800293,-4.82202529907227,
-24.6305236816406,-12.3654689788818,
-9.79621791839600,11.1462316513062,
17.9492073059082,34.2173957824707,
3.22513341903687,35.2134437561035,
-53.4211807250977,27.9973239898682,
-79.2221145629883,25.6554946899414,
-31.2274208068848,19.4833850860596,
30.9321022033691,4.83691406250000,
35.3439140319824,3.79679846763611,
2.61213684082031,26.3591880798340,
4.66287040710449,37.9719886779785,
40.1785011291504,4.99385070800781,
50.4084777832031,-41.3263549804688,
21.0022239685059,-39.2975463867188,
8.08447837829590,11.6712007522583,
36.2993698120117,39.3837432861328,
56.2640419006348,7.22790193557739,
22.7254161834717,-32.3632621765137,
-23.5598983764648,-20.2454128265381,
-19.9733638763428,16.4194126129150,
17.8642311096191,9.32467269897461,
21.0716438293457,-39.8621978759766,
-24.5910873413086,-58.0188369750977,
-59.5547676086426,-9.29464817047119,
-48.6030845642090,51.6937065124512,
-34.0690002441406,53.6627311706543,
-52.0217742919922,0.745662689208984,
-69.9071807861328,-43.0015792846680,
-48.3256530761719,-46.2831726074219,
-5.53440189361572,-34.3479728698731,
8.24760532379150,-36.3098640441895,
-18.2700920104980,-44.4255180358887,
-42.2914047241211,-39.3383064270020,
-33.6085357666016,-18.9931297302246,
-5.77384948730469,0.454294323921204,
16.9517288208008,5.10915374755859,
37.7116241455078,-5.17649173736572,
59.0350837707520,-12.5866098403931,
65.0651473999023,0.684975981712341,
50.1330184936523,33.7857437133789,
29.3284454345703,60.7283554077148,
13.5225343704224,52.6080932617188,
-9.83052635192871,7.95558547973633,
-43.4219207763672,-32.0654296875000,
-60.2492942810059,-31.9011650085449,
-35.6630287170410,-2.85653185844421,
9.26117229461670,16.0577106475830,
26.1593036651611,7.28097581863403,
7.14181566238403,-11.8110904693604,
-7.27874660491943,-25.6769771575928,
10.6694202423096,-31.1274929046631,
32.0199890136719,-35.2490348815918,
20.2614803314209,-30.4038944244385,
-8.37528610229492,-12.7078275680542,
-8.43351650238037,4.69704008102417,
29.1203899383545,5.27725410461426,
62.8210868835449,-3.17044472694397,
58.3889579772949,2.28851842880249,
22.6058940887451,24.2363357543945,
-10.2781047821045,43.1085662841797,
-26.2930488586426,42.7873458862305,
-32.7072029113770,36.6504211425781,
-36.1109733581543,32.4571914672852,
-38.0220298767090,17.0026721954346,
-37.1833114624023,-19.8392448425293,
-30.8132286071777,-59.8014793395996,
-8.85593318939209,-72.1021423339844,
25.8046321868897,-53.0499038696289,
44.8695144653320,-29.8479099273682,
23.1463356018066,-20.8126850128174,
-20.9382610321045,-15.3154315948486,
-42.5591697692871,0.153535962104797,
-20.1311588287354,13.3648748397827,
15.8013820648193,10.6131153106689,
24.7774753570557,-0.435352087020874,
3.97666072845459,-11.6786403656006,
-9.81255149841309,-24.4005413055420,
-1.74149870872498,-41.1974639892578,
13.5110225677490,-44.3993949890137,
18.6069965362549,-24.6962337493897,
14.6239166259766,1.04416465759277,
9.74178791046143,1.61830484867096,
2.17905926704407,-13.6422948837280,
-8.06098747253418,-4.71491622924805,
-7.09937095642090,32.3111228942871,
11.6397142410278,43.8836250305176,
33.4617881774902,4.99279975891113,
38.0827102661133,-35.9717788696289,
28.6146564483643,-15.1670541763306,
25.8719768524170,49.5771980285645,
34.2023010253906,77.0231018066406,
29.9647617340088,36.1559638977051,
0.308229923248291,-19.9154376983643,
-32.3560600280762,-35.4711074829102,
-36.6423339843750,-27.2740745544434,
-16.0963897705078,-40.1949043273926,
3.81109571456909,-63.2638473510742,
4.15804529190064,-46.1303520202637,
-6.49526691436768,14.3342266082764,
-14.5212287902832,54.3119812011719,
-20.0055904388428,30.4820270538330,
-30.0688800811768,-25.0316905975342,
-37.4775161743164,-51.1851196289063,
-32.2836799621582,-30.8394145965576,
-14.2503767013550,12.4492778778076,
4.36751222610474,44.6841201782227,
11.6795835494995,51.7843704223633,
-1.29888737201691,34.0141944885254,
-30.0375614166260,-0.201342433691025,
-52.6137619018555,-31.0691108703613,
-39.7395629882813,-40.6536788940430,
12.8919572830200,-34.9871635437012,
67.1161346435547,-35.0513420104981,
75.8139419555664,-33.9272651672363,
38.2827262878418,-14.4328718185425,
3.78589868545532,12.4289665222168,
14.2127237319946,15.1879005432129,
51.9198112487793,-1.60812079906464,
63.2334976196289,1.09713137149811,
30.2982749938965,40.4527282714844,
-6.74202108383179,76.6849899291992,
-11.2918624877930,60.1511688232422,
6.23852252960205,3.72797250747681,
5.70718288421631,-38.1708526611328,
-20.4078884124756,-48.0786628723145,
-33.1229476928711,-52.2526321411133,
-4.95582580566406,-56.9514389038086,
39.1061325073242,-30.4642982482910,
46.9328460693359,24.9697227478027,
3.59491419792175,50.2507286071777,
-47.5773162841797,10.8049945831299,
-55.9174575805664,-43.2596397399902,
-18.2021713256836,-36.6990928649902,
24.9032020568848,19.7080726623535,
29.6165390014648,46.9339408874512,
-3.35965490341187,15.3911275863647,
-34.4435958862305,-17.9881668090820,
-36.1708106994629,-5.29186153411865,
-16.2949638366699,19.6971359252930,
4.80670738220215,-0.569741725921631,
19.5901317596436,-41.9906959533691,
36.0944671630859,-37.8930282592773,
47.8668937683106,13.8729896545410,
32.0063514709473,49.4430809020996,
-16.2323532104492,26.8278694152832,
-53.4796142578125,-12.6533832550049,
-36.0535697937012,-19.2406902313232,
16.7614059448242,4.35225820541382,
42.1458206176758,16.9519348144531,
18.4334888458252,3.44599962234497,
-12.7967634201050,-11.6902465820313,
-9.23312568664551,-12.2660646438599,
8.68293666839600,-5.53368568420410,
-3.40480279922485,5.10091876983643,
-39.2449951171875,23.7878761291504,
-53.5886993408203,31.8903427124023,
-30.7475166320801,11.8693504333496,
-11.1587495803833,-22.0930442810059,
-22.0104885101318,-41.6320114135742,
-35.8125419616699,-45.3634414672852,
-22.4500637054443,-56.4357070922852,
2.93702483177185,-77.3997344970703,
14.7729473114014,-77.2686767578125,
23.3898258209229,-38.0643577575684,
48.7261848449707,0.661735653877258,
69.1356658935547,-6.10449171066284,
46.3814964294434,-34.1062088012695,
-4.11287498474121,-30.0008316040039,
-26.5473365783691,-0.651077985763550,
-2.38809084892273,0.157621622085571,
18.4841613769531,-39.2212753295898,
-5.19070577621460,-60.7506256103516,
-36.9528846740723,-20.3028945922852,
-25.8285408020020,35.9701194763184,
7.24746751785278,41.1199760437012,
1.68771553039551,5.02981996536255,
-45.2579460144043,-5.27393531799316,
-68.5662384033203,28.2625427246094,
-32.0283813476563,49.9866104125977,
23.8532428741455,27.1908035278320,
40.2094650268555,1.18700897693634,
10.7578830718994,22.9106140136719,
-24.8228034973145,60.1022148132324,
-40.9892921447754,42.3192634582520,
-39.2788543701172,-27.2839717864990,
-23.0188007354736,-71.4997100830078,
11.5293197631836,-37.3361701965332,
44.8997344970703,36.0833854675293,
50.5286102294922,67.8167877197266,
34.4902915954590,36.0705413818359,
22.0372085571289,-5.38251113891602,
17.5960407257080,-5.98814535140991,
4.05440473556519,22.7321548461914,
-13.7106838226318,38.4426269531250,
-7.07406330108643,21.0966815948486,
25.9256916046143,-2.47868061065674,
43.3244323730469,-1.34493362903595,
9.05511093139648,23.6417694091797,
-42.7144927978516,29.7039813995361,
-51.6413803100586,-11.3069667816162,
-17.4973945617676,-71.0574645996094,
-0.107648074626923,-90.9071273803711,
-23.0712203979492,-51.7323455810547,
-42.9476318359375,4.95927858352661,
-15.1852779388428,21.5931682586670,
37.6791152954102,-9.64016723632813,
61.9273300170898,-37.1862602233887,
47.6879158020020,-25.3340511322022,
28.1778373718262,8.56109523773193,
23.2353458404541,33.1903915405273,
16.2346115112305,46.4355545043945,
-6.27891874313355,61.8259506225586,
-29.8215198516846,70.7876815795898,
-40.5522232055664,44.7857284545898,
-46.3171386718750,-7.41571378707886,
-54.7471733093262,-40.0887145996094,
-49.5725860595703,-25.7649250030518,
-16.0926418304443,4.49157905578613,
20.0410594940186,2.85332918167114,
25.7147045135498,-23.0596885681152,
2.45058822631836,-29.2418613433838,
-16.5646553039551,5.41190528869629,
-11.0194969177246,42.1069335937500,
-0.472455441951752,39.4618415832520,
-7.85985183715820,7.57242155075073,
-23.4005317687988,-18.2104244232178,
-21.4163093566895,-16.8583679199219,
1.87367582321167,6.25240850448608,
20.1714267730713,36.7773094177246,
17.4088420867920,61.2225151062012,
-5.80640411376953,56.9782638549805,
-39.4907226562500,13.4059658050537,
-60.4719810485840,-50.3508872985840,
-47.4870986938477,-87.6329040527344,
1.48951923847198,-76.4586181640625,
45.5012359619141,-38.9933586120606,
40.4402008056641,-6.51805210113525,
-12.7808856964111,11.1918020248413,
-62.5403976440430,12.8336553573608,
-64.1136245727539,-7.01986789703369,
-29.6197681427002,-43.6897087097168,
5.15701627731323,-67.2982254028320,
34.8446960449219,-55.8582153320313,
68.7550201416016,-21.8291702270508,
85.6432876586914,-5.13683176040649,
55.6247100830078,-12.0608959197998,
-5.61078405380249,-10.9466400146484,
-45.2917213439941,17.8354225158691,
-38.0056915283203,49.5801124572754,
-14.3481512069702,52.2604598999023,
-8.90549659729004,35.0362167358398,
-5.22779083251953,27.1806297302246,
20.1091346740723,30.2496013641357,
43.1533393859863,22.3930473327637,
23.2969284057617,-6.15807008743286,
-20.9069938659668,-31.9435653686523,
-29.9544048309326,-36.3865509033203,
6.62266063690186,-33.2278938293457,
27.7591056823730,-39.3244361877441,
-0.684744119644165,-47.7230606079102,
-34.6032524108887,-42.1507759094238,
-15.7074661254883,-29.3304443359375,
27.8294429779053,-30.7869548797607,
28.7760391235352,-47.4592666625977,
-18.2882499694824,-48.5170631408691,
-43.5405464172363,-14.7176074981689,
-7.98105382919312,31.5819530487061,
35.1977500915527,54.2288208007813,
19.2634277343750,33.5877571105957,
-38.3574714660645,-10.9187316894531,
-60.5227050781250,-49.5001907348633,
-19.1129055023193,-66.4628829956055,
30.3452701568604,-64.9580230712891,
32.7694358825684,-52.3649024963379,
0.231372475624084,-33.6152992248535,
-11.6833581924438,-14.5280647277832,
17.3462142944336,-0.575486063957214,
48.1727790832520,-1.02623033523560,
40.1958961486816,-18.7584438323975,
6.23957681655884,-37.4419250488281,
-6.76809835433960,-30.8286323547363,
13.4419040679932,9.89348411560059,
37.2349510192871,53.9816932678223,
30.6965560913086,60.1417770385742,
1.78693318367004,23.9919548034668,
-13.7040576934814,-15.6150436401367,
-3.22396039962769,-17.9414348602295,
8.24454975128174,10.9823627471924,
-3.74204730987549,32.8313140869141,
-25.0971240997314,29.5789852142334,
-30.0939292907715,14.5875062942505,
-16.3993587493897,9.92150402069092,
-2.80528974533081,8.03900718688965,
-1.91475367546082,-5.76051092147827,
-0.691242456436157,-31.0210285186768,
18.1646823883057,-46.5614433288574,
48.7244377136231,-35.4858703613281,
65.6840515136719,-4.51513719558716,
59.5847167968750,26.2482128143311,
39.6445426940918,37.8869056701660,
17.1516780853272,28.0054054260254,
-8.39936256408691,2.92472600936890,
-34.4299087524414,-24.1990108489990,
-40.3875083923340,-41.1220283508301,
-14.4026823043823,-46.5799026489258,
23.7095832824707,-46.9304199218750,
31.1857757568359,-38.5058403015137,
-2.03883886337280,-13.1013221740723,
-33.2684783935547,19.4899063110352,
-23.7821254730225,32.6315612792969,
9.36555099487305,13.4912157058716,
13.6865701675415,-13.0322980880737,
-21.6065654754639,-14.2818813323975,
-52.9445838928223,5.14754915237427,
-48.1932144165039,3.39640259742737,
-28.9651317596436,-38.3619308471680,
-27.6983680725098,-79.8070983886719,
-30.6613445281982,-74.6111679077148,
2.27424550056458,-34.3240699768066,
60.9393043518066,-8.01404190063477,
85.7597427368164,-13.3804626464844,
47.2896499633789,-23.7533302307129,
-11.0447654724121,-15.6927995681763,
-32.1786842346191,2.44885849952698,
-14.4254684448242,14.8358039855957,
3.05117821693420,22.8619308471680,
4.17226934432983,28.1068744659424,
7.99478149414063,14.9104871749878,
17.7580013275147,-20.5768623352051,
14.1825189590454,-43.3996162414551,
-12.5915832519531,-24.4587688446045,
-35.7760963439941,5.43591594696045,
-26.9541816711426,-3.80168795585632,
1.06766402721405,-41.5656013488770,
17.6446800231934,-49.2652511596680,
14.7445755004883,-9.93661594390869,
17.5724086761475,31.7567958831787,
36.7279319763184,37.5405807495117,
45.5031089782715,31.5016975402832,
20.5218334197998,48.2622184753418,
-26.5591030120850,63.2610702514648,
-55.6322708129883,33.0807342529297,
-38.8584861755371,-15.5155735015869,
8.03599548339844,-16.0374450683594,
46.6617050170898,32.9975662231445,
56.9281997680664,55.1915817260742,
43.3597106933594,12.2102527618408,
20.7962226867676,-36.2272605895996,
-3.61399364471436,-20.7584590911865,
-28.3260498046875,30.0988845825195,
-47.3682556152344,42.4090385437012,
-47.2132301330566,5.75586700439453,
-22.5156955718994,-16.1243743896484,
7.64868879318237,14.5621623992920,
12.0194301605225,51.1106376647949,
-18.2328872680664,36.6894340515137,
-50.2307510375977,-15.1779270172119,
-41.4308776855469,-49.7469596862793,
11.8795900344849,-46.2042465209961,
65.1004409790039,-26.2121696472168,
69.6830520629883,-5.41454935073853,
30.8144474029541,16.4238071441650,
-6.77036714553833,35.3933906555176,
-11.0667343139648,39.1641731262207,
5.36178016662598,31.8174877166748,
8.32023143768311,29.8906383514404,
-8.32478427886963,38.0961303710938,
-26.7184123992920,40.1675720214844,
-28.1915512084961,19.3870277404785,
-16.3624572753906,-7.60055351257324,
-6.13551616668701,-20.5785331726074,
-9.00763416290283,-25.1696434020996,
-19.3443527221680,-37.7483940124512,
-26.4092063903809,-49.0872573852539,
-23.0053119659424,-41.0148162841797,
-14.6358880996704,-12.7958889007568,
-11.2289628982544,12.1656312942505,
-13.4012804031372,15.3356294631958,
-7.57680845260620,1.92978942394257,
16.0756645202637,-13.1825485229492,
31.6226959228516,-21.7964229583740,
11.4383068084717,-16.6413478851318,
-30.5059165954590,7.78138542175293,
-46.6673622131348,45.1441078186035,
-17.1117134094238,62.9984207153320,
17.2495727539063,42.2885131835938,
3.68000984191895,7.82258510589600,
-44.2405624389648,0.226439118385315,
-63.7624549865723,21.2624988555908,
-29.2546806335449,38.5699615478516,
15.1242990493774,35.9267501831055,
21.9205856323242,33.4758682250977,
4.42797279357910,45.4393539428711,
7.85496377944946,52.6713752746582,
31.5193614959717,30.2007350921631,
38.8028030395508,-8.49457740783691,
16.8018188476563,-27.3635807037354,
-1.73746275901794,-25.4743995666504,
6.99820899963379,-30.7797298431397,
21.6763439178467,-43.9430465698242,
8.57645606994629,-33.6499099731445,
-25.8388576507568,7.18430900573731,
-46.4756202697754,38.9220504760742,
-35.7347946166992,28.9455184936523,
-10.6373701095581,3.57369732856751,
12.2957801818848,4.00101184844971,
24.7229804992676,24.2198314666748,
12.6492042541504,25.8581809997559,
-21.9358501434326,3.30192947387695,
-52.4318771362305,-0.805946111679077,
-50.5046501159668,25.0479373931885,
-22.3143997192383,40.4325942993164,
-4.12776803970337,10.5644044876099,
-6.45708322525024,-31.8678264617920,
-0.500279426574707,-35.8875083923340,
30.3512878417969,-7.26500082015991,
52.4732704162598,7.24100017547607,
30.6028804779053,-9.00110530853272,
-6.06962490081787,-23.3917102813721,
0.432915806770325,-12.8930263519287,
44.6178894042969,6.61397838592529,
56.8313140869141,7.83383417129517,
6.46609354019165,0.586879611015320,
-53.7371520996094,11.7933816909790,
-56.5178985595703,38.4592132568359,
-9.09557056427002,51.8562088012695,
28.9586162567139,42.4610748291016,
25.5490989685059,21.8476696014404,
1.31414377689362,0.0932804644107819,
-16.1664180755615,-18.1192550659180,
-28.2006034851074,-26.4732227325439,
-33.9356651306152,-27.7104492187500,
-20.7180957794189,-32.6602516174316,
3.76787900924683,-44.8247184753418,
12.2237367630005,-44.0424423217773,
-3.18353056907654,-6.29719400405884,
-6.49929857254028,46.8274345397949,
21.8792114257813,59.5617294311523,
51.5282325744629,14.6694593429565,
40.0511474609375,-28.3168430328369,
3.39067220687866,-10.7660093307495,
-5.62162780761719,35.9520606994629,
23.9181404113770,36.8484153747559,
41.4897613525391,-15.0074911117554,
10.8875141143799,-48.6330375671387,
-27.9142913818359,-11.4450807571411,
-19.6798057556152,50.0356712341309,
27.0457172393799,59.1848526000977,
53.6813087463379,11.2767753601074,
30.8917446136475,-32.7294616699219,
-7.84988784790039,-30.7105121612549,
-26.5460624694824,-5.84225511550903,
-26.4565010070801,12.7366685867310,
-32.0476608276367,21.5416526794434,
-45.4247589111328,25.8418312072754,
-45.9833297729492,11.4269456863403,
-19.3187656402588,-25.2799510955811,
21.1998310089111,-49.6843719482422,
55.8707313537598,-32.9471206665039,
69.2109832763672,10.8938055038452,
53.1271705627441,41.3192405700684,
18.8686447143555,39.2769966125488,
-5.83679294586182,21.3115634918213,
-9.83985614776611,3.67268109321594,
-10.0910949707031,-20.1873817443848,
-17.8923797607422,-46.8536109924316,
-17.1561927795410,-48.8365516662598,
7.98178577423096,-15.4947338104248,
43.2600173950195,25.7828464508057,
48.2189216613770,41.1400375366211,
20.9428062438965,29.9445686340332,
10.7899074554443,13.9379472732544,
43.2121391296387,5.45085096359253,
73.6677017211914,-5.53033971786499,
45.8113861083984,-16.9672164916992,
-14.2709188461304,-14.1949014663696,
-36.6580162048340,5.36867046356201,
-3.00263786315918,19.3935050964355,
21.8507099151611,4.34885644912720,
-5.02599859237671,-22.7156028747559,
-37.8198242187500,-33.0819015502930,
-12.5049457550049,-17.0430927276611,
53.0696983337402,4.44990587234497,
80.5763854980469,11.9221506118774,
40.3626976013184,4.32513093948364,
-11.9403438568115,-11.4529209136963,
-21.0277214050293,-28.9437980651855,
-2.76662778854370,-43.2495155334473,
1.07697618007660,-51.0784912109375,
-5.85719347000122,-49.3796615600586,
8.66763496398926,-42.3687362670898,
46.8181114196777,-28.6333312988281,
66.5199661254883,0.163878440856934,
45.0566291809082,41.1988754272461,
-1.61337065696716,68.8633804321289,
-32.7761993408203,66.6711807250977,
-30.1018676757813,47.8523406982422,
-3.82520198822022,36.1751289367676,
28.1123847961426,34.6835098266602,
45.0896301269531,30.2968025207520,
32.1533012390137,27.3651065826416,
3.04501724243164,40.2574806213379,
-4.33787727355957,61.6287384033203,
20.3215408325195,56.6693267822266,
45.8110656738281,11.6006431579590,
38.3101768493652,-30.0925235748291,
4.21366834640503,-22.8321857452393,
-26.4581756591797,15.0584678649902,
-40.4508132934570,22.1543636322022,
-50.9730377197266,-17.3475131988525,
-58.9813957214356,-54.2681503295898,
-41.8209838867188,-46.1258163452148,
3.70882511138916,-11.7030458450317,
37.1965599060059,17.1333999633789,
27.4937610626221,36.7651405334473,
-4.24382734298706,60.8657836914063,
-16.7682800292969,68.7425918579102,
-6.56251525878906,30.9943237304688,
-1.92962443828583,-32.2374343872070,
-7.47034978866577,-52.8799781799316,
-3.25558352470398,-11.0606412887573,
11.8268299102783,39.1696624755859,
4.46430873870850,38.7867813110352,
-35.4067459106445,-1.47193682193756,
-64.3910827636719,-32.1092033386231,
-37.2427406311035,-36.2646980285645,
19.1955738067627,-28.5301513671875,
43.0031738281250,-11.8984565734863,
21.8315219879150,19.1126022338867,
1.07718288898468,48.4262161254883,
11.4477243423462,41.7144393920898,
22.9419021606445,2.25496387481689,
3.66580057144165,-16.8770751953125,
-23.4261245727539,14.1588153839111,
-13.9743652343750,57.0041732788086,
26.7793445587158,56.9015884399414,
47.8299484252930,19.7228794097900,
24.3291854858398,-1.65211701393127,
-10.2209281921387,13.8640270233154,
-12.9351196289063,39.4428291320801,
4.10395526885986,43.2326545715332,
-2.56639957427979,25.7126693725586,
-37.9312896728516,2.85146379470825,
-60.8103523254395,-18.2365226745605,
-38.3658638000488,-36.0326271057129,
13.0331935882568,-33.8115806579590,
41.1685523986816,-7.23121881484985,
18.4108943939209,17.7072849273682,
-21.7481155395508,9.82434654235840,
-29.5398941040039,-25.0722064971924,
3.78558826446533,-48.3673286437988,
35.2717781066895,-44.3338470458984,
19.9043235778809,-28.6236820220947,
-32.7147026062012,-19.9910163879395,
-64.5158767700195,-23.3269081115723,
-39.9358520507813,-28.6589393615723,
6.38231658935547,-29.2423553466797,
13.5302238464355,-18.7002105712891,
-25.5248603820801,5.23730325698853,
-57.0738143920898,36.3956298828125,
-35.1937065124512,48.4584693908691,
14.3654346466064,32.8267631530762,
28.3722000122070,9.80539894104004,
-12.6701278686523,0.392065554857254,
-55.3447265625000,-8.56503772735596,
-46.8254470825195,-39.5501365661621,
0.507684707641602,-72.0271911621094,
29.4536628723145,-64.6859893798828,
10.1178359985352,-17.9093551635742,
-24.8963623046875,22.7367877960205,
-31.7708663940430,22.9216880798340,
-15.5079956054688,8.34883975982666,
-14.0488872528076,18.5618495941162,
-31.9073905944824,41.6034393310547,
-38.9288558959961,30.3632144927979,
-12.0580387115479,-14.0674381256104,
22.0091571807861,-45.6537704467773,
22.6379203796387,-41.1136512756348,
-6.55670595169067,-28.3474349975586,
-18.6249408721924,-33.7877426147461,
5.27215480804443,-31.6296215057373,
33.1177940368652,-0.434577941894531,
25.3947811126709,29.2722816467285,
-8.79674625396729,12.8089799880981,
-27.3278770446777,-29.3680419921875,
-13.8347845077515,-36.8245277404785,
-0.865056514739990,6.77733039855957,
-16.4788284301758,40.2235260009766,
-48.2603225708008,10.9244689941406,
-62.6919364929199,-45.8270568847656,
-47.8037414550781,-66.1012191772461,
-23.6111278533936,-43.9721565246582,
-11.4671068191528,-26.2950248718262,
-13.7848548889160,-36.7558364868164,
-14.6121053695679,-55.6754112243652,
-2.05538845062256,-57.9154548645020,
22.0120563507080,-43.6442527770996,
45.1986351013184,-27.0056076049805,
57.3617362976074,-11.4347877502441,
53.8365440368652,-5.66290664672852,
42.6745948791504,-17.7335491180420,
34.7345008850098,-36.2455177307129,
32.5051689147949,-22.6785964965820,
31.7654895782471,28.3293476104736,
26.4885978698730,64.6570358276367,
16.9529514312744,41.6478805541992,
5.54693126678467,-9.04034900665283,
-4.40151977539063,-23.5604038238525,
-13.8866291046143,4.11327648162842,
-25.8726844787598,23.2676353454590,
-39.4786605834961,1.55662655830383,
-39.2279396057129,-25.6170806884766,
-13.6504678726196,-16.7906112670898,
27.0903263092041,14.0630874633789,
52.1050338745117,23.3120956420898,
44.1797370910645,18.6571941375732,
21.4557266235352,33.5040473937988,
13.7988576889038,64.8021926879883,
19.4776954650879,70.9262771606445,
9.89313793182373,40.8488311767578,
-19.8070049285889,14.8140716552734,
-31.3998031616211,13.5683441162109,
1.94984555244446,10.3059730529785,
49.3899116516113,-15.0279455184937,
53.4898338317871,-32.3148269653320,
5.16553974151611,-9.74498081207275,
-43.8593101501465,27.3807163238525,
-45.5536041259766,22.0248508453369,
-14.5512504577637,-25.0403327941895,
1.53493237495422,-47.1051216125488,
-3.58716034889221,-12.0822029113770,
-1.44928455352783,33.8129768371582,
23.5987071990967,39.9441032409668,
45.8615570068359,15.4474868774414,
35.9652252197266,-5.55952310562134,
7.51215171813965,-16.5045108795166,
-5.53267860412598,-30.2243022918701,
-2.58753347396851,-42.7807426452637,
-7.93779468536377,-38.9670028686523,
-23.0293254852295,-34.2323341369629,
-17.1239452362061,-48.7544441223145,
22.6513328552246,-63.9357986450195,
57.0074806213379,-35.4764976501465,
35.9926795959473,30.2539272308350,
-23.4114952087402,63.4302291870117,
-50.3001747131348,27.8024921417236,
-14.4958095550537,-23.2519569396973,
38.0446128845215,-27.6919918060303,
44.0525741577148,-0.626497149467468,
6.59972810745239,4.48744630813599,
-13.6728363037109,-16.7429809570313,
14.5076007843018,-16.4122848510742,
58.3414802551270,28.4950866699219,
63.7857208251953,74.0907058715820,
29.0757865905762,79.6438903808594,
-3.48068046569824,62.1711120605469,
-4.51665210723877,50.3118476867676,
11.0783290863037,33.9713249206543,
16.2009773254395,-0.442966938018799,
0.411440610885620,-24.5566539764404,
-22.9426116943359,-5.84946393966675,
-33.8915557861328,25.7668094635010,
-35.4720497131348,18.0841140747070,
-34.0058898925781,-19.7675762176514,
-28.1949501037598,-29.7639293670654,
-19.6314277648926,5.05899190902710,
-18.5049285888672,27.3946208953857,
-33.5227394104004,-7.73626279830933,
-53.1525421142578,-53.7374420166016,
-46.8694610595703,-39.0172042846680,
-8.67298030853272,22.5805053710938,
24.1343917846680,55.7570419311523,
5.76872491836548,37.7171096801758,
-45.9566268920898,19.8611202239990,
-65.6910171508789,28.6084671020508,
-15.7504415512085,28.9308223724365,
60.0452766418457,-3.00721216201782,
88.6814346313477,-33.3444023132324,
54.3685188293457,-20.8454055786133,
4.50125360488892,13.6250839233398,
-20.7046413421631,21.8495483398438,
-18.1852817535400,4.55307340621948,
-5.94419527053833,4.94694805145264,
5.47794246673584,24.6805763244629,
9.79445171356201,19.2471733093262,
-4.37943458557129,-16.8233585357666,
-33.7070198059082,-32.8652839660645,
-51.7392234802246,-10.3324537277222,
-44.3751068115234,4.08906698226929,
-28.9376506805420,-24.3944778442383,
-25.8891162872314,-50.7968864440918,
-22.4705562591553,-20.9337120056152,
-4.81578779220581,40.6991233825684,
6.32599973678589,59.8500823974609,
-15.0159854888916,23.2162303924561,
-47.1336860656738,-2.65125250816345,
-43.6499671936035,23.5144710540772,
-0.777389049530029,55.7091255187988,
18.9400177001953,44.5226860046387,
-22.2514934539795,15.4007196426392,
-77.1675415039063,13.4198150634766,
-74.8265075683594,27.0145626068115,
-23.3813152313232,11.0758876800537,
7.01499509811401,-35.2372436523438,
-12.3996257781982,-67.0529403686523,
-29.7311382293701,-65.9461059570313,
5.63574314117432,-54.9044151306152,
62.8437423706055,-50.3325691223145,
74.1372528076172,-34.8549728393555,
28.6584205627441,-1.61760354042053,
-18.3845329284668,14.5511941909790,
-20.1691875457764,-9.43072605133057,
10.8529710769653,-32.0917778015137,
34.9923286437988,-11.5462455749512,
41.7828140258789,30.5541343688965,
47.0096054077148,41.4956512451172,
52.3925399780273,19.2912464141846,
39.8505287170410,6.93319368362427,
6.39967536926270,25.4371833801270,
-18.3612766265869,45.1945343017578,
-13.9795722961426,41.1890144348145,
6.40037631988525,29.2362518310547,
9.62436771392822,28.0447559356689,
-14.4277315139771,18.8641681671143,
-38.2240829467773,-17.4932689666748,
-34.9659652709961,-45.6442337036133,
-11.1738281250000,-22.8616752624512,
8.60114002227783,31.6939735412598,
20.3194274902344,53.9165725708008,
33.7267112731934,20.4891242980957,
45.6342010498047,-17.8988151550293,
36.4678878784180,-15.5511741638184,
-0.130316078662872,7.96950626373291,
-29.8817386627197,4.52726745605469,
-21.1499977111816,-29.8227424621582,
16.3475608825684,-50.9610214233398,
33.2350311279297,-36.0474967956543,
5.12685489654541,-11.8938570022583,
-35.7230682373047,-11.7246913909912,
-44.6419944763184,-23.2224903106689,
-22.6915893554688,-15.3535614013672,
-10.2741470336914,12.7391881942749,
-30.6764354705811,25.7237205505371,
-59.1767616271973,0.845971584320068,
-53.8291320800781,-40.6475105285645,
-15.0719318389893,-58.0887298583984,
22.2360820770264,-33.9083061218262,
35.5487785339356,-0.724304437637329,
37.9243392944336,7.06042385101318,
38.0787353515625,-6.67158269882202,
25.1943721771240,-14.5874567031860,
-5.18689632415772,-2.93089866638184,
-29.1575756072998,8.45556640625000,
-16.0430850982666,-3.00000190734863,
18.0237083435059,-30.3310527801514,
21.2844333648682,-37.6061859130859,
-15.0923919677734,-12.5046606063843,
-39.1590385437012,18.1598358154297,
-9.31536674499512,19.3467540740967,
42.6386146545410,-0.989759802818298,
48.0780868530273,-7.59639310836792,
4.32852888107300,18.0909004211426,
-22.4555339813232,46.8366546630859,
7.18712997436523,36.9853057861328,
44.6276855468750,-6.77507352828980,
24.1895599365234,-41.0350303649902,
-40.8160095214844,-38.4444351196289,
-71.5218429565430,-20.1820793151855,
-33.7947540283203,-18.0286178588867,
21.4573001861572,-29.0057926177979,
26.1957702636719,-27.4854564666748,
-17.6203975677490,-8.45411109924316,
-51.5597915649414,7.59638786315918,
-41.1040344238281,11.7937135696411,
-8.30883598327637,22.0237598419189,
14.3150596618652,46.8577957153320,
20.0886936187744,65.9605712890625,
23.4603519439697,56.2561607360840,
31.0805644989014,28.6203231811523,
30.5970516204834,8.96274375915527,
13.1457386016846,2.94683933258057,
-10.0109939575195,-6.14551544189453,
-17.7904434204102,-17.5865688323975,
-2.71038007736206,-12.2381248474121,
21.4662761688232,7.56175422668457,
34.3477287292481,18.9894695281982,
24.1700630187988,8.47185039520264,
7.37035083770752,-4.58249664306641,
1.18102288246155,2.34270071983337,
2.31517720222473,20.8448963165283,
-6.98727798461914,26.1979904174805,
-31.8824558258057,17.3660240173340,
-51.4873962402344,16.2242050170898,
-37.6061820983887,27.3938751220703,
7.18006420135498,34.8510551452637,
46.9471855163574,28.3891754150391,
50.5359649658203,19.6275863647461,
20.2708263397217,11.3623971939087,
-11.2045392990112,-6.16536283493042,
-23.9269123077393,-33.3449401855469,
-25.9988040924072,-44.9888381958008,
-33.9395866394043,-23.3114967346191,
-45.1732215881348,14.1929807662964,
-41.7512588500977,32.8536224365234,
-16.8655662536621,22.9440155029297,
10.4925212860107,9.68505382537842,
16.4670028686523,9.60531711578369,
1.24145674705505,8.27474975585938,
-14.8648223876953,-4.88404273986816,
-14.3428754806519,-16.4400539398193,
-1.53213667869568,-13.2480325698853,
1.30388987064362,-1.38870692253113,
-11.4140958786011,1.07031726837158,
-31.1114234924316,-5.45830869674683,
-35.9478836059570,-8.96879196166992,
-17.0073471069336,-9.91090202331543,
10.3615875244141,-15.6035518646240,
17.7086467742920,-17.4731483459473,
-7.20518493652344,1.99658322334290,
-41.7249145507813,33.8804206848145,
-50.3891868591309,37.5749740600586,
-18.3065490722656,-5.72488927841187,
23.8234100341797,-58.2162246704102,
35.7924842834473,-66.6844940185547,
11.2722253799438,-31.3567848205566,
-14.2086629867554,-3.00894737243652,
-3.24986505508423,-16.7628002166748,
40.5595169067383,-45.7330093383789,
77.1322555541992,-44.0786514282227,
77.0926895141602,-4.64506101608276,
52.0356674194336,32.7553558349609,
31.8648052215576,37.4517860412598,
29.4923458099365,20.0620594024658,
31.2852153778076,12.1602287292480,
17.3513278961182,18.5780372619629,
-9.50166797637940,19.4742813110352,
-30.5522632598877,0.743518471717835,
-32.0790596008301,-23.4385795593262,
-16.9989318847656,-37.1450920104981,
-1.51627564430237,-40.3623008728027,
1.65163218975067,-45.1894836425781,
-7.47099685668945,-51.4257583618164,
-17.8434543609619,-36.5459823608398,
-17.5793228149414,0.0503435134887695,
-10.7891016006470,32.3195953369141,
-12.2180957794189,33.2802124023438,
-25.0797634124756,15.4003181457520,
-30.4042758941650,10.2302904129028,
-16.2082862854004,27.8152236938477,
7.64560651779175,46.1777954101563,
14.6353378295898,43.0116691589356,
1.44364380836487,32.0105743408203,
-6.26274013519287,36.6309700012207,
6.45724105834961,49.5266761779785,
23.6183452606201,40.9781761169434,
22.2251491546631,4.06560707092285,
3.88333845138550,-35.6536483764648,
-9.11639308929443,-53.1158638000488,
-6.90064859390259,-52.9704513549805,
-4.48378849029541,-53.2350769042969,
-14.0119628906250,-53.3800582885742,
-23.8142433166504,-30.6891403198242,
-19.5811252593994,10.0569076538086,
-6.30215978622437,27.4040298461914,
-1.10669672489166,-3.74717283248901,
-6.11189365386963,-53.9944877624512,
-5.55312871932983,-62.3625679016113,
12.2133903503418,-16.8428058624268,
32.9663314819336,25.7887630462647,
32.8409767150879,12.9743347167969,
12.6835613250732,-32.4791069030762,
0.992800712585449,-38.5080299377441,
14.3568143844605,14.2482976913452,
33.6963539123535,64.2746887207031,
25.9087009429932,49.4919013977051,
-5.76851320266724,-12.9529314041138,
-23.8956470489502,-46.0685272216797,
-4.80508708953857,-17.6760597229004,
29.1955509185791,34.8375091552734,
41.2413063049316,51.0299339294434,
28.5100498199463,23.9453716278076,
16.2471218109131,-12.7795066833496,
10.3555784225464,-29.7640991210938,
-2.07437920570374,-20.0542736053467,
-19.1716136932373,8.41076660156250,
-16.1005420684814,40.0563964843750,
12.7104883193970,55.4173812866211,
34.6972236633301,36.3066520690918,
25.4768619537354,-5.02766704559326,
5.90867948532105,-32.8490486145020,
10.8635931015015,-33.6194038391113,
31.7183780670166,-28.0776062011719,
31.2402305603027,-39.2487869262695,
6.56231594085693,-60.7296028137207,
-2.80842018127441,-59.4619483947754,
21.6208572387695,-18.2998466491699,
39.2657356262207,33.4958229064941,
10.0012207031250,52.4545707702637,
-40.7952995300293,27.4643135070801,
-61.4327583312988,-13.4084997177124,
-37.5085258483887,-29.9911308288574,
-5.54930400848389,-7.71170902252197,
4.37868595123291,26.9053249359131,
3.92845845222473,35.1259193420410,
9.84430313110352,6.12040805816650,
16.5476570129395,-30.5846252441406,
8.62344837188721,-34.9824333190918,
-7.74552297592163,-11.4734001159668,
-18.9178504943848,5.89418888092041,
-25.8658866882324,-4.92206764221191,
-31.3086051940918,-24.9178466796875,
-20.0044364929199,-26.2983169555664,
18.2037601470947,-9.51138210296631,
59.5721817016602,-5.61678504943848,
61.6428756713867,-20.2480010986328,
24.7310619354248,-29.0244331359863,
-9.14964580535889,-19.0361442565918,
-3.94737696647644,-0.766021966934204,
27.6615161895752,8.60854339599609,
44.1404991149902,8.61527442932129,
36.8482589721680,5.07260990142822,
27.8047409057617,-10.2849264144897,
26.3037128448486,-40.6870918273926,
18.9486713409424,-55.9412117004395,
-0.801955580711365,-29.4143714904785,
-20.6554889678955,16.3595409393311,
-24.1623802185059,24.7960796356201,
-6.51047277450562,-19.1923732757568,
27.3792648315430,-60.9523010253906,
61.2082252502441,-43.3050460815430,
68.7754669189453,12.7011423110962,
32.2910270690918,37.7397270202637,
-22.3178787231445,6.10949230194092,
-44.5475654602051,-31.5092887878418,
-11.4111700057983,-23.0641994476318,
30.5917854309082,17.1348361968994,
25.3249511718750,31.2772388458252,
-16.6825447082520,-0.958197355270386,
-34.8920249938965,-36.2262191772461,
-8.21282958984375,-29.8473167419434,
21.9311504364014,8.48420333862305,
21.1393203735352,29.8776130676270,
9.18999481201172,14.1702604293823,
22.1876220703125,-15.3336992263794,
51.4089279174805,-27.4382572174072,
58.0584869384766,-15.8736066818237,
38.2717285156250,-0.301290333271027,
27.4823398590088,-1.04050707817078,
37.0617752075195,-12.3931169509888,
38.2038230895996,-24.9279747009277,
9.81697654724121,-36.5765151977539,
-22.8060054779053,-47.4737815856934,
-26.4043045043945,-50.5720558166504,
-11.4165058135986,-39.4199180603027,
-2.02321219444275,-16.3101272583008,
1.93235135078430,0.150493264198303,
17.3803424835205,-6.26731491088867,
37.2051963806152,-25.7584114074707,
34.9038734436035,-23.2966976165772,
8.40686702728272,8.78790855407715,
-8.73587894439697,37.1201477050781,
0.724299550056458,21.0818157196045,
12.4628162384033,-28.9429626464844,
-1.12902796268463,-62.4848518371582,
-24.6674365997314,-49.8107833862305,
-29.6537609100342,-20.6367340087891,
-18.9863452911377,-18.3255348205566,
-16.4144935607910,-36.5566024780273,
-19.7677783966064,-40.2290573120117,
-3.35780310630798,-17.6381473541260,
35.6959991455078,1.83611273765564,
60.2421531677246,7.29260063171387,
41.0492553710938,18.1967544555664,
-0.136657238006592,47.8704490661621,
-18.1866397857666,67.9872360229492,
-2.86127424240112,48.7730789184570,
16.2237358093262,13.1778907775879,
14.7106504440308,9.24495506286621,
0.770533859729767,46.2472496032715,
-11.2377538681030,73.6360549926758,
-20.4823894500732,49.0396003723145,
-28.3246517181397,-12.8227024078369,
-31.7377395629883,-58.4127807617188,
-29.6874599456787,-59.6965408325195,
-22.8508968353272,-28.3440971374512,
-18.3888645172119,11.2441768646240,
-17.8661289215088,41.8795433044434,
-19.9209842681885,49.6827278137207,
-23.4390525817871,35.5090141296387,
-25.0530872344971,12.0981445312500,
-14.6105651855469,-5.24563884735107,
2.21139049530029,-14.8168783187866,
1.28891348838806,-29.8210926055908,
-25.8225097656250,-53.4353637695313,
-42.4242782592773,-70.8812789916992,
-14.4671764373779,-67.7379608154297,
35.3955268859863,-46.1124343872070,
40.7810134887695,-16.6697311401367,
-16.4029064178467,17.5979843139648,
-69.9901733398438,43.0095367431641,
-54.8253364562988,36.0073585510254,
6.29648494720459,-3.35054445266724,
30.6708850860596,-40.8085975646973,
-6.75406789779663,-33.6882476806641,
-40.7789192199707,10.3163824081421,
-13.3134756088257,35.3529891967773,
48.1557846069336,11.6185626983643,
77.5176239013672,-26.3977279663086,
59.6809310913086,-24.5649375915527,
37.1205024719238,16.6205749511719,
39.4882621765137,48.3900909423828,
50.5278015136719,41.1157989501953,
46.6289634704590,17.7634925842285,
26.1406021118164,8.82380485534668,
4.62872695922852,8.74864292144775,
-11.9416341781616,-7.21244955062866,
-17.4541378021240,-34.4810600280762,
-1.33067536354065,-42.2226943969727,
32.3784561157227,-15.6869239807129,
47.5196609497070,24.2559757232666,
22.9858779907227,45.7568016052246,
-17.6621398925781,43.4813880920410,
-34.4844284057617,36.4464187622070,
-24.3419952392578,32.5627861022949,
-12.3315277099609,25.1463680267334,
-13.0742874145508,7.62074756622314,
-16.1198348999023,-15.0771045684814,
-11.0318708419800,-25.3523597717285,
-15.7879772186279,-12.2683134078980,
-40.3365631103516,16.4753265380859,
-61.7854652404785,30.5980491638184,
-55.0662193298340,10.9095115661621,
-29.5310001373291,-25.9240322113037,
-15.6455554962158,-42.2011070251465,
-19.5188159942627,-18.2157688140869,
-25.4647884368897,19.0158939361572,
-28.2169609069824,20.3910446166992,
-36.1774482727051,-19.3028888702393,
-44.3525962829590,-57.8954277038574,
-33.6830978393555,-60.2372474670410,
-3.29075336456299,-34.2666740417481,
16.2461910247803,-16.7060394287109,
0.490114212036133,-21.3625946044922,
-24.9913730621338,-38.4679794311523,
-18.4533443450928,-54.0228500366211,
18.8980827331543,-57.9728736877441,
45.2722358703613,-41.1260871887207,
42.8546485900879,2.15659928321838,
35.3842658996582,50.0491828918457,
39.6228485107422,61.6970787048340,
39.1609725952148,22.0326633453369,
11.5185661315918,-32.2017517089844,
-24.6978473663330,-49.9314460754395,
-35.3302497863770,-28.5760002136230,
-16.5351047515869,1.45897781848907,
1.02726721763611,14.8419780731201,
1.47400641441345,6.39014959335327,
-0.254448711872101,-19.1248531341553,
7.74525547027588,-44.7762298583984,
9.71667385101318,-45.5458183288574,
-1.13890480995178,-3.61829900741577,
-4.78129529953003,49.2676887512207,
11.1833715438843,58.3370208740234,
25.0001621246338,12.0186548233032,
13.2872085571289,-26.0995693206787,
-12.5320873260498,-9.12909412384033,
-27.4631309509277,25.9214286804199,
-27.6975383758545,5.56533670425415,
-29.7013549804688,-62.9939460754395,
-29.4173316955566,-96.4056091308594,
-4.52804565429688,-47.9853668212891,
34.4135742187500,26.2566871643066,
37.6306610107422,40.6296424865723,
-2.22914195060730,-6.42261266708374,
-30.2710838317871,-44.0661430358887,
-3.23988842964172,-30.3197708129883,
41.7923049926758,6.67577981948853,
45.9443244934082,30.2893962860107,
10.8071517944336,40.3037490844727,
-8.58207130432129,51.6556930541992,
2.86097383499146,51.8488273620606,
2.87284541130066,28.4109039306641,
-28.2467155456543,2.28092527389526,
-47.2991142272949,2.41862487792969,
-18.5287036895752,25.6049365997314,
15.2821340560913,39.9035072326660,
0.240380167961121,24.4496135711670,
-48.5245704650879,-6.46821975708008,
-66.9768295288086,-20.0895195007324,
-42.7108078002930,-15.4146842956543,
-28.0240345001221,-8.75091743469238,
-43.0703544616699,-14.8714265823364,
-46.6391754150391,-39.9987525939941,
-1.27107143402100,-69.8827743530273,
57.6161460876465,-71.5267257690430,
69.1477050781250,-23.1278228759766,
31.0553436279297,44.5792541503906,
0.816772460937500,71.3052978515625,
4.57671451568604,30.4876384735107,
10.6617355346680,-23.5641098022461,
-12.0515556335449,-27.8375453948975,
-46.5178451538086,13.4024343490601,
-58.2287445068359,28.8436203002930,
-38.9621849060059,-18.7576694488525,
-4.37062168121338,-79.4812850952148,
32.0688095092773,-82.8989715576172,
59.4924125671387,-24.7900543212891,
71.3248672485352,35.5709915161133,
59.3390846252441,57.1224441528320,
31.8707256317139,52.0130538940430,
5.48206233978272,49.3482398986816,
-14.0882759094238,50.7639732360840,
-33.4975776672363,36.6612701416016,
-50.1380043029785,4.40032863616943,
-45.8538665771484,-30.0537929534912,
-23.9899597167969,-51.4555206298828,
-3.11736869812012,-57.1084938049316,
7.48657369613648,-51.9375152587891,
12.6564445495605,-39.8159942626953,
12.3049087524414,-23.8517894744873,
-4.87567329406738,-8.25578689575195,
-37.7632789611816,10.4044532775879,
-55.1888313293457,33.6162948608398,
-32.9572029113770,49.2328872680664,
10.1615562438965,46.1076202392578,
32.8141250610352,28.4672775268555,
23.5791873931885,15.9365520477295,
13.3890380859375,20.5956878662109,
12.1804943084717,27.8947486877441,
-2.40287971496582,17.3947048187256,
-36.1151390075684,-7.85482597351074,
-53.7822456359863,-18.4836254119873,
-22.2571086883545,0.621108770370483,
27.5467720031738,31.1792907714844,
41.1063270568848,44.3977012634277,
12.8081455230713,29.8746604919434,
-11.1561679840088,8.33562088012695,
-6.05425691604614,-0.445536792278290,
-2.19177842140198,9.11081695556641,
-26.4648513793945,23.6282424926758,
-48.0320014953613,26.0061473846436,
-25.1021347045898,7.80186939239502,
23.2349395751953,-23.4012527465820,
38.7210159301758,-47.8457794189453,
12.3314666748047,-46.7223815917969,
-10.3448266983032,-25.3159465789795,
4.71739816665649,-4.24211263656616,
38.0926551818848,1.59834313392639,
51.0035629272461,-0.418034881353378,
36.3329696655273,2.43386578559876,
12.0172729492188,11.1467514038086,
-9.98747920989990,17.7107563018799,
-24.3958511352539,20.9905281066895,
-18.0187377929688,26.8026103973389,
12.3532886505127,32.4006805419922,
41.3945693969727,20.4668159484863,
40.8910865783691,-11.9267454147339,
26.7482109069824,-38.3937988281250,
32.4397087097168,-34.4071884155273,
50.7358932495117,-2.27395915985107,
39.4813880920410,24.7487220764160,
-11.4318675994873,22.6768379211426,
-53.4446372985840,5.13333511352539,
-38.2279243469238,-5.52309417724609,
15.3233270645142,-9.23849964141846,
42.3889999389648,-20.4419231414795,
17.6192607879639,-34.8629074096680,
-18.7768707275391,-30.2750530242920,
-24.0165252685547,-0.782006502151489,
2.90017676353455,21.5902671813965,
33.3141593933106,8.94479084014893,
48.3989715576172,-17.4382190704346,
48.9895172119141,-9.57993412017822,
38.8800277709961,39.1138877868652,
23.3915157318115,76.8797225952148,
9.86297225952148,56.1526908874512,
2.78749728202820,-2.76536059379578,
-3.39124584197998,-30.0905475616455,
-15.9760389328003,3.33976030349731,
-32.9456253051758,46.5986938476563,
-39.4294738769531,32.2046089172363,
-30.5084018707275,-35.4303894042969,
-20.6252689361572,-84.7573623657227,
-19.1040401458740,-63.9408226013184,
-18.0813980102539,0.0188597440719605,
-7.74155521392822,39.1817474365234,
6.25074434280396,26.5608177185059,
11.8366537094116,3.16134834289551,
3.20024991035461,10.4369020462036,
-8.32641410827637,32.4205818176270,
-16.9277935028076,31.2912845611572,
-25.4025764465332,7.93504953384399,
-32.0112762451172,-6.30435657501221,
-24.8527412414551,-0.325120627880096,
1.24185776710510,-5.39094161987305,
27.4032707214355,-34.9664726257324,
30.2331752777100,-51.0162811279297,
9.15121841430664,-17.1200218200684,
-14.8008975982666,34.4150276184082,
-28.1404170989990,43.1023674011231,
-31.5369911193848,4.55740404129028,
-28.5731372833252,-26.8737964630127,
-11.4849796295166,-13.1674385070801,
20.8913230895996,10.1691465377808,
54.1016731262207,-1.40648031234741,
67.2260742187500,-29.9380683898926,
60.7971496582031,-26.4704246520996,
45.7770919799805,10.9814777374268,
27.0773906707764,33.6432876586914,
2.26094722747803,16.5107898712158,
-20.1177864074707,-7.67803812026978,
-21.7806282043457,4.32547473907471,
-3.93094754219055,38.2342643737793,
12.4447307586670,48.3321495056152,
10.0593442916870,15.9161930084229,
-4.39544248580933,-25.1684703826904,
-14.6020565032959,-39.7215538024902,
-16.5843944549561,-30.1639938354492,
-16.7414360046387,-15.6664676666260,
-10.0324764251709,-10.4923801422119,
11.3133563995361,-9.76943492889404,
41.5037727355957,-1.28420066833496,
58.3418502807617,13.1665353775024,
50.5330047607422,21.8842067718506,
32.8397979736328,16.4102897644043,
16.5833950042725,-3.80843496322632,
1.21285116672516,-29.2218227386475,
-16.8214225769043,-47.6674118041992,
-30.2661666870117,-55.2840003967285,
-33.9450111389160,-53.7597427368164,
-29.2725028991699,-37.7188415527344,
-23.1826190948486,-0.340378463268280,
-16.9773349761963,46.0431175231934,
-8.00919246673584,68.2169265747070,
-6.82529449462891,43.2454299926758,
-22.7945289611816,-9.77576637268066,
-41.5109825134277,-39.7636489868164,
-39.5148124694824,-21.9227466583252,
-22.2644901275635,11.0835075378418,
-16.0475063323975,11.3321132659912,
-25.5070896148682,-25.0629425048828,
-17.9035186767578,-50.9990081787109,
15.8212633132935,-30.8807468414307,
39.1800765991211,13.7678527832031,
13.6351661682129,33.0321044921875,
-34.9542617797852,9.21339035034180,
-42.6769218444824,-25.7942790985107,
4.22804927825928,-34.2306442260742,
46.9338111877441,-20.5896472930908,
38.3442306518555,-8.99856758117676,
6.53825283050537,-4.84911155700684,
5.17254877090454,6.21905565261841,
33.5698852539063,33.4619941711426,
46.9981803894043,54.6569252014160,
26.3939228057861,45.6756477355957,
-3.77441835403442,12.3117532730103,
-21.1723155975342,-19.7940082550049,
-31.2720260620117,-28.2858047485352,
-40.5087623596191,-10.8274478912354,
-33.8340911865234,18.9510269165039,
-4.59469079971314,39.4588546752930,
21.8313350677490,39.3526840209961,
20.9156436920166,15.4703960418701,
9.56412506103516,-14.0440835952759,
18.0715274810791,-21.8221282958984,
35.4496803283691,-1.67031359672546,
27.7528953552246,28.7789726257324,
1.14215040206909,38.6331787109375,
-4.12514495849609,16.8695640563965,
28.1052589416504,-18.4522247314453,
61.5406112670898,-33.4191589355469,
58.5634498596191,-9.91603279113770,
28.0234031677246,26.6105613708496,
7.44507503509522,41.4215202331543,
1.70407116413116,28.4708728790283,
-10.4012498855591,20.6984844207764,
-22.8663520812988,42.4579391479492,
-12.4025039672852,68.0327911376953,
17.3667240142822,52.2420196533203,
27.8442726135254,-3.34520626068115,
10.0611782073975,-48.5827560424805,
-0.933389663696289,-47.9422912597656,
13.9673032760620,-28.8705406188965,
27.8318881988525,-28.6731986999512,
11.0042896270752,-33.2692909240723,
-17.3614234924316,-8.55817031860352,
-13.0720729827881,39.9775886535645,
20.5031013488770,62.5427513122559,
36.6811637878418,39.9686470031738,
21.0762710571289,7.43271493911743,
10.4752130508423,-0.293356001377106,
25.8336944580078,6.52853965759277,
39.5976943969727,0.0480237007141113,
29.9665203094482,-16.3014640808105,
16.8741416931152,-18.1880779266357,
27.3399600982666,-10.6915683746338,
35.9576873779297,-12.4569578170776,
2.63809728622437,-20.9263248443604,
-51.6481666564941,-7.44185256958008,
-59.4734344482422,26.1464309692383,
-5.17165184020996,47.2962799072266,
44.5451812744141,40.2025947570801,
27.1844234466553,31.9359989166260,
-33.9641532897949,41.4437103271484,
-68.2128372192383,45.3684272766113,
-54.9666671752930,13.8124885559082,
-37.5121078491211,-39.5787925720215,
-39.7937316894531,-62.7246932983398,
-29.9943332672119,-40.5272445678711,
21.2557659149170,-11.4942979812622,
78.7245483398438,-14.3369703292847,
82.3864669799805,-37.8824577331543,
25.7762718200684,-48.1144638061523,
-24.6564216613770,-32.5129508972168,
-14.4036302566528,-6.08218097686768,
28.3639736175537,10.2761011123657,
35.6815376281738,9.08640575408936,
-5.46484947204590,-6.84578609466553,
-40.7478103637695,-20.1507663726807,
-21.7778244018555,-16.0206165313721,
27.8709163665772,6.61111545562744,
45.2230873107910,27.7293930053711,
10.7332000732422,30.6286563873291,
-26.2037715911865,21.1483993530273,
-25.2068519592285,20.5324783325195,
-3.59225273132324,30.6374244689941,
-5.90117454528809,26.7539443969727,
-32.6337394714356,3.61695575714111,
-42.1276588439941,-18.3074207305908,
-8.51496696472168,-19.3726215362549,
39.3894119262695,-3.98664426803589,
52.4158592224121,11.1071472167969,
22.9251251220703,20.1636676788330,
-10.7871198654175,28.3506450653076,
-18.6874561309814,29.3004665374756,
-11.2651195526123,12.0750646591187,
-14.6596946716309,-10.8385782241821,
-31.3224258422852,-14.7376585006714,
-37.3165245056152,2.40691614151001,
-15.0686197280884,9.45102119445801,
13.1521835327148,-16.5320377349854,
17.7266273498535,-49.9059906005859,
-1.80292773246765,-52.4044494628906,
-15.7260475158691,-26.6514282226563,
-1.05115032196045,-12.4105882644653,
32.3393783569336,-26.6848373413086,
56.7911300659180,-46.7760658264160,
58.5444793701172,-39.8234634399414,
43.1875534057617,-11.1121425628662,
18.5084857940674,5.76465129852295,
-9.93045234680176,-3.75522637367249,
-26.2137088775635,-23.0977916717529,
-13.8123416900635,-34.3059997558594,
24.8054008483887,-26.9530506134033,
56.1457595825195,-0.630964994430542,
55.7013282775879,27.3419170379639,
31.9021263122559,26.6712856292725,
15.4230928421021,-5.30381298065186,
16.8742580413818,-28.0187091827393,
23.6964988708496,-3.12904882431030,
22.0462646484375,43.0871734619141,
9.78448009490967,43.6517524719238,
-7.99916505813599,-19.3445339202881,
-26.8442382812500,-70.4031829833984,
-34.8993949890137,-44.4499511718750,
-19.4241733551025,18.2175292968750,
12.1168212890625,25.2000236511230,
22.8125381469727,-30.0954971313477,
-8.16590499877930,-58.5195808410645,
-52.8485870361328,-15.0317935943604,
-65.8018035888672,35.3612442016602,
-38.9369201660156,16.2977008819580,
-12.2297677993774,-42.4445381164551,
-15.1335744857788,-52.1121864318848,
-29.8925590515137,0.858051657676697,
-20.6695728302002,38.7011756896973,
14.9136810302734,8.38681983947754,
47.0090446472168,-44.3719329833984,
55.5769157409668,-49.2633857727051,
50.1111335754395,-7.84874343872070,
44.6597480773926,23.5590877532959,
35.8775215148926,16.8512744903564,
16.8186511993408,-11.7494859695435,
0.0498152077198029,-39.7848930358887,
4.94429588317871,-56.4816017150879,
28.1521854400635,-50.7112007141113,
44.5872116088867,-21.8496665954590,
33.1723442077637,7.15978622436523,
-2.28032445907593,7.85859966278076,
-35.0298843383789,-13.0221138000488,
-39.6571426391602,-16.9597129821777,
-21.0779571533203,13.6808013916016,
-6.34887123107910,37.6575736999512,
-13.0888872146606,18.3599777221680,
-28.5791110992432,-20.0170593261719,
-23.6331596374512,-22.2285804748535,
4.94079065322876,19.6027221679688,
21.6355304718018,61.7429924011231,
0.926434993743897,60.0115661621094,
-33.3338584899902,17.8363857269287,
-33.4809570312500,-24.7077350616455,
0.137058734893799,-42.5538597106934,
21.8289051055908,-37.4185867309570,
6.27988958358765,-22.7796440124512,
-15.1798458099365,-15.2910623550415,
-2.27505850791931,-25.0276908874512,
32.2949600219727,-46.1289901733398,
40.7471771240234,-53.1620025634766,
15.2974672317505,-35.3792953491211,
-8.17600917816162,-19.8600215911865,
-10.4902296066284,-32.1803321838379,
-13.6600685119629,-54.0612258911133,
-34.1860771179199,-43.3450851440430,
-41.7013893127441,4.28523969650269,
-4.88159561157227,42.1728515625000,
44.9459571838379,31.4142208099365,
50.6006584167481,-7.58410453796387,
8.73529815673828,-23.9245128631592,
-25.3753890991211,-14.3531513214111,
-11.7255725860596,-11.5078010559082,
25.9087066650391,-21.5128707885742,
37.7592010498047,-17.9495868682861,
15.6777572631836,8.74792671203613,
-8.88826656341553,20.7735519409180,
-10.1458377838135,-6.06815338134766,
10.2790546417236,-39.9344329833984,
40.4363594055176,-40.1516036987305,
58.5505409240723,-12.7345256805420,
42.0570945739746,-0.482488334178925,
-8.73919486999512,-12.1578769683838,
-50.6254081726074,-12.5440607070923,
-38.9386177062988,16.8341884613037,
12.8939180374146,44.9654922485352,
47.2285041809082,36.7652854919434,
31.2012481689453,9.20602512359619,
-3.07567858695984,-2.90338921546936,
-5.10675811767578,6.81636238098145,
23.9954586029053,22.9506874084473,
39.2880821228027,32.4177818298340,
23.1922492980957,33.6091308593750,
3.75617551803589,18.9944229125977,
3.51023507118225,-15.2725114822388,
18.0635757446289,-44.0032997131348,
31.6786537170410,-38.1625976562500,
40.3474044799805,1.86772251129150,
46.1236877441406,35.0877761840820,
36.6875648498535,39.9720611572266,
5.98718643188477,38.5487632751465,
-27.0351142883301,49.9570312500000,
-41.3966598510742,52.1247673034668,
-34.6471519470215,22.9931354522705,
-23.8079586029053,-11.2510643005371,
-12.7277803421021,-10.2221717834473,
10.5232982635498,26.2145538330078,
35.3987045288086,50.5627250671387,
29.5283756256104,33.4475250244141,
-14.1990299224854,-6.31130456924439,
-53.4882202148438,-36.6332855224609,
-47.2735061645508,-56.0564765930176,
-2.77478408813477,-69.4800262451172,
30.5839748382568,-61.6813316345215,
22.0963516235352,-21.2475624084473,
-12.0566539764404,15.2647647857666,
-41.0318298339844,9.67672729492188,
-51.8055458068848,-19.4859237670898,
-45.6544151306152,-21.3723678588867,
-23.7831192016602,15.7572040557861,
-1.75053322315216,48.9670906066895,
-6.88713264465332,47.7723922729492,
-41.3875579833984,27.5836544036865,
-70.4250183105469,16.5931415557861,
-59.6748237609863,4.00591087341309,
-26.0978374481201,-24.5375785827637,
-13.5674943923950,-40.1223678588867,
-30.0405445098877,-11.2858028411865,
-40.9323272705078,26.9780635833740,
-22.9195652008057,11.8937263488770,
-2.31270670890808,-46.0125122070313,
-12.0491170883179,-68.0102233886719,
-35.0706672668457,-25.8211765289307,
-28.1859493255615,15.3076601028442,
9.01795959472656,-4.60728263854981,
37.4968223571777,-46.2053260803223,
31.4901256561279,-28.4284629821777,
6.04273700714111,46.5816192626953,
-13.1343250274658,90.9327239990234,
-18.1244697570801,59.0662040710449,
-13.1306991577148,9.01537322998047,
1.90001857280731,1.09723627567291,
17.3015003204346,22.8814315795898,
15.6590967178345,29.5372524261475,
-9.45149993896484,16.7723560333252,
-32.1828384399414,8.85542106628418,
-31.0725784301758,2.29284787178040,
-24.3067741394043,-21.4738616943359,
-40.5798568725586,-42.0175743103027,
-60.7788200378418,-26.0547046661377,
-39.2419319152832,13.5125379562378,
20.0816402435303,22.1133804321289,
60.6049270629883,-13.9550447463989,
42.8284988403320,-35.4451942443848,
-5.31598806381226,-1.35102653503418,
-26.0088253021240,38.8431510925293,
-9.08430290222168,13.8734989166260,
12.9256067276001,-55.2294692993164,
18.0991954803467,-84.3426666259766,
13.7933368682861,-35.5684356689453,
7.40962409973145,29.3004608154297,
-7.10930633544922,34.4546394348145,
-20.6728935241699,-17.7739276885986,
-13.0846242904663,-55.8803291320801,
8.00645637512207,-42.6279830932617,
7.12667179107666,0.0320479869842529,
-23.3238525390625,32.1701889038086,
-45.1895141601563,40.6788520812988,
-27.5190620422363,35.4311370849609,
11.9496879577637,24.0574417114258,
34.0258979797363,13.4000921249390,
30.4561786651611,14.2195167541504,
29.2155399322510,27.4702033996582,
30.4584140777588,31.6607341766357,
9.94342041015625,7.69042158126831,
-27.0716419219971,-33.5387573242188,
-39.6579551696777,-59.3429870605469,
-10.2658920288086,-54.7234001159668,
21.6095695495605,-48.3421821594238,
17.0307235717773,-66.4478836059570,
-6.74138689041138,-89.1941146850586,
-10.7133407592773,-71.9739379882813,
6.54172182083130,-12.7833328247070,
9.59073638916016,35.7259635925293,
-11.0738668441772,27.6072216033936,
-19.0871028900147,-10.8313159942627,
13.1522617340088,-18.2177066802979,
59.0961151123047,22.6244201660156,
71.3583602905273,55.0447311401367,
40.3956260681152,33.2096099853516,
-4.31248903274536,-16.0871658325195,
-27.3377189636230,-29.6834812164307,
-17.8982219696045,3.92464542388916,
15.1445426940918,36.5510482788086,
47.6552581787109,29.5579452514648,
48.2204093933106,3.38900828361511,
6.40236949920654,3.86802673339844,
-47.5972862243652,29.5285358428955,
-67.7985458374023,40.2756881713867,
-34.9066886901856,13.1119804382324,
18.3194541931152,-19.4686622619629,
42.0366973876953,-16.1911849975586,
24.7526626586914,23.6488437652588,
-2.46734213829041,58.5079154968262,
-6.21149826049805,54.3989067077637,
10.2803144454956,21.5807075500488,
23.5908451080322,-3.04898953437805,
15.6750001907349,-1.82758998870850,
-1.00431656837463,11.7422981262207,
-8.30980014801025,17.7288322448730,
-5.48044204711914,11.8712415695190,
-9.39488124847412,5.82102537155151,
-28.8994712829590,7.78515768051148,
-53.1598587036133,10.7643384933472,
-58.8742599487305,7.68751859664917,
-42.3047561645508,-1.03173482418060,
-14.9753026962280,-9.89824485778809,
8.91843032836914,-14.1451568603516,
24.6954574584961,-7.63028335571289,
34.9147186279297,9.41428661346436,
40.1426200866699,25.0850658416748,
36.0874061584473,23.7368202209473,
25.7911281585693,-1.87842965126038,
17.5931053161621,-31.2918300628662,
19.5531616210938,-37.5227432250977,
30.4893112182617,-17.9064350128174,
38.6167068481445,7.20424079895020,
31.7739353179932,16.4581336975098,
9.49162769317627,7.36916875839233,
-17.3247985839844,-6.32010650634766,
-35.6811828613281,-10.5069665908813,
-42.0690841674805,-4.20181274414063,
-41.7025299072266,5.28261804580689,
-41.7838897705078,7.68913269042969,
-40.3197059631348,-0.435179769992828,
-36.4907684326172,-7.42076826095581,
-31.2575950622559,0.410746276378632,
-28.5222377777100,19.5832939147949,
-26.8020687103272,22.8106746673584,
-22.3498744964600,-4.54003334045410,
-13.1502590179443,-39.4031715393066,
-8.76265525817871,-44.1469688415527,
-9.85632324218750,-17.4588527679443,
-10.3871965408325,3.57942819595337,
-2.73534345626831,-12.6114130020142,
8.24470901489258,-47.0161361694336,
10.4463872909546,-56.2669296264648,
-5.41236686706543,-26.5254173278809,
-30.9609355926514,9.68486976623535,
-41.5873603820801,22.3451690673828,
-25.9538345336914,9.08341026306152,
5.74049949645996,-12.8266506195068,
25.0691623687744,-35.0005035400391,
22.3159580230713,-50.9421310424805,
15.4091567993164,-48.8926811218262,
34.7945327758789,-26.5111732482910,
71.6114349365234,-3.47027301788330,
82.6348648071289,-0.504463195800781,
48.3008880615234,-13.5757503509521,
1.71756553649902,-22.3682880401611,
-11.6495895385742,-21.5946712493897,
4.15705299377441,-30.8546752929688,
6.83401584625244,-55.4151268005371,
-18.8377227783203,-64.3515090942383,
-36.3777809143066,-32.0057716369629,
-14.7352972030640,21.1567516326904,
19.5102958679199,58.7019805908203,
23.3269081115723,66.3923645019531,
4.85175037384033,53.6340713500977,
11.2181921005249,30.5274848937988,
47.6436462402344,2.69943928718567,
65.8027267456055,-14.2227602005005,
32.3844642639160,-3.59997415542603,
-18.4840240478516,19.7445793151855,
-32.9704055786133,18.5033264160156,
-12.3018760681152,-7.96320438385010,
3.47374057769775,-14.7364635467529,
-4.28678226470947,18.7318134307861,
-12.7922668457031,47.9715270996094,
-4.01890182495117,28.2993125915527,
9.88625335693359,-15.8301334381104,
18.6475963592529,-23.0787220001221,
30.6148834228516,6.12328624725342,
46.9019355773926,20.7745666503906,
39.4059410095215,-2.21242523193359,
-7.80938720703125,-19.1070632934570,
-57.7342491149902,4.19428539276123,
-61.1779251098633,27.6667289733887,
-19.4004344940186,1.72600698471069,
15.9335269927979,-50.9697227478027,
10.4783210754395,-61.1408996582031,
-14.6757450103760,-16.9356861114502,
-20.1318073272705,22.9618568420410,
-2.20725727081299,19.3982563018799,
10.3660764694214,-2.54444408416748,
-0.783291935920715,-6.24755144119263,
-21.9510898590088,-5.58559226989746,
-33.4713249206543,-29.6142635345459,
-20.6572132110596,-66.7762680053711,
16.0382690429688,-72.4759674072266,
57.4635276794434,-30.5612659454346,
77.3539123535156,21.9949607849121,
59.4157333374023,45.6334190368652,
20.3977642059326,38.3533096313477,
-6.04178190231323,20.3455410003662,
-3.67062854766846,-0.135277926921844,
18.8588027954102,-18.7750892639160,
38.6013793945313,-24.4190731048584,
47.0950736999512,-9.36904335021973,
40.8429298400879,16.5115470886230,
10.4140567779541,35.7670249938965,
-37.7136688232422,37.5151214599609,
-73.6961975097656,22.7377834320068,
-67.6343154907227,1.22514367103577,
-23.1139755249023,-16.9686508178711,
22.1121387481689,-25.6020240783691,
39.0666427612305,-20.3512020111084,
34.4841079711914,-7.32359790802002,
31.0219383239746,1.32976257801056,
32.3151245117188,9.24275016784668,
32.4722862243652,23.6620998382568,
27.3823394775391,36.5396347045898,
29.4516696929932,34.3373107910156,
36.8878784179688,15.4742221832275,
31.1353797912598,0.553290307521820,
3.64530086517334,-2.03751349449158,
-26.9089298248291,-9.73085689544678,
-35.3957939147949,-32.4154510498047,
-14.5038690567017,-47.5074157714844,
15.8062515258789,-19.0352554321289,
33.5294952392578,42.4115142822266,
32.0007743835449,80.1508941650391,
23.0274829864502,58.5633850097656,
21.3846111297607,9.96499824523926,
31.7282848358154,-14.2892904281616,
42.4608230590820,-6.97683620452881,
33.1654281616211,1.16061341762543,
1.21761488914490,-9.13475990295410,
-31.3324127197266,-25.1992683410645,
-31.5069274902344,-29.6259899139404,
-3.93533229827881,-29.8337688446045,
15.8333225250244,-26.5931911468506,
5.80408382415772,-6.53838109970093,
-16.8276023864746,27.9625911712647,
-22.4296493530273,43.4602851867676,
-1.78519296646118,16.4368019104004,
26.1955814361572,-22.6248264312744,
39.5278930664063,-16.1982154846191,
32.6858863830566,36.5314407348633,
7.13051605224609,66.3901672363281,
-24.1237716674805,32.2408866882324,
-29.8689136505127,-25.5025234222412,
6.42989540100098,-30.9292030334473,
50.3685684204102,19.6301517486572,
48.7985649108887,52.5240821838379,
-1.61370968818665,16.3391799926758,
-36.1376838684082,-47.9402313232422,
-7.18429899215698,-58.8808441162109,
45.2646980285645,-5.40436983108521,
44.5754470825195,48.8418884277344,
-9.17274093627930,43.3864173889160,
-39.6606178283691,-4.98212718963623,
0.0876245498657227,-33.1579742431641,
56.6599617004395,-12.5461044311523,
45.9928703308106,29.6268501281738,
-25.5062961578369,47.9311637878418,
-76.3175125122070,37.6793327331543,
-54.2924270629883,28.4911079406738,
0.508056402206421,30.8338165283203,
21.0155906677246,29.4499149322510,
3.44822883605957,8.67201614379883,
-4.87883949279785,-21.8813037872314,
18.2284431457520,-28.3293018341064,
40.7599372863770,2.44142532348633,
21.1811332702637,42.5604324340820,
-32.8175659179688,56.1590843200684,
-70.6364746093750,39.5411415100098,
-60.9408454895020,11.3110218048096,
-20.8892631530762,-11.9800262451172,
16.0286560058594,-30.0288486480713,
33.4143562316895,-43.6895561218262,
35.9248657226563,-34.4604110717773,
32.6826438903809,4.73698186874390,
21.4149398803711,44.1577415466309,
-0.700560808181763,42.8847579956055,
-17.7550849914551,-6.72160148620606,
-18.4768791198730,-58.6647682189941,
-8.30236721038818,-67.8512878417969,
0.0636719912290573,-36.5347023010254,
1.85095024108887,-4.63529586791992,
5.74724483489990,1.40565013885498,
16.7738475799561,-3.43339896202087,
25.6857395172119,4.05131673812866,
19.6631946563721,23.0603275299072,
2.84697175025940,30.9206905364990,
-7.94540977478027,10.7757797241211,
-7.76995468139648,-24.9090747833252,
-6.25927209854126,-47.2023086547852,
-16.9344062805176,-39.2774353027344,
-36.1432418823242,-5.28990888595581,
-43.5360832214356,29.4792366027832,
-25.2915897369385,39.9549674987793,
7.79427337646484,20.5464401245117,
30.2063255310059,-9.19185352325440,
26.5835475921631,-27.6122035980225,
6.41029071807861,-30.1282863616943,
-11.1857357025146,-28.1180210113525,
-17.3083839416504,-31.1160087585449,
-15.7949686050415,-34.5337677001953,
-13.3459920883179,-28.7301025390625,
-10.0922861099243,-14.6476469039917,
-8.18218994140625,-0.0598560571670532,
-8.83671188354492,14.2009105682373,
-9.93832492828369,31.7631206512451,
-8.11648464202881,41.5955543518066,
-3.05302548408508,28.2068424224854,
-1.87503004074097,-6.37334108352661,
-3.12170147895813,-34.9992713928223,
1.04881632328033,-28.5181846618652,
16.6819152832031,7.89111900329590,
30.8534927368164,44.4875602722168,
28.8928127288818,58.8056793212891,
12.5544137954712,52.7732505798340,
-11.6976833343506,40.2843093872070,
-40.2465133666992,23.8112411499023,
-61.5538978576660,9.22252845764160,
-52.7457199096680,3.64532184600830,
-7.65729427337647,10.6251087188721,
39.0686340332031,13.1869592666626,
41.4805297851563,-0.938912868499756,
-4.03986024856567,-25.1345539093018,
-46.1498870849609,-32.8671417236328,
-48.5410003662109,-16.5623455047607,
-32.6933708190918,4.00302267074585,
-32.5630722045898,8.99935150146484,
-37.0874023437500,1.85035431385040,
-17.1284770965576,-2.71353578567505,
15.1060037612915,-6.97993469238281,
17.9199256896973,-22.8953399658203,
-9.91808795928955,-47.3177032470703,
-22.0153293609619,-59.2939910888672,
6.96024274826050,-51.3089981079102,
36.4670906066895,-44.4890060424805,
23.8870429992676,-53.0855941772461,
-5.95674562454224,-61.7978782653809,
-0.113114833831787,-41.1139907836914,
39.1321411132813,9.06209850311279,
52.8619689941406,51.9467544555664,
16.0719718933105,57.5517272949219,
-22.7549552917480,36.4868927001953,
-17.3912792205811,21.2569427490234,
12.6916732788086,23.8253593444824,
19.2298393249512,25.2419052124023,
-4.77616596221924,1.89900040626526,
-20.4815006256104,-40.7309112548828,
-3.78305506706238,-71.2167510986328,
23.5526371002197,-60.9015541076660,
34.6811027526856,-14.8162317276001,
32.5569953918457,25.3112869262695,
33.8128967285156,31.3115215301514,
41.0657272338867,8.84845352172852,
44.8994483947754,-7.09572649002075,
46.7334060668945,0.230291545391083,
49.2110900878906,17.6610450744629,
42.6439170837402,18.4378604888916,
13.0405750274658,1.87951707839966,
-23.7254772186279,-14.2908220291138,
-37.6769332885742,-18.9091243743897,
-15.1436424255371,-10.0977134704590,
14.8104763031006,10.0998678207397,
13.7245788574219,33.4382247924805,
-19.6708049774170,39.1223335266113,
-41.7248115539551,12.0604963302612,
-22.6127052307129,-35.6922111511231,
17.7381649017334,-59.6624832153320,
37.8640022277832,-42.7633361816406,
22.1105022430420,-11.3362913131714,
1.24451673030853,-4.44119167327881,
8.56913757324219,-23.9114074707031,
40.5591087341309,-35.0903015136719,
52.3381576538086,-18.5013732910156,
22.3956813812256,6.26076650619507,
-27.2845973968506,14.7037525177002,
-49.5527801513672,12.1012077331543,
-35.6529884338379,16.3848724365234,
-19.0822105407715,27.9811992645264,
-32.3420066833496,26.4218864440918,
-62.0166740417481,0.974652767181397,
-60.6296157836914,-33.1840400695801,
-14.8724575042725,-56.2757301330566,
31.6927185058594,-59.0804481506348,
34.4220466613770,-45.7132720947266,
5.83921623229981,-26.2386322021484,
0.234029233455658,-7.35604333877564,
41.7952156066895,-1.43102753162384,
87.4140472412109,-5.61196327209473,
80.8956909179688,-4.07627677917481,
22.6688156127930,16.7480945587158,
-35.2161483764648,39.7167778015137,
-59.6354179382324,39.8502044677734,
-55.7991409301758,11.3790969848633,
-43.7214393615723,-23.2375507354736,
-25.8763465881348,-34.3189964294434,
6.41442680358887,-15.4845991134644,
35.1576347351074,15.7369108200073,
36.6168251037598,34.7955932617188,
13.9077253341675,26.7668685913086,
-2.37728857994080,-4.38344526290894,
3.38443636894226,-35.6737556457520,
10.6634988784790,-45.4210739135742,
-3.68982291221619,-38.1261940002441,
-24.4998855590820,-41.9624938964844,
-15.4253158569336,-62.8083496093750,
26.7219200134277,-70.1267547607422,
55.6694602966309,-41.3004646301270,
39.9574203491211,-0.201843261718750,
1.06659555435181,9.86894035339356,
-12.8061895370483,-13.8794307708740,
16.0979003906250,-30.9684505462647,
49.0565185546875,-13.7919378280640,
52.5191116333008,15.1897296905518,
30.0640068054199,23.6081256866455,
10.4955492019653,24.8414363861084,
3.50928139686584,40.9244194030762,
-2.82241821289063,55.1329803466797,
-16.5113620758057,35.3437194824219,
-25.5726490020752,-8.50593090057373,
-17.5211296081543,-24.7327880859375,
2.95733642578125,2.18636560440063,
13.6808691024780,31.5973930358887,
-2.88695859909058,19.1517105102539,
-35.6440811157227,-16.2303352355957,
-51.2881660461426,-34.1120452880859,
-28.1636562347412,-30.8709316253662,
22.6996078491211,-32.8121871948242,
61.0621337890625,-37.7272720336914,
58.5421180725098,-12.6116485595703,
29.6805648803711,42.0520706176758,
11.5356273651123,69.7384567260742,
16.5938205718994,39.8499031066895,
34.4908409118652,-9.25385093688965,
45.6448020935059,-23.1568241119385,
45.6695289611816,-4.98789215087891,
33.7742538452148,-0.196514546871185,
11.9474430084229,-28.3602504730225,
-10.2865858078003,-54.8881072998047,
-15.2319793701172,-44.2308883666992,
1.02495861053467,-7.18839359283447,
15.5540924072266,25.6442661285400,
9.07813739776611,43.7619705200195,
-6.12033605575562,49.7457427978516,
-2.99564456939697,44.6324729919434,
17.9773159027100,35.8209419250488,
23.5010986328125,39.9916114807129,
-4.30494976043701,58.2323799133301,
-41.7665824890137,61.3711967468262,
-55.2348365783691,32.2107162475586,
-43.6172981262207,-3.09721732139587,
-30.9555091857910,-3.22939395904541,
-27.0853862762451,28.2505035400391,
-19.6787986755371,42.3231506347656,
0.122499585151672,11.6689968109131,
17.0608749389648,-29.1000099182129,
20.1492290496826,-33.5568656921387,
19.4454631805420,-4.90514755249023,
31.7720661163330,23.9358634948730,
44.3515930175781,39.2747039794922,
28.9981803894043,43.8292236328125,
-13.6587677001953,32.0242996215820,
-43.8822097778320,-5.18123674392700,
-28.7031059265137,-44.5262756347656,
17.2466278076172,-42.8450126647949,
52.2767944335938,7.03551673889160,
48.9814186096191,56.4810829162598,
21.1511611938477,60.2817230224609,
-0.357814550399780,30.6006031036377,
-8.51388072967529,11.8124132156372,
-16.4598140716553,11.4235849380493,
-33.5045623779297,8.27646446228027,
-49.2684936523438,0.870152175426483,
-47.5377922058106,12.6476850509644,
-26.7726001739502,40.6592216491699,
-12.7137918472290,45.4790916442871,
-19.5743083953857,5.62829732894898,
-26.7025356292725,-44.7598114013672,
1.28153920173645,-53.1267280578613,
52.5357818603516,-18.6114349365234,
72.7571411132813,18.8528175354004,
35.0067710876465,35.9842834472656,
-21.3068275451660,44.5885620117188,
-32.0818138122559,53.5362243652344,
2.81767034530640,41.1573791503906,
21.1946716308594,-3.17095851898193,
-6.52483463287354,-48.1320152282715,
-35.6046218872070,-59.5595436096191,
-13.2686014175415,-36.4266395568848,
41.8142967224121,-8.54023170471191,
65.8191909790039,6.63571834564209,
41.2156372070313,15.6565113067627,
15.1441698074341,22.5741386413574,
19.4122428894043,18.7904415130615,
31.1982192993164,1.26402914524078,
10.6221532821655,-13.3650817871094,
-32.2415161132813,-14.2316484451294,
-53.6716651916504,-13.5817003250122,
-35.8637390136719,-21.1754550933838,
-1.83002901077271,-26.4010391235352,
17.8341751098633,-14.3212366104126,
16.9218463897705,4.44061613082886,
8.23058414459229,2.60037231445313,
0.682892799377441,-21.6792030334473,
3.96108150482178,-39.4746818542481,
22.7107715606689,-28.3322315216064,
42.6223258972168,-1.09745657444000,
33.0051422119141,7.25844621658325,
-8.21548271179199,-6.64347457885742,
-52.1960792541504,-15.7913541793823,
-61.3798294067383,0.790139555931091,
-32.2042884826660,24.7875995635986,
0.822767734527588,27.4770584106445,
4.25540494918823,3.99792242050171,
-19.1797447204590,-21.5238323211670,
-37.7570266723633,-19.0247230529785,
-30.3649616241455,11.7272291183472,
2.41032171249390,39.9740486145020,
36.2946395874023,39.3998527526856,
42.3359451293945,18.6921157836914,
21.5208797454834,7.09462833404541,
3.90167164802551,20.7407989501953,
18.3352127075195,39.9277648925781,
49.8975830078125,36.7590141296387,
54.6245727539063,15.8563776016235,
16.0269279479980,15.2666883468628,
-26.9083347320557,43.1671295166016,
-29.8872089385986,53.7164192199707,
-5.40547084808350,12.9153156280518,
-6.85049486160278,-42.6276969909668,
-41.3949012756348,-46.6530227661133,
-56.2827835083008,7.71305465698242,
-16.8471336364746,51.5978126525879,
32.0032768249512,30.6062297821045,
23.9297237396240,-19.3184051513672,
-35.9682350158691,-31.6516799926758,
-76.2118072509766,-4.88180780410767,
-55.1152458190918,12.9929256439209,
-15.3248643875122,4.34055709838867,
-10.8717813491821,4.30729675292969,
-35.2093963623047,25.5368614196777,
-39.0611572265625,28.8276977539063,
-10.0863838195801,-7.95057678222656,
15.9619350433350,-40.6234741210938,
10.2060661315918,-18.5646286010742,
-8.68390274047852,29.9708881378174,
-16.5813236236572,33.2270812988281,
-13.3062763214111,-20.2712707519531,
-9.05653381347656,-64.4937667846680,
2.44921016693115,-42.6080780029297,
30.9691333770752,12.7538585662842,
63.6568183898926,35.9692916870117,
71.4982070922852,15.9563446044922,
42.2830734252930,-9.65772342681885,
0.203851699829102,-16.7895603179932,
-24.1392822265625,-12.5351324081421,
-25.2309494018555,-5.20587396621704,
-13.7861146926880,9.47818565368652,
-3.89154505729675,31.5491981506348,
-7.42744731903076,42.8331336975098,
-26.1060733795166,32.8758811950684,
-42.4720268249512,5.39470720291138,
-35.8924026489258,-22.6108188629150,
-5.74093437194824,-45.0747528076172,
24.3416786193848,-59.1891555786133,
32.3323783874512,-52.5763778686523,
27.4224033355713,-27.6534957885742,
34.6139373779297,-10.0994863510132,
54.1877937316895,-13.9949207305908,
61.6797714233398,-23.2665729522705,
41.3072776794434,-20.9545974731445,
10.1942911148071,-12.2792387008667,
-11.3182353973389,-10.5084733963013,
-21.3834514617920,-16.4738388061523,
-28.3717918395996,-18.9331512451172,
-28.3703498840332,-23.7885990142822,
-12.9038562774658,-49.1760978698731,
6.87739181518555,-76.2880020141602,
8.41059017181397,-60.6889877319336,
-11.6402101516724,0.950942039489746,
-24.0497817993164,46.6802330017090,
-5.73750257492065,30.4769802093506,
26.2531147003174,-5.58109235763550,
36.3660774230957,6.75686120986939,
16.3455314636230,50.8292884826660,
-14.8407859802246,48.6504249572754,
-34.4464187622070,-21.3948192596436,
-40.0786743164063,-79.6797485351563,
-34.0457382202148,-56.2041664123535,
-22.1352138519287,8.63295173645020,
-12.4754524230957,20.0874080657959,
-15.3617792129517,-31.0428619384766,
-25.1871089935303,-70.2620697021484,
-15.7425403594971,-51.2880592346191,
21.1480026245117,-8.03004550933838,
54.7042350769043,16.0493431091309,
48.6760139465332,29.0575771331787,
9.98929405212402,50.0875740051270,
-15.5980157852173,56.1838531494141,
-3.13477373123169,22.3773231506348,
24.2767295837402,-24.5015563964844,
30.1537780761719,-31.0881633758545,
13.4974298477173,2.37747788429260,
1.82535517215729,24.4116859436035,
5.41586303710938,7.72596359252930,
7.30746507644653,-9.67759704589844,
0.314741551876068,14.1632671356201,
-1.14195013046265,52.7957344055176,
14.4853763580322,52.8807678222656,
28.2545661926270,9.47175121307373,
14.1290826797485,-31.7234611511230,
-20.2901573181152,-34.4472465515137,
-37.1855278015137,-6.31771278381348,
-21.2587833404541,15.0080528259277,
-0.568964004516602,11.2358980178833,
-6.09318351745606,-0.0109558701515198,
-29.1822738647461,3.80085730552673,
-35.9538726806641,20.0785198211670,
-14.5688982009888,26.3750667572022,
7.16525983810425,6.87235307693481,
7.99842691421509,-24.7372608184814,
-3.86662697792053,-33.3044700622559,
-9.29728698730469,-8.16072750091553,
-10.3263053894043,18.9387264251709,
-21.1484088897705,13.4441280364990,
-34.1713256835938,-13.9797782897949,
-29.0247097015381,-20.7424678802490,
-3.77481365203857,5.21898221969605,
13.0746698379517,28.1178188323975,
5.06056308746338,9.08468151092529,
-7.33499288558960,-38.7203140258789,
3.21195507049561,-63.8217506408691,
32.1703376770020,-41.0182647705078,
50.2069396972656,1.86903643608093,
45.2685356140137,19.7357463836670,
31.7083911895752,1.58497405052185,
23.1730098724365,-23.9497814178467,
10.6080055236816,-28.7062053680420,
-12.3864631652832,-14.4012851715088,
-33.0266418457031,-2.12315011024475,
-28.5995635986328,-3.51499509811401,
3.39489054679871,-9.73015213012695,
39.1184120178223,-5.53763294219971,
56.3342514038086,7.57386112213135,
54.8107032775879,11.1715803146362,
41.9180603027344,-2.30727934837341,
19.3355083465576,-20.2054500579834,
-13.3762731552124,-20.6939582824707,
-40.6727142333984,0.136398553848267,
-39.5006828308106,18.7014598846436,
-8.88876724243164,10.8425350189209,
16.2661685943604,-20.6822185516357,
-1.36070954799652,-40.4837036132813,
-47.6645278930664,-22.4942073822022,
-66.2987136840820,15.5820074081421,
-30.6919002532959,30.9698638916016,
22.1936416625977,8.43822765350342,
37.2488517761231,-18.6785812377930,
10.1378421783447,-11.1055040359497,
-15.9705381393433,17.4067478179932,
-18.0660152435303,16.3896312713623,
-13.1639041900635,-22.7487964630127,
-14.8178148269653,-53.0193862915039,
-6.70285320281982,-32.8059043884277,
23.0220870971680,17.2235717773438,
38.8393478393555,44.0289764404297,
4.60118198394775,29.8230037689209,
-54.0614395141602,4.52084779739380,
-75.2254486083984,-10.0565176010132,
-39.0457305908203,-16.7966194152832,
10.8814630508423,-16.7443695068359,
28.3479003906250,7.22274017333984,
19.5051784515381,48.9430770874023,
5.00408935546875,62.6075210571289,
-5.71302461624146,15.5931377410889,
-12.8119916915894,-54.6766738891602,
-4.33045101165772,-81.4394149780273,
28.5946884155273,-48.2158393859863,
56.8834114074707,-3.51387858390808,
42.2638130187988,8.29998397827148,
-0.194899082183838,-1.64615511894226,
-20.3825454711914,-2.53165292739868,
0.720487117767334,11.9867897033691,
24.9318027496338,23.7766132354736,
16.0085372924805,31.1822948455811,
-10.2770357131958,47.5989952087402,
-30.3818740844727,64.7527618408203,
-42.1562957763672,57.0919876098633,
-60.4311218261719,22.2956008911133,
-71.8863449096680,-2.38367390632629,
-43.8987770080566,10.1713752746582,
9.98494911193848,37.6132049560547,
36.9202690124512,36.9550170898438,
8.11969947814941,-1.04124665260315,
-40.8628082275391,-38.9369850158691,
-55.8112449645996,-36.5433692932129,
-27.9710102081299,-2.66736507415772,
6.42706394195557,24.3829383850098,
21.3573722839355,23.5699310302734,
16.6933956146240,8.57696342468262,
-0.467560291290283,2.31462860107422,
-30.8716144561768,9.48755073547363,
-63.2085227966309,14.6389122009277,
-68.0310287475586,2.89171218872070,
-26.9786586761475,-17.1627712249756,
37.2743682861328,-26.6053256988525,
74.2730331420898,-23.9894962310791,
59.6604347229004,-19.8162269592285,
21.3235263824463,-20.0072746276855,
-0.341583997011185,-12.6782999038696,
5.59521818161011,7.06045913696289,
17.0827503204346,22.4575786590576,
15.3287973403931,8.83827686309815,
6.36318016052246,-29.1952629089355,
7.61097431182861,-47.7204704284668,
10.6692972183228,-20.6888294219971,
-1.75667953491211,23.2173309326172,
-27.5367527008057,33.7147521972656,
-35.8861007690430,-1.70886468887329,
-6.22434520721436,-40.0622367858887,
43.3075561523438,-38.1707763671875,
70.5543746948242,-1.88248431682587,
57.4951667785645,29.5929012298584,
23.9743576049805,36.7732887268066,
0.936432123184204,31.0248394012451,
-8.73698329925537,26.2553501129150,
-17.7730636596680,15.6160984039307,
-30.6870517730713,-12.5980262756348,
-33.1183547973633,-45.7204933166504,
-14.2048091888428,-58.9323883056641,
17.6035594940186,-46.8651275634766,
41.0336112976074,-27.7699871063232,
45.0511093139648,-19.8391819000244,
38.6543655395508,-21.8561496734619,
36.5298080444336,-23.1306228637695,
37.8446197509766,-15.3711147308350,
35.5267791748047,-0.756095767021179,
30.9804000854492,6.09465312957764,
28.5828304290772,-1.31780362129211,
26.2720222473145,-14.0263319015503,
13.6808109283447,-12.6180715560913,
-6.69387340545654,18.3257408142090,
-14.1529216766357,55.3836555480957,
2.98021316528320,54.7731132507324,
24.0104675292969,10.8833732604980,
14.9336986541748,-28.7788963317871,
-18.3526515960693,-26.8414268493652,
-36.1975975036621,-4.81128978729248,
-21.2003803253174,-1.55304884910584,
-3.42488193511963,-15.5240478515625,
-15.3129940032959,-13.2794456481934,
-38.5271644592285,5.08455562591553,
-33.6771011352539,-5.38340568542481,
-0.489101052284241,-51.4069824218750,
22.9998931884766,-68.2634277343750,
15.6912527084351,-13.5039463043213,
1.40662384033203,52.4211387634277,
4.93513441085815,42.2515411376953,
7.76132726669312,-27.7293491363525,
-13.4882946014404,-61.1226692199707,
-39.5823898315430,-20.0368423461914,
-32.4265441894531,27.0204582214355,
6.66334438323975,20.8932437896729,
36.3063659667969,-6.62485361099243,
29.5235900878906,2.37317347526550,
3.85711693763733,25.4518833160400,
-13.2782468795776,0.373789310455322,
-12.8510599136353,-60.7183799743652,
2.94955110549927,-81.8178100585938,
36.4888687133789,-40.0759811401367,
74.9373626708984,-0.331415057182312,
81.7608413696289,-8.35769367218018,
34.8056564331055,-20.8443355560303,
-29.4382972717285,10.1097965240479,
-49.0498352050781,49.5581207275391,
-11.2937278747559,35.5769691467285,
26.0631885528564,-17.6740245819092,
16.0191383361816,-35.4609146118164,
-22.3442344665527,13.7015991210938,
-42.6187362670898,70.1578216552734,
-26.8719444274902,66.8966751098633,
-2.45454597473145,17.1795139312744,
4.35412597656250,-20.4367885589600,
4.29413747787476,-21.6914234161377,
16.8016242980957,-5.75269508361816,
36.8322448730469,7.16726398468018,
39.8521881103516,6.10276556015015,
17.9889163970947,-13.4475126266480,
-11.8868322372437,-41.9661064147949,
-14.9222660064697,-54.1786651611328,
23.1184883117676,-34.9552688598633,
74.5379486083984,-0.979023456573486,
84.0158386230469,14.5583515167236,
27.6215934753418,6.42939472198486,
-46.6887321472168,6.58112430572510,
-70.0394973754883,23.5911407470703,
-29.9419345855713,26.0064868927002,
17.7056617736816,-5.60196304321289,
21.3633785247803,-32.4570426940918,
0.0783522054553032,-8.30051422119141,
-2.40043401718140,54.6115798950195,
12.0597124099731,91.6534881591797,
-2.18119192123413,67.8390426635742,
-51.2517318725586,15.4046840667725,
-80.0755538940430,-19.3606853485107,
-49.0468673706055,-33.6539421081543,
14.5340709686279,-47.9421691894531,
50.3780021667481,-54.2175559997559,
42.0435142517090,-24.2122859954834,
21.4578094482422,38.5040168762207,
12.6045417785645,84.3278579711914,
7.33789587020874,75.0753479003906,
-1.09607875347137,28.7996177673340,
-8.03245639801025,-9.37629699707031,
-12.9117794036865,-17.2579059600830,
-30.9307842254639,-1.39003467559814,
-59.6985130310059,17.0663757324219,
-68.4516296386719,24.8224258422852,
-39.3161582946777,21.7871398925781,
-7.77069282531738,14.6922788619995,
-18.0397739410400,10.9448041915894,
-61.2306709289551,14.5875120162964,
-82.6668777465820,14.0899400711060,
-53.4285774230957,-0.499007225036621,
-5.12691307067871,-16.4803161621094,
15.9568128585815,-19.4727210998535,
8.32653999328613,-15.3318099975586,
6.10245418548584,-19.6939811706543,
23.2823925018311,-24.5681190490723,
37.7540626525879,-4.21299457550049,
26.9779663085938,40.0429115295410,
-2.61555814743042,64.0970153808594,
-32.1531715393066,35.3228950500488,
-51.5944824218750,-17.8750076293945,
-55.6680374145508,-41.0630760192871,
-41.3594322204590,-27.7992401123047,
-19.9985637664795,-20.6241016387939,
-7.51530122756958,-42.4077186584473,
-18.5706577301025,-57.8563613891602,
-46.9411888122559,-30.5949230194092,
-68.0726928710938,15.1088275909424,
-59.3143005371094,23.7833709716797,
-23.1411247253418,-13.0608186721802,
22.1170902252197,-47.7011032104492,
45.9042816162109,-38.8852272033691,
25.6637153625488,-2.89619421958923,
-17.9894351959229,18.0920810699463,
-30.8244209289551,11.0490074157715,
10.9883308410645,-1.57508301734924,
61.3130073547363,-1.76896357536316,
53.4060821533203,5.72668695449829,
-12.3675136566162,9.52068138122559,
-56.6134529113770,4.77617597579956,
-26.2830848693848,-9.81748771667481,
36.2960624694824,-23.9556007385254,
50.4729270935059,-22.8286399841309,
7.23973941802979,1.71643805503845,
-28.3809623718262,27.3299770355225,
-15.8982362747192,22.5097427368164,
6.13350391387939,-14.8541841506958,
-4.42261028289795,-46.8616905212402,
-32.8647270202637,-41.4529266357422,
-35.1175613403320,-11.4094953536987,
-8.85944175720215,-2.30590605735779,
5.53913021087647,-24.7490329742432,
-9.67795467376709,-46.5169219970703,
-25.2221260070801,-40.2686309814453,
-13.9887075424194,-17.3099956512451,
13.3568792343140,-7.81950712203980,
26.4124660491943,-22.3905429840088,
19.9410610198975,-38.0784416198731,
11.1342906951904,-29.3962707519531,
9.01659393310547,5.22381877899170,
12.3132619857788,40.6524200439453,
20.7455215454102,52.0616378784180,
31.3837337493897,36.0340614318848,
30.7344875335693,19.9882850646973,
9.38299655914307,29.3438529968262,
-18.5927429199219,59.1222267150879,
-21.2133731842041,68.9032287597656,
9.71702289581299,32.3369560241699,
43.9394187927246,-19.8124179840088,
44.3194694519043,-32.6352233886719,
14.8447360992432,1.02681350708008,
-6.16774320602417,38.0057754516602,
2.67432689666748,35.3793106079102,
21.1988773345947,12.7332725524902,
17.2118911743164,15.5423574447632,
-13.1161565780640,49.8046226501465,
-43.9058189392090,71.8490829467773,
-53.2667579650879,48.1537322998047,
-46.4539070129395,-5.03791618347168,
-36.2640953063965,-47.5495567321777,
-23.8911819458008,-58.0278511047363,
-4.13685083389282,-47.6198806762695,
20.1066303253174,-30.8503952026367,
28.7221736907959,-14.9422140121460,
16.2157688140869,-7.04137229919434,
-3.35099148750305,-19.5421905517578,
-10.7795648574829,-48.3251075744629,
-3.53931975364685,-72.5681915283203,
6.50308227539063,-68.7422332763672,
4.94418191909790,-37.4465408325195,
-5.92974185943604,-2.53948783874512,
-17.5905513763428,15.6228218078613,
-31.8868656158447,15.8163728713989,
-48.9588317871094,11.9671916961670,
-54.3259849548340,8.98508644104004,
-30.6071472167969,8.33668041229248,
16.4206504821777,6.61250448226929,
43.3626251220703,7.75674343109131,
18.2765369415283,13.2273674011230,
-42.1639823913574,15.4509248733521,
-74.4594039916992,10.3188304901123,
-49.1029357910156,1.59732210636139,
-8.98282623291016,-3.68165516853333,
-7.38134574890137,-9.27023887634277,
-39.1791000366211,-19.9272117614746,
-47.1647644042969,-30.7049789428711,
-8.28887176513672,-29.2519969940186,
33.1637191772461,-7.61829757690430,
29.5057430267334,21.6393795013428,
-2.46991896629334,40.9212760925293,
-12.4670867919922,42.2257575988770,
0.919122457504273,28.9664573669434,
-7.28969955444336,11.6801595687866,
-43.4213104248047,-5.80341672897339,
-55.3162727355957,-20.5585823059082,
-6.75109291076660,-32.7083435058594,
56.6161499023438,-38.4056243896484,
58.9336280822754,-32.1976318359375,
-0.0754851102828980,-10.0574731826782,
-50.0213699340820,15.8153762817383,
-45.8855476379395,27.1061668395996,
-18.4901905059814,18.0086746215820,
-14.5821485519409,0.0784158706665039,
-24.8881320953369,-15.9776992797852,
-11.0149812698364,-25.2567806243897,
30.1470794677734,-22.4395809173584,
52.9749488830566,0.798259735107422,
35.5126228332520,38.3953704833984,
2.28388428688049,60.2882423400879,
-13.2618513107300,50.6370887756348,
-8.21629810333252,29.7139606475830,
-4.10407733917236,32.8749694824219,
-8.77896785736084,56.5264167785645,
-21.0388202667236,59.9696769714356,
-36.5799446105957,30.1763362884522,
-57.3062095642090,-1.52102077007294,
-70.0710525512695,-5.60595273971558,
-57.0537414550781,0.851958453655243,
-21.1427574157715,-10.5672588348389,
12.7335662841797,-31.2472667694092,
32.7332878112793,-32.5498046875000,
44.0110969543457,-9.82561779022217,
52.6281623840332,9.58710670471191,
46.5989952087402,11.9178962707520,
16.9643573760986,13.5346708297730,
-22.6493301391602,23.8493595123291,
-46.2141532897949,22.0205249786377,
-50.6934280395508,-7.57964611053467,
-49.3573036193848,-42.7541198730469,
-42.8867454528809,-58.8974418640137,
-11.9111509323120,-54.0399322509766,
44.2672996520996,-44.3098793029785,
86.9883422851563,-27.2159938812256,
78.9058609008789,-1.94622492790222,
30.5835151672363,13.0555772781372,
0.0802739262580872,-2.99095153808594,
14.5985193252563,-31.9983024597168,
48.3568496704102,-28.9254112243652,
50.7521247863770,11.5331764221191,
15.3548078536987,39.7929420471191,
-17.2113609313965,13.4274425506592,
-12.9908008575439,-39.1823387145996,
17.3944511413574,-53.4523200988770,
39.7658958435059,-11.3472757339478,
40.6558036804199,43.1499061584473,
28.0234832763672,63.5090751647949,
15.8385477066040,48.1601600646973,
1.97645008563995,21.6434669494629,
-11.7635641098022,3.54080533981323,
-15.2310075759888,-10.1123142242432,
2.76443600654602,-17.7821941375732,
36.4859008789063,-14.9058732986450,
61.7679214477539,0.0136826634407043,
65.5033721923828,16.8178882598877,
47.6084632873535,24.1057071685791,
21.8171195983887,16.5405216217041,
-0.872409701347351,-0.384727716445923,
-17.4651203155518,-19.0581340789795,
-29.1845760345459,-28.5674896240234,
-35.4367828369141,-25.3857765197754,
-36.0841598510742,-18.9269981384277,
-32.9850387573242,-19.4260101318359,
-27.5053634643555,-30.9526023864746,
-23.7651977539063,-48.7272338867188,
-15.0589103698730,-60.5072708129883,
6.33319187164307,-61.2964897155762,
38.4764900207520,-51.5251884460449,
58.9983749389648,-35.8558387756348,
44.6462593078613,-17.8482170104980,
-2.56792855262756,1.65134727954865,
-44.8240547180176,20.5318546295166,
-45.7088737487793,31.5467700958252,
-5.98960971832275,28.2736148834229,
30.5455837249756,10.6778335571289,
30.6870822906494,-6.93146371841431,
2.02624130249023,-12.5984210968018,
-13.4925403594971,-4.69454717636108,
5.66872882843018,5.40976619720459,
36.0284767150879,9.76282501220703,
39.8981742858887,3.25913548469543,
20.8770198822022,-7.86743783950806,
16.2889652252197,-16.0448951721191,
39.6293678283691,-13.7030582427979,
54.4498634338379,-0.633009433746338,
22.6351699829102,14.4016656875610,
-35.3734283447266,16.8121528625488,
-60.7718429565430,5.97810745239258,
-29.0651836395264,-11.5328397750855,
8.95661354064941,-27.4465827941895,
0.224314212799072,-37.4950218200684,
-33.1684951782227,-35.9427299499512,
-37.2830886840820,-19.6498126983643,
-5.80495595932007,-6.84988117218018,
13.1744670867920,-18.7687702178955,
-1.91443920135498,-51.3389244079590,
-14.0349254608154,-66.1343917846680,
10.9315538406372,-34.5972061157227,
43.3835639953613,24.1007804870605,
35.4040718078613,58.6546440124512,
-3.77437758445740,43.6184043884277,
-21.7395229339600,-0.622612953186035,
-11.3078880310059,-35.1010208129883,
-15.3015537261963,-39.8521652221680,
-43.1089591979981,-20.4130764007568,
-45.3423080444336,6.95023202896118,
4.63257503509522,22.5300140380859,
54.0979461669922,10.7426185607910,
45.5990600585938,-17.0070590972900,
7.04439496994019,-35.1612777709961,
7.75023126602173,-30.9390106201172,
47.9335823059082,-19.5881195068359,
55.8207740783691,-16.1926727294922,
4.32724189758301,-20.5003261566162,
-40.3368682861328,-24.2566757202148,
-19.4693031311035,-25.0416107177734,
25.4939270019531,-21.8343372344971,
12.9398937225342,-7.07035970687866,
-48.7920150756836,16.4460849761963,
-76.9007339477539,21.2524662017822,
-32.3042335510254,-9.42142391204834,
27.6331939697266,-43.6616058349609,
35.4205398559570,-35.3238410949707,
-0.0850667953491211,12.6648139953613,
-24.6467952728272,41.3068161010742,
-18.4313163757324,22.6291198730469,
-12.9957656860352,-4.73614549636841,
-26.0275478363037,2.31051731109619,
-34.9598350524902,32.9745368957520,
-22.0311813354492,50.5108680725098,
-0.0656547546386719,42.8628234863281,
13.0241184234619,26.9348278045654,
20.6823329925537,10.2136211395264,
30.8089485168457,-17.2759876251221,
40.1987342834473,-40.0634651184082,
40.3121910095215,-32.9652709960938,
33.7118568420410,-5.46587133407593,
32.5514450073242,0.422599077224731,
35.4166374206543,-20.4942188262939,
28.2888622283936,-18.2932281494141,
16.9093399047852,23.5193080902100,
23.5593070983887,50.7673110961914,
45.6225318908691,22.7512989044189,
49.6561355590820,-19.8516407012939,
20.8991088867188,-11.4014797210693,
-14.3895759582520,34.6924285888672,
-25.6843643188477,41.9973030090332,
-18.3410415649414,-12.1421813964844,
-17.8279247283936,-57.9810523986816,
-25.0580120086670,-49.1461944580078,
-13.4401912689209,-27.5371837615967,
22.2643146514893,-34.7717361450195,
51.0376243591309,-34.9444007873535,
45.2943000793457,18.6193046569824,
18.5987167358398,75.9782180786133,
-5.93029737472534,54.3903923034668,
-19.5436496734619,-29.0059299468994,
-22.5922298431397,-66.4096984863281,
-3.86629676818848,-11.8881244659424,
27.6095027923584,53.6038970947266,
37.0555267333984,45.4157981872559,
2.72869586944580,-0.678912043571472,
-38.7792015075684,1.26965618133545,
-38.7262458801270,45.3838539123535,
0.362493276596069,49.4008140563965,
22.7802066802979,-7.68578577041626,
4.27382373809814,-52.3302803039551,
-18.0347061157227,-42.3255386352539,
-6.48820114135742,-18.3537044525147,
19.8313503265381,-26.1550979614258,
26.8760967254639,-38.9135169982910,
25.5324821472168,-11.1830005645752,
37.9365119934082,34.6159744262695,
46.2230491638184,43.1297645568848,
17.9939613342285,10.9231433868408,
-32.7956619262695,-2.24817800521851,
-54.8977737426758,29.8475284576416,
-31.8183498382568,57.2608985900879,
-8.30291461944580,39.6603813171387,
-19.9799919128418,4.11000299453735,
-45.8344993591309,-11.7213125228882,
-49.4750213623047,-9.71574974060059,
-35.1207313537598,-14.0674343109131,
-29.1360321044922,-19.7499294281006,
-22.8796234130859,-7.66944932937622,
0.00900799036026001,19.4557437896729,
20.3776149749756,35.7561683654785,
2.61468362808228,36.5118484497070,
-37.9453468322754,37.3179588317871,
-47.8151359558106,40.2139968872070,
-8.63885402679443,22.4734859466553,
25.9952259063721,-14.0733795166016,
7.40857267379761,-29.2265205383301,
-38.5223426818848,-6.92275428771973,
-49.1031188964844,14.5395488739014,
-14.1040840148926,-2.58178019523621,
15.0788106918335,-40.9511260986328,
9.91787052154541,-53.4929656982422,
-1.64326572418213,-28.6397209167480,
13.6524801254272,2.21402740478516,
41.6839828491211,11.2841148376465,
47.6770935058594,7.43741607666016,
33.7641754150391,1.70238614082336,
28.9532947540283,-11.6472768783569,
39.6253051757813,-30.4720249176025,
38.0004081726074,-32.5562477111816,
7.29778575897217,-7.95675516128540,
-28.0387496948242,15.0187788009644,
-28.6531105041504,2.54131174087524,
3.77932119369507,-31.2042865753174,
29.1556930541992,-40.5663833618164,
25.6147975921631,-10.8141059875488,
12.8657207489014,26.9642925262451,
13.1566896438599,40.3646087646484,
21.1090354919434,34.2994613647461,
7.27652502059937,35.5507659912109,
-35.1487083435059,50.2042007446289,
-68.3419876098633,52.0908508300781,
-57.7006340026856,25.0004959106445,
-17.3782730102539,-17.5563068389893,
8.36391544342041,-48.5528526306152,
-5.72332763671875,-48.3904762268066,
-28.5041007995605,-25.5822219848633,
-18.7475872039795,-5.83908319473267,
22.0059013366699,-7.81675243377686,
46.8796844482422,-20.4021129608154,
20.5397663116455,-12.6177139282227,
-28.5129566192627,22.8896064758301,
-43.8812370300293,51.7632026672363,
-8.71946144104004,42.0801849365234,
32.5187988281250,1.64377975463867,
27.4497318267822,-22.7983646392822,
-20.5619106292725,-2.05095243453980,
-55.3675460815430,28.8903903961182,
-33.9014205932617,22.0171680450439,
23.7710571289063,-21.3878459930420,
64.8848266601563,-53.3516693115234,
64.6293258666992,-48.3526344299316,
35.8363113403320,-18.0917739868164,
2.30657482147217,10.0069379806519,
-24.1839103698730,30.3555889129639,
-38.3449249267578,36.8696556091309,
-37.6437911987305,10.8789787292480,
-27.2222061157227,-46.5601806640625,
-23.8804759979248,-81.4677734375000,
-23.6949481964111,-45.5530014038086,
-7.58480739593506,27.5919132232666,
25.5720634460449,52.9048995971680,
47.3012084960938,5.63218688964844,
28.0949611663818,-39.0980682373047,
-12.4137239456177,-18.8527202606201,
-29.6116142272949,24.3737354278564,
-12.2462806701660,10.4341573715210,
3.17780923843384,-55.8353576660156,
-5.64166021347046,-86.9907531738281,
-16.8870754241943,-42.6128120422363,
-3.32847094535828,11.6271200180054,
30.2558097839355,5.67506837844849,
55.2834548950195,-35.7599105834961,
61.2514419555664,-43.8544692993164,
54.0117721557617,-7.06994915008545,
34.0673217773438,19.1198558807373,
-3.51620149612427,2.33993482589722,
-35.6723213195801,-24.1483440399170,
-28.1531047821045,-30.1849498748779,
16.5788917541504,-25.0644893646240,
55.5943145751953,-24.4876194000244,
56.5833587646484,-19.9605140686035,
36.1974716186523,5.38452053070068,
21.3296127319336,38.5119285583496,
5.33986330032349,41.9238014221191,
-28.4334487915039,11.8898248672485,
-65.2891159057617,-14.5097169876099,
-65.5817337036133,-11.5470228195190,
-23.2975788116455,13.7401905059814,
14.1809368133545,34.1115646362305,
6.27976560592651,29.3988018035889,
-24.7174549102783,-3.17637395858765,
-29.1372661590576,-34.9802436828613,
4.85632896423340,-32.1530952453613,
36.5976219177246,8.30616950988770,
30.6962318420410,48.3470382690430,
-1.29012560844421,46.8782958984375,
-25.6152381896973,13.3120737075806,
-21.9911651611328,2.32490563392639,
0.756912112236023,36.7683372497559,
22.3563613891602,69.4166030883789,
31.2484779357910,49.1120681762695,
23.6053199768066,-4.72807455062866,
4.23949527740479,-30.6287803649902,
-12.0644149780273,-15.7815656661987,
-15.8568134307861,-9.47955894470215,
-11.9229192733765,-39.0341758728027,
-12.0602884292603,-63.8535041809082,
-15.6155376434326,-35.5348968505859,
-15.8084697723389,19.5803546905518,
-15.9594001770020,37.6136703491211,
-23.3477191925049,7.53950691223145,
-34.1350326538086,-16.5003395080566,
-35.8064308166504,3.17668938636780,
-20.5189971923828,33.3598136901856,
-0.803450822830200,18.9075565338135,
8.89043235778809,-26.3523502349854,
13.3645668029785,-47.6402740478516,
24.1938705444336,-18.3627204895020,
35.6517906188965,26.8916549682617,
38.3164100646973,45.2765083312988,
34.7574348449707,28.3113746643066,
35.1427955627441,5.87856817245483,
32.9974403381348,6.85438203811646,
14.0941419601440,28.1558609008789,
-14.1673851013184,44.7163276672363,
-16.8204288482666,34.4525299072266,
16.7683849334717,2.39194512367249,
47.8014984130859,-13.1890106201172,
31.7138080596924,15.7402362823486,
-20.5098495483398,58.0690727233887,
-55.5003890991211,51.5480041503906,
-44.3934669494629,-11.7385540008545,
-21.4217166900635,-67.2092056274414,
-26.2221221923828,-60.8800086975098,
-47.7892341613770,-15.4245929718018,
-46.2643966674805,2.34760975837708,
-12.3025255203247,-18.8082523345947,
21.2182750701904,-23.2376537322998,
20.7357940673828,21.4487571716309,
-11.6561002731323,65.8312225341797,
-40.3483238220215,55.1382484436035,
-38.0522308349609,7.87336492538452,
-8.11812686920166,-17.5132274627686,
20.6280879974365,-5.97164201736450,
21.0333175659180,-2.16391515731812,
-6.36519861221314,-26.2860260009766,
-33.3259811401367,-40.4880180358887,
-32.4949760437012,-12.9682779312134,
-14.2530918121338,21.2756366729736,
-11.9692420959473,11.1999263763428,
-25.1193103790283,-36.7656593322754,
-19.5555458068848,-66.2906494140625,
16.0773410797119,-47.8591003417969,
45.6812286376953,-19.7893009185791,
29.9454879760742,-23.4399223327637,
-15.8887338638306,-41.5716476440430,
-39.3690910339356,-30.2011528015137,
-22.0281314849854,10.5775156021118,
0.171730697154999,43.1401138305664,
1.67774605751038,38.7011184692383,
-3.18709778785706,13.2699785232544,
1.99474108219147,3.28049397468567,
3.83228921890259,13.4981632232666,
-12.8890905380249,21.1925735473633,
-24.5526084899902,14.8217592239380,
-2.52121424674988,9.91743469238281,
31.0193023681641,22.6567592620850,
22.6784057617188,42.0302429199219,
-36.2289695739746,41.2344474792481,
-84.3629074096680,6.84132099151611,
-72.1777267456055,-36.5098228454590,
-22.7682285308838,-43.6399688720703,
1.00065732002258,-2.87356472015381,
-16.4814014434814,44.8073997497559,
-31.3031749725342,45.7414855957031,
-10.7271757125855,-2.54912137985230,
21.6377105712891,-51.0961189270020,
28.9944076538086,-51.7382087707520,
12.6249284744263,-13.3147258758545,
7.97836875915527,20.6599121093750,
26.6075096130371,28.0970516204834,
37.8596992492676,28.6272811889648,
14.8450946807861,37.8138198852539,
-31.6519813537598,44.2250251770020,
-62.1155090332031,31.8612117767334,
-55.4229049682617,7.92435550689697,
-26.0061893463135,-10.4499406814575,
4.25854110717773,-19.1175594329834,
29.1190338134766,-25.8091220855713,
39.6983222961426,-25.5653438568115,
31.7232456207275,-6.35662078857422,
8.47556972503662,19.5322704315186,
-5.83640861511231,23.4614601135254,
8.70903587341309,3.32774400711060,
38.8065147399902,-10.0662279129028,
41.0541534423828,8.84999561309815,
-1.63939499855042,40.2404479980469,
-53.3803749084473,42.0013122558594,
-65.9564971923828,9.97815322875977,
-31.0300064086914,-22.0568542480469,
10.6476888656616,-27.7104396820068,
20.8472328186035,-17.0272312164307,
4.88471412658691,-9.66404819488525,
2.35275745391846,-10.0592088699341,
26.6199226379395,-6.05564546585083,
53.5464057922363,6.91215276718140,
51.6064529418945,13.4735822677612,
23.2322349548340,2.67334032058716,
3.42845344543457,-18.9499416351318,
15.1624460220337,-29.7738418579102,
38.7188415527344,-13.2580585479736,
34.0866546630859,29.9699726104736,
-9.34260177612305,68.8821640014648,
-54.2449836730957,62.6528358459473,
-66.5008010864258,11.8629341125488,
-52.0419082641602,-30.5315723419189,
-40.0208511352539,-23.1816768646240,
-46.1802062988281,12.7075862884521,
-47.3929748535156,16.9621162414551,
-29.1733169555664,-30.2747097015381,
-8.87097454071045,-73.9661941528320,
-9.64412117004395,-62.8970031738281,
-23.1151924133301,-19.4706954956055,
-18.1965293884277,-0.400780916213989,
8.22122955322266,-10.0148696899414,
28.5758266448975,0.177302837371826,
24.6465110778809,38.2292518615723,
15.4349613189697,52.5871810913086,
23.6652545928955,15.5810832977295,
38.0127601623535,-27.4340877532959,
27.4127750396729,-15.9885063171387,
-12.1452093124390,30.5531806945801,
-51.6704597473145,40.8950271606445,
-66.1322250366211,-5.58483314514160,
-58.7218437194824,-49.2013702392578,
-37.0494613647461,-40.9619178771973,
-3.51059556007385,-0.878544092178345,
34.8318824768066,22.6529598236084,
52.8038711547852,19.5877342224121,
34.6568679809570,7.18280506134033,
2.73241949081421,-14.4883289337158,
-4.08858823776245,-45.6624221801758,
16.5243377685547,-58.4541358947754,
28.5418682098389,-22.6954803466797,
8.67517089843750,36.3177947998047,
-22.2754192352295,51.2659721374512,
-22.4116554260254,3.13057065010071,
15.8044099807739,-46.2284545898438,
49.7685699462891,-30.0382347106934,
40.7160835266113,36.6081962585449,
0.813079357147217,77.9158096313477,
-22.1618061065674,58.3882713317871,
2.08929157257080,18.4336433410645,
43.0976867675781,10.0401086807251,
48.0924034118652,33.2168960571289,
1.57447171211243,51.1390075683594,
-53.6038208007813,44.4834175109863,
-67.4318618774414,31.3487510681152,
-45.3563957214356,26.8669052124023,
-28.0369987487793,19.0475940704346,
-31.2943191528320,-3.99284601211548,
-29.9468250274658,-26.1251678466797,
-5.09656429290772,-18.6926631927490,
24.1923103332520,15.2122764587402,
25.5340785980225,37.3453445434570,
4.85120820999146,23.7090816497803,
-4.98792123794556,-11.0374984741211,
2.49147105216980,-24.2471446990967,
3.66666913032532,2.30733466148376,
-11.8138628005981,41.8241386413574,
-21.3569011688232,56.9580764770508,
-8.75457859039307,39.0775070190430,
3.22746562957764,9.60446071624756,
-15.4061203002930,-3.72430396080017,
-45.9521026611328,4.51716566085815,
-47.2981567382813,15.0336856842041,
-14.3616161346436,8.95787429809570,
13.1325273513794,-11.0069103240967,
2.48143291473389,-24.1266403198242,
-27.1025257110596,-24.1255741119385,
-39.6072311401367,-21.4520454406738,
-29.3394565582275,-22.2113018035889,
-16.1734104156494,-23.7286586761475,
-9.61049747467041,-19.9358081817627,
-1.93582856655121,-20.1571617126465,
2.82258319854736,-36.1809349060059,
-3.85846424102783,-55.7635803222656,
-9.69270610809326,-60.6522750854492,
8.76811981201172,-52.3727226257324,
46.9972839355469,-47.3630828857422,
66.1161651611328,-44.7647819519043,
41.6902694702148,-23.8963775634766,
-1.58751428127289,9.84375095367432,
-20.3663768768311,16.6174945831299,
-6.96145629882813,-16.9081821441650,
3.98671054840088,-46.8156509399414,
-3.50319457054138,-23.2884330749512,
-16.4381942749023,33.4673080444336,
-23.8485469818115,58.7037582397461,
-33.5362586975098,26.8839759826660,
-43.4903221130371,-17.8743190765381,
-35.3266296386719,-32.8704032897949,
-4.20184850692749,-33.8785591125488,
23.5328884124756,-46.1605987548828,
22.7104358673096,-53.7314910888672,
10.3569192886353,-28.2066116333008,
16.4703044891357,4.76168537139893,
35.1261520385742,1.76647818088532,
31.8993053436279,-36.9088859558106,
1.37783908843994,-54.5254859924316,
-9.78088760375977,-25.0168304443359,
20.2476863861084,16.6660594940186,
55.7694778442383,29.1797351837158,
52.5340347290039,22.4212303161621,
18.8250446319580,24.3588180541992,
-1.12553215026855,26.4064178466797,
4.40468311309814,0.587287187576294,
7.45201349258423,-39.5432510375977,
-9.42906284332275,-45.6017913818359,
-29.2520370483398,-11.9832172393799,
-33.5763015747070,11.9723901748657,
-31.3493938446045,-9.02562046051025,
-33.1895332336426,-51.7395439147949,
-20.7878055572510,-72.8252563476563,
20.0497322082520,-58.5727539062500,
62.0017471313477,-31.9224624633789,
62.2909507751465,-5.42817974090576,
21.7897834777832,21.7308959960938,
-15.4008235931396,41.6893730163574,
-18.1999797821045,34.7161750793457,
5.00448513031006,6.70681810379028,
25.2956333160400,-12.3297128677368,
25.9264221191406,-11.9764699935913,
12.8422307968140,-6.63434123992920,
-3.25211787223816,-5.00504446029663,
-10.5968189239502,11.3553771972656,
-2.21621656417847,49.0582771301270,
14.6828565597534,69.9015045166016,
15.5095281600952,35.7376289367676,
-3.76112413406372,-35.7162628173828,
-18.0436401367188,-78.4298171997070,
-11.3563385009766,-59.5140647888184,
-9.82480430603027,-18.6183929443359,
-35.1702537536621,-2.33653783798218,
-65.2769088745117,-7.46876811981201,
-63.5531768798828,0.559966802597046,
-30.7035999298096,23.2377662658691,
-5.81401109695435,24.3308963775635,
-7.36219215393066,-8.31547164916992,
-7.75847959518433,-39.7138137817383,
10.4179162979126,-33.0442352294922,
12.1629333496094,1.02653527259827,
-23.7454147338867,24.5219554901123,
-54.8564224243164,23.6443405151367,
-29.8763980865479,20.9215660095215,
23.9755401611328,30.3326797485352,
26.9028949737549,37.6657333374023,
-35.7280082702637,26.2090969085693,
-86.0289382934570,6.86896324157715,
-59.9709930419922,-4.69512939453125,
-1.52161347866058,-1.70119321346283,
5.24259662628174,6.32960605621338,
-40.4362907409668,12.5854616165161,
-66.9017028808594,16.4658241271973,
-38.4785156250000,19.2087497711182,
-7.93557262420654,19.2761878967285,
-27.2773189544678,13.0768280029297,
-64.8210220336914,-0.551153004169464,
-57.8047714233398,-20.2305259704590,
-6.56045007705689,-43.1019439697266,
28.1117286682129,-58.0735092163086,
13.9985485076904,-59.5333557128906,
-9.11822319030762,-55.9192886352539,
4.64355611801148,-53.4530296325684,
46.6031532287598,-42.2322082519531,
61.6903800964356,-20.8760147094727,
26.6903038024902,-5.93698692321777,
-16.2583961486816,-10.8063926696777,
-24.3888969421387,-20.6720695495605,
7.21967697143555,-12.8663721084595,
43.9873542785645,5.30890941619873,
50.0037612915039,5.65740489959717,
19.8784980773926,-12.5595741271973,
-17.8627872467041,-12.9297838211060,
-32.7479591369629,20.6730308532715,
-18.4597682952881,42.3980751037598,
6.08104562759399,14.5738945007324,
20.7664375305176,-29.6042156219482,
24.9071121215820,-23.9994049072266,
32.7238807678223,28.0493354797363,
40.4839439392090,54.3282356262207,
21.5089378356934,19.5352687835693,
-30.4833393096924,-20.5955638885498,
-72.5775527954102,-11.9697427749634,
-61.3741531372070,21.0054168701172,
-5.66429758071899,13.2255392074585,
37.6362838745117,-32.5586318969727,
30.2546081542969,-48.3312149047852,
-6.07437849044800,-4.05786132812500,
-28.1710529327393,40.9099693298340,
-30.5401020050049,27.7140045166016,
-33.0751266479492,-26.7412319183350,
-41.4902763366699,-62.5927467346191,
-38.3997879028320,-58.9656333923340,
-17.4254379272461,-41.9945297241211,
0.297145187854767,-31.5020637512207,
1.81721127033234,-25.4355468750000,
0.553377091884613,-27.3935737609863,
9.46328639984131,-42.2143936157227,
19.6250991821289,-59.9333076477051,
14.6445865631104,-51.1731109619141,
1.69505167007446,-14.9208860397339,
-4.12532377243042,4.05599164962769,
2.30449819564819,-25.3045749664307,
8.43254852294922,-70.2342147827148,
8.62231159210205,-74.7656326293945,
12.8951826095581,-35.7597427368164,
20.3140392303467,4.51287698745728,
18.4342079162598,16.6141262054443,
7.66068983078003,6.99853849411011,
6.33040952682495,0.843547165393829,
18.7795047760010,5.18975830078125,
22.8561477661133,15.5628986358643,
1.48662090301514,31.7810325622559,
-31.3597049713135,44.0749740600586,
-46.2155532836914,36.1337585449219,
-36.4781150817871,6.66940116882324,
-24.2817726135254,-15.9575309753418,
-20.8989734649658,-7.95726442337036,
-13.2305803298950,5.21509075164795,
5.46431207656860,-7.29009628295898,
21.7532138824463,-28.3350257873535,
23.0087108612061,-15.0969295501709,
16.9519672393799,38.4764785766602,
14.6115932464600,84.9383239746094,
4.37704753875732,76.7572555541992,
-26.5749320983887,27.1012496948242,
-58.5065498352051,-18.4855270385742,
-55.4902076721191,-36.1116561889648,
-16.4429950714111,-31.2244663238525,
16.4150524139404,-8.38300228118897,
4.77911472320557,23.0151252746582,
-35.7943954467773,33.5786285400391,
-52.2558517456055,-1.28641772270203,
-24.2210941314697,-52.0582351684570,
20.4723243713379,-55.7537345886231,
39.1520652770996,8.16790962219238,
18.9511871337891,78.8579864501953,
-20.2687683105469,86.3468399047852,
-45.9133033752441,35.4952697753906,
-41.3457450866699,-13.2616748809814,
-17.8970012664795,-27.2167606353760,
0.00783510506153107,-31.6321468353272,
1.05725264549255,-54.0755577087402,
3.56214308738709,-69.3729934692383,
26.8656654357910,-43.0574684143066,
56.3877143859863,9.34035015106201,
54.2340812683106,41.5310783386231,
7.44357776641846,33.4432678222656,
-44.2269706726074,15.8711719512939,
-51.0344848632813,24.2237033843994,
-17.8292865753174,46.9883155822754,
9.22510147094727,50.4008789062500,
1.13802123069763,21.0914039611816,
-22.7876873016357,-11.3134031295776,
-29.6786098480225,-15.7171020507813,
-14.4805660247803,3.65531134605408,
3.39388132095337,16.6608772277832,
15.3052158355713,2.57670998573303,
25.6675243377686,-26.9695510864258,
35.3724327087402,-37.7403602600098,
32.3818511962891,-11.4785919189453,
15.1460599899292,34.3883972167969,
-5.61295604705811,57.4676551818848,
-17.4187602996826,36.2373428344727,
-22.8333911895752,-13.1035270690918,
-32.6985473632813,-53.0408973693848,
-43.0739288330078,-57.5752906799316,
-42.6536560058594,-32.8769035339356,
-34.5647315979004,-6.32860517501831,
-31.5197219848633,-1.66447627544403,
-35.3248596191406,-24.1992568969727,
-28.8125762939453,-56.0803909301758,
-2.99480772018433,-66.7126083374023,
17.7161064147949,-42.5176925659180,
4.51289463043213,-6.43388509750366,
-32.6230812072754,4.10728502273560,
-44.1135406494141,-20.1108837127686,
-3.29436826705933,-47.6750564575195,
50.7623786926270,-50.1467628479004,
61.5898551940918,-35.0988235473633,
25.8707199096680,-25.1655178070068,
-5.31623077392578,-20.6105079650879,
4.71373271942139,-4.36166000366211,
29.1700210571289,21.9693660736084,
25.9819068908691,26.2226428985596,
-0.840948462486267,-4.83963775634766,
-14.1414585113525,-33.0349693298340,
-1.74769341945648,-24.3434467315674,
9.50913333892822,3.16164398193359,
-4.39516925811768,10.4316272735596,
-30.0123310089111,-2.86347627639771,
-34.0228424072266,5.62220954895020,
-12.2321386337280,44.1112823486328,
6.39996433258057,64.1962127685547,
-2.60243415832520,33.4443130493164,
-26.1741580963135,-11.1336536407471,
-32.1564636230469,-14.1180381774902,
-2.96463894844055,17.8270301818848,
38.2861137390137,24.3085632324219,
44.3944587707520,-11.3621044158936,
0.580600261688232,-35.2464599609375,
-48.4574737548828,-9.26966667175293,
-49.5365982055664,29.7049007415772,
-2.90711307525635,26.1275997161865,
33.7244415283203,-16.1868457794189,
17.7424545288086,-40.7953872680664,
-25.4195346832275,-19.0176277160645,
-39.5726394653320,21.0309867858887,
-14.6004247665405,41.5409393310547,
3.48011350631714,37.6811065673828,
-13.5673961639404,22.9388542175293,
-41.0766639709473,1.18313741683960,
-39.9234619140625,-25.0212726593018,
-11.9350290298462,-38.6912727355957,
10.6037206649780,-37.5980491638184,
14.9564704895020,-40.1575202941895,
19.9399356842041,-54.8391876220703,
39.4852027893066,-55.5254402160645,
57.3306121826172,-14.8583641052246,
56.0297660827637,46.0576667785645,
38.6274261474609,76.9607238769531,
21.2889995574951,57.9670562744141,
9.00158500671387,20.8448066711426,
-4.12891054153442,3.51409816741943,
-18.4520492553711,-1.73721706867218,
-25.0076828002930,-17.4836921691895,
-19.7669086456299,-33.8656044006348,
-9.03477096557617,-23.8932628631592,
1.84384965896606,14.6352195739746,
14.1424398422241,46.2628059387207,
20.7426624298096,46.0847511291504,
15.7944879531860,26.1939296722412,
-1.41017723083496,13.1872158050537,
-17.9826927185059,19.0532627105713,
-21.6263732910156,28.9887161254883,
-13.6278429031372,31.7482910156250,
-9.85660171508789,22.6640663146973,
-22.1106700897217,4.06186628341675,
-41.0024108886719,-16.8605651855469,
-43.2226867675781,-26.3987407684326,
-14.1603097915649,-11.8529109954834,
31.4378299713135,11.7533798217773,
51.5751075744629,21.3071613311768,
20.9662532806397,15.5503072738647,
-36.7314033508301,14.9562044143677,
-68.3960647583008,25.2539997100830,
-52.7399406433106,21.8587093353272,
-20.2203235626221,-19.6317138671875,
-7.00431108474731,-77.8580703735352,
-6.16340923309326,-99.9176788330078,
7.61099624633789,-67.1661453247070,
34.6952743530273,-13.9823493957520,
45.6983833312988,10.8646011352539,
30.2334117889404,1.07702994346619,
16.3068542480469,-19.2022132873535,
27.6008663177490,-29.6362915039063,
49.2563056945801,-29.8083000183105,
52.0597305297852,-21.8518333435059,
39.6790466308594,-5.55206060409546,
35.6211357116699,13.7171707153320,
39.5904655456543,18.4088497161865,
29.8345317840576,0.401751518249512,
6.78718948364258,-25.8690319061279,
2.07355594635010,-36.4980621337891,
26.3713893890381,-23.4552021026611,
52.2779464721680,5.79641151428223,
41.6577453613281,37.1605186462402,
0.202260017395020,53.0068626403809,
-34.6702346801758,37.1537933349609,
-43.1099853515625,3.84403038024902,
-31.7464752197266,-17.1240425109863,
-13.5913276672363,-7.38265800476074,
11.6244182586670,13.5248546600342,
32.6112442016602,9.01459407806397,
25.6976566314697,-21.5543289184570,
-8.51901531219482,-40.3396377563477,
-36.8817291259766,-29.6902160644531,
-36.0026588439941,-16.7322444915772,
-19.0668334960938,-31.6558418273926,
-14.7124681472778,-53.6104927062988,
-30.9472942352295,-39.6355247497559,
-43.2671394348145,6.25730895996094,
-27.6045742034912,31.9176692962647,
10.2630729675293,3.74181842803955,
41.3475227355957,-41.5458869934082,
44.0642509460449,-47.5012474060059,
8.89633941650391,-17.6837768554688,
-39.2568244934082,1.25187659263611,
-48.1284294128418,-16.7896499633789,
0.727260351181030,-39.2972831726074,
59.7442932128906,-28.2508182525635,
58.2243041992188,5.15381050109863,
-6.42410135269165,24.5703582763672,
-53.7179679870606,18.9521007537842,
-26.2447586059570,7.29267454147339,
32.1135368347168,5.65342569351196,
32.7694740295410,4.78987026214600,
-24.5938873291016,-8.07321453094482,
-50.9169883728027,-27.3086719512939,
8.54994392395020,-28.0667381286621,
86.6952743530273,2.89674258232117,
87.6276321411133,46.8439216613770,
11.0442905426025,67.3836212158203,
-52.9148750305176,48.1240043640137,
-43.6537666320801,5.33320808410645,
0.266660332679749,-18.8777065277100,
11.9362268447876,-2.50428295135498,
-10.3466091156006,26.7192115783691,
-22.8641490936279,31.9746513366699,
-7.33751344680786,14.9037466049194,
7.43901634216309,1.77395200729370,
-5.04552698135376,1.87590444087982,
-28.2973098754883,1.29927909374237,
-34.7154960632324,-5.76734018325806,
-30.4692916870117,-0.805100381374359,
-30.5898532867432,18.6624832153320,
-34.2402572631836,15.1021366119385,
-25.3849124908447,-33.6154975891113,
-5.89429569244385,-83.6421737670898,
0.921897828578949,-70.2232589721680,
-19.6841926574707,-7.44652986526489,
-42.1393051147461,23.9474315643311,
-34.1073493957520,-17.5919628143311,
-0.553272962570190,-71.8332748413086,
27.5165786743164,-60.3696479797363,
28.4419918060303,1.04970455169678,
10.1572093963623,31.9756793975830,
-3.44223022460938,0.236305117607117,
4.51842355728149,-42.2117919921875,
33.2919044494629,-38.9746932983398,
64.8162307739258,0.696115732192993,
76.5182723999023,29.5952663421631,
58.5349693298340,34.1677398681641,
23.4906654357910,38.0060043334961,
-4.21184825897217,48.8123474121094,
-10.6534729003906,46.2552986145020,
-5.02529239654541,23.6090583801270,
1.24106907844543,4.79284906387329,
7.00441884994507,7.86409950256348,
12.7780714035034,31.6987724304199,
11.0158348083496,55.0059051513672,
4.10728883743286,55.7738380432129,
-2.16280198097229,33.5248718261719,
-5.24280405044556,7.25576210021973,
-11.4410266876221,-0.841269850730896,
-19.8435344696045,21.2068557739258,
-12.1928787231445,44.5760383605957,
19.7216148376465,29.2542076110840,
48.0296401977539,-17.5587329864502,
39.5446777343750,-36.6149864196777,
0.403678894042969,-0.0616161823272705,
-21.3452224731445,43.3744659423828,
-4.10370349884033,27.7338199615479,
14.3953151702881,-32.3230476379395,
-6.62401390075684,-55.8323554992676,
-51.5302619934082,-13.0215721130371,
-68.4861984252930,24.1910400390625,
-40.3283500671387,-12.5171298980713,
0.603736817836762,-81.0225677490234,
18.9375000000000,-77.4388275146484,
15.0258493423462,15.3126802444458,
7.87870550155640,96.5192871093750,
4.05414867401123,82.4496459960938,
1.13328599929810,10.5403556823730,
2.59418010711670,-24.0226764678955,
6.16395044326782,5.41498661041260,
1.96397960186005,33.4217567443848,
-15.2014045715332,6.09264945983887,
-25.6825542449951,-49.9669837951660,
-15.5822448730469,-71.3946380615234,
-5.56614828109741,-37.8089523315430,
-14.8108987808228,10.4372901916504,
-25.4629230499268,27.8143596649170,
-2.60002088546753,11.8667736053467,
47.1909790039063,-11.0733919143677,
74.2271347045898,-5.87399816513062,
46.3823966979981,35.8967819213867,
-3.31638646125793,80.9979019165039,
-21.1567535400391,78.6809692382813,
-3.27676916122437,23.0296401977539,
14.7806196212769,-38.0445861816406,
21.2312297821045,-53.9308547973633,
27.1830673217773,-22.8823699951172,
30.5189609527588,10.9605550765991,
9.62324523925781,18.2777976989746,
-34.1459121704102,12.3631467819214,
-58.2938919067383,7.05680370330811,
-38.0560913085938,-8.97752380371094,
1.09778523445129,-40.8865737915039,
16.5014400482178,-63.4943122863770,
11.5266323089600,-49.8835487365723,
15.0130805969238,-17.5449695587158,
27.9447040557861,-5.26827621459961,
21.3709716796875,-19.4459991455078,
-10.8588705062866,-26.7416419982910,
-19.4277782440186,-4.47569751739502,
23.2170314788818,23.2571926116943,
78.7103271484375,28.9813728332520,
85.7932891845703,12.6144227981567,
33.3186416625977,-0.355303347110748,
-26.5128326416016,0.511325716972351,
-47.4530067443848,8.16593360900879,
-36.1932334899902,19.8059463500977,
-28.3343753814697,33.9801559448242,
-39.7119636535645,32.7941017150879,
-53.5040931701660,-0.00750690698623657,
-47.5870552062988,-45.4515304565430,
-14.5370855331421,-60.4136581420898,
34.4099044799805,-30.8929824829102,
69.3175277709961,11.1915779113770,
61.2680282592773,20.1426239013672,
12.7508516311646,-4.11873626708984,
-33.1618957519531,-28.6111564636230,
-33.6242828369141,-31.1621303558350,
7.20937061309814,-23.9116458892822,
44.0754127502441,-20.8854064941406,
42.8486480712891,-24.3719196319580,
12.7246770858765,-30.8359127044678,
-6.84861612319946,-39.6710472106934,
1.05466032028198,-42.3672485351563,
20.0868587493897,-26.5754146575928,
28.4215373992920,9.08666133880615,
23.3270950317383,35.6540031433106,
11.2633857727051,23.3776550292969,
2.74161434173584,-18.9787406921387,
-1.48473346233368,-55.2184677124023,
-5.00886726379395,-52.3070755004883,
-9.13204002380371,-20.0346546173096,
-13.9338493347168,14.5333509445190,
-11.4994831085205,39.7588920593262,
-3.60448074340820,58.8630790710449,
0.570452630519867,68.8321304321289,
-4.23782444000244,61.2709655761719,
-9.34057617187500,36.7095451354981,
-0.203566938638687,20.7369689941406,
20.3893642425537,30.4562377929688,
24.8674640655518,52.6931228637695,
-1.02836501598358,51.5528450012207,
-34.8892211914063,10.0154113769531,
-41.8228607177734,-47.8477783203125,
-14.3823480606079,-79.5209808349609,
20.1106700897217,-69.5436096191406,
34.6865615844727,-34.5251655578613,
29.4923915863037,-2.95800852775574,
16.8301906585693,5.30361175537109,
3.57130837440491,-0.662567138671875,
-11.8445968627930,-4.79968833923340,
-22.4874687194824,1.80827224254608,
-18.0186824798584,18.5219726562500,
-5.71600198745728,36.7316856384277,
-0.837527394294739,50.0014953613281,
-8.82645034790039,47.4731369018555,
-15.0139617919922,26.4767360687256,
-7.63441801071167,-1.57991003990173,
2.87864398956299,-11.4620351791382,
2.94874095916748,12.0700626373291,
-6.62364578247070,42.1614646911621,
-14.4694833755493,35.3589439392090,
-18.9930572509766,-12.0690212249756,
-33.0996589660645,-56.8962020874023,
-49.4827384948731,-53.5203170776367,
-39.1987228393555,-14.6535968780518,
5.98569250106812,18.0740871429443,
50.4625129699707,31.2214412689209,
47.6833839416504,42.3767051696777,
-2.04143285751343,57.5479202270508,
-48.3342437744141,54.8903617858887,
-52.4488983154297,23.8576717376709,
-24.8295631408691,-4.95689487457275,
1.44967663288116,2.18828368186951,
18.9927310943604,26.5480384826660,
35.8897171020508,32.2354965209961,
42.7783508300781,14.3724069595337,
17.6538467407227,-0.344295203685761,
-32.0853424072266,-2.16229128837585,
-59.8914718627930,-10.9916057586670,
-38.6306915283203,-29.1540660858154,
2.10834527015686,-24.3380527496338,
11.6187534332275,12.1128387451172,
-9.12110614776611,41.1459999084473,
-20.1050949096680,19.7438468933105,
3.42498779296875,-31.1932640075684,
35.8372688293457,-48.1339149475098,
37.4977378845215,-16.2752246856689,
14.2631788253784,13.6094932556152,
4.68288755416870,-6.06528997421265,
19.7914676666260,-49.6931343078613,
31.8112850189209,-58.1871070861816,
12.3991289138794,-19.1915283203125,
-26.2648468017578,20.7105636596680,
-43.0359268188477,19.2103042602539,
-19.7342948913574,-15.6459894180298,
8.28163719177246,-45.1255035400391,
-3.41691207885742,-45.7527236938477,
-45.5722274780273,-26.3981723785400,
-67.5539703369141,-5.11540365219116,
-40.0197944641113,9.92541599273682,
4.62260818481445,10.9238958358765,
13.1594524383545,-6.47897768020630,
-13.1572017669678,-32.2134780883789,
-24.6278991699219,-44.7795677185059,
4.49210548400879,-29.5393657684326,
34.0030937194824,2.47638440132141,
17.3683605194092,23.1119556427002,
-27.6861972808838,17.9479942321777,
-41.5196266174316,-1.26227211952209,
-5.08030176162720,-7.24178171157837,
37.4633216857910,5.41916751861572,
39.2687454223633,26.4927406311035,
7.17947196960449,36.2757034301758,
-18.5671253204346,23.1020088195801,
-15.3601036071777,-9.07473468780518,
5.95968198776245,-41.6351966857910,
31.4453773498535,-47.1648979187012,
50.0982894897461,-15.8068161010742,
50.7527313232422,32.0165557861328,
25.9567260742188,60.6387176513672,
-5.55395555496216,50.4041366577148,
-13.4237995147705,18.9679431915283,
8.70766162872315,1.44179773330688,
30.2007427215576,11.7754945755005,
22.8461227416992,37.8062438964844,
2.10992646217346,56.8193054199219,
-2.42001914978027,58.2979202270508,
8.91879558563232,50.6891250610352,
7.90417385101318,43.2637252807617,
-20.2634220123291,37.2910614013672,
-45.4265022277832,23.9678745269775,
-33.3695144653320,0.460813701152802,
5.98875522613525,-18.7419586181641,
24.3093109130859,-13.4589109420776,
-3.25367784500122,14.3147048950195,
-46.1121253967285,39.2381477355957,
-54.5207252502441,34.9507217407227,
-20.7441463470459,3.52755188941956,
17.2460842132568,-21.6956729888916,
17.5042209625244,-19.6992549896240,
-18.5889205932617,1.85813653469086,
-48.5314445495606,17.3071308135986,
-42.3726348876953,11.7883987426758,
-8.82049751281738,-13.6624526977539,
19.5452747344971,-41.1758613586426,
24.8344860076904,-53.1673889160156,
21.3681335449219,-40.5651321411133,
27.9983196258545,-17.5120792388916,
40.9282150268555,-6.22143745422363,
30.6314468383789,-12.8667621612549,
-6.39168405532837,-13.0593118667603,
-33.8360252380371,10.9832696914673,
-21.1078567504883,41.6948966979981,
10.6863708496094,41.3928031921387,
13.0684480667114,9.91504478454590,
-27.1309013366699,-8.99863243103027,
-63.2914123535156,9.18366241455078,
-48.2586631774902,30.5209655761719,
1.91757130622864,15.2714900970459,
33.5151214599609,-24.4057502746582,
28.7117824554443,-39.6518402099609,
6.21809625625610,-14.0000629425049,
-14.9348821640015,13.9588537216187,
-36.8957481384277,7.87682390213013,
-56.6015739440918,-16.6737232208252,
-49.1316337585449,-29.5906085968018,
-10.6754102706909,-30.3790168762207,
15.8018474578857,-35.9543380737305,
0.146682977676392,-44.5610923767090,
-26.2481708526611,-39.8401184082031,
-11.6047687530518,-27.2120075225830,
39.0897178649902,-28.6224174499512,
59.9864349365234,-41.1031570434570,
17.4398193359375,-39.3281745910645,
-33.6306838989258,-15.0669822692871,
-20.3830471038818,2.34838652610779,
42.3306045532227,-7.09368133544922,
76.7434005737305,-22.1060123443604,
37.8862113952637,-8.26288795471191,
-33.8496398925781,24.1661491394043,
-64.1224441528320,31.9040603637695,
-28.4468231201172,4.31263732910156,
29.1029930114746,-24.0822620391846,
51.3746452331543,-23.1441898345947,
23.1752758026123,-8.18179798126221,
-21.2420520782471,-7.65520381927490,
-35.5519447326660,-17.4800872802734,
-8.76188087463379,-13.1710147857666,
26.8786487579346,13.1643695831299,
24.4834938049316,36.4766883850098,
-20.3131561279297,39.7730369567871,
-63.7796401977539,29.6726512908936,
-73.6055068969727,21.1457405090332,
-57.4700469970703,10.1947259902954,
-36.6764411926270,-10.3494844436646,
-16.5289001464844,-26.4763278961182,
6.46349954605103,-19.2968826293945,
22.9977855682373,8.65141582489014,
13.9115619659424,34.4714279174805,
-14.7821187973022,38.4836769104004,
-29.9336929321289,25.6762351989746,
-23.6916103363037,9.24692058563232,
-24.9807872772217,-3.74392247200012,
-48.0171775817871,-15.5978279113770,
-63.8047523498535,-25.3587455749512,
-37.2472801208496,-28.7571697235107,
10.8628177642822,-26.3509788513184,
29.7722702026367,-14.9280853271484,
9.79355335235596,6.40769481658936,
-9.67352676391602,27.6120643615723,
-0.792338848114014,27.8775539398193,
16.4868297576904,-0.747028827667236,
11.6793451309204,-31.6126117706299,
-1.82407331466675,-29.8916110992432,
5.74009323120117,7.78619050979614,
26.5382843017578,48.8251762390137,
21.1702175140381,63.3713150024414,
-18.7438087463379,53.1030960083008,
-52.6468391418457,40.7540321350098,
-51.9402732849121,30.3308792114258,
-31.3476200103760,10.4174327850342,
-23.9550952911377,-21.5849914550781,
-23.9964523315430,-51.9201202392578,
-8.71966552734375,-68.1494674682617,
22.8447875976563,-62.2169227600098,
44.3269653320313,-34.7897949218750,
44.4592666625977,3.57010865211487,
44.6538810729981,26.3548488616943,
59.1466598510742,20.6468296051025,
68.0276947021484,2.98795413970947,
50.5927963256836,-3.63957524299622,
23.1882266998291,-1.00188553333282,
10.3866891860962,-12.4888124465942,
10.4851007461548,-41.8502693176270,
-2.67009210586548,-53.7675743103027,
-36.2957687377930,-27.0717506408691,
-63.2582511901856,5.80871391296387,
-59.8995933532715,6.21384334564209,
-35.5267295837402,-14.4202022552490,
-11.5247364044189,-19.5065040588379,
1.49081254005432,-10.4994125366211,
5.38476181030273,-23.9183349609375,
-1.87063765525818,-65.7144927978516,
-16.0267066955566,-77.3405609130859,
-15.2264804840088,-24.7190322875977,
5.86282920837402,49.0366401672363,
22.3395748138428,72.8507614135742,
-0.0616267882287502,38.1204643249512,
-45.0931472778320,9.36424732208252,
-62.8287010192871,21.3434848785400,
-25.6797180175781,42.6356086730957,
30.6211853027344,34.6152534484863,
50.3092193603516,7.69220972061157,
24.3277244567871,1.79583668708801,
-10.0099792480469,21.4462985992432,
-25.9528694152832,39.9816284179688,
-24.7208271026611,29.1091823577881,
-16.1386623382568,-9.09158992767334,
1.89268100261688,-52.2350311279297,
24.6387329101563,-72.4885940551758,
40.4005928039551,-48.0009193420410,
37.1226921081543,8.79227638244629,
14.8839807510376,49.3012466430664,
-17.5376796722412,22.5643711090088,
-47.1591606140137,-50.1665420532227,
-53.5124549865723,-89.9946746826172,
-24.0261230468750,-56.6866798400879,
23.6754798889160,7.63292980194092,
46.4005622863770,36.7901344299316,
21.7150611877441,28.4492168426514,
-12.9258890151978,26.1742687225342,
-13.0083208084106,48.6417388916016,
5.94127893447876,63.5724754333496,
-6.47048950195313,42.5013275146484,
-56.1386871337891,10.3600540161133,
-84.7866134643555,-1.54079198837280,
-52.8045158386231,-6.82701253890991,
5.74050521850586,-29.2978916168213,
30.8621749877930,-59.3750648498535,
20.2560844421387,-64.8739318847656,
23.9807567596436,-43.0066680908203,
56.2850761413574,-25.5802898406982,
74.5699462890625,-25.8030357360840,
52.1974601745606,-28.1998901367188,
17.6023902893066,-25.5169696807861,
11.0327262878418,-29.0177669525147,
22.8426742553711,-36.1979064941406,
20.8015003204346,-19.0102882385254,
5.27447652816773,33.3515090942383,
-0.542521476745606,69.2026290893555,
4.83760261535645,36.9248733520508,
-1.97451198101044,-32.7316474914551,
-25.2038688659668,-59.2439880371094,
-35.3063812255859,-14.9878711700439,
-14.5077896118164,45.8599357604981,
9.02755928039551,61.1949958801270,
3.82856655120850,34.2416687011719,
-20.9106826782227,3.92827844619751,
-35.3527374267578,-9.85547542572022,
-33.9207382202148,-21.0266323089600,
-28.6465167999268,-33.9284629821777,
-16.4066543579102,-42.5875549316406,
6.84621953964233,-49.0745735168457,
28.9400749206543,-62.8294410705566,
23.5531749725342,-65.6303710937500,
-6.55241680145264,-34.9170227050781,
-22.7322673797607,12.9891433715820,
-1.42224717140198,28.7754383087158,
33.2697868347168,-3.88123464584351,
43.4885139465332,-38.8860054016113,
28.3181037902832,-37.1231613159180,
9.71497154235840,-8.06321048736572,
-9.41718578338623,4.85354375839233,
-38.8331451416016,-10.0559482574463,
-60.6425285339356,-21.7508411407471,
-44.1308364868164,-16.2075099945068,
9.26461315155029,-7.44550323486328,
55.7555084228516,-3.61355209350586,
56.8888893127441,10.4765968322754,
28.8320655822754,37.3448982238770,
12.1268367767334,47.3595504760742,
17.2489948272705,23.4637451171875,
24.7878017425537,-10.1898908615112,
23.0415458679199,-18.1627120971680,
22.0734214782715,-9.59362792968750,
23.8392925262451,-18.4099788665772,
17.6340732574463,-46.2576828002930,
11.2045726776123,-56.2984695434570,
22.5522785186768,-26.9654445648193,
51.4474105834961,13.7997331619263,
64.6626052856445,30.5337028503418,
38.5711784362793,26.7981109619141,
-4.27236080169678,26.2575263977051,
-25.6101131439209,23.3689994812012,
-19.0603103637695,0.980816841125488,
-14.9445304870605,-31.6465129852295,
-26.7737655639648,-43.8932800292969,
-31.3856372833252,-27.8592815399170,
-19.1479358673096,-7.15910911560059,
-7.69893789291382,-4.22653055191040,
-11.9610919952393,-13.4274730682373,
-15.7516679763794,-17.1787452697754,
2.62096166610718,-10.8903923034668,
29.7244701385498,1.33244681358337,
32.4582252502441,19.1188125610352,
12.9639625549316,31.4353504180908,
3.52654552459717,12.9250946044922,
14.9410552978516,-30.7428588867188,
18.7710304260254,-53.8874816894531,
-7.16899204254150,-28.4891586303711,
-31.8105831146240,10.8659124374390,
-14.2904958724976,10.5057201385498,
29.9136543273926,-22.0230541229248,
49.1385993957520,-24.9058570861816,
24.6216945648193,21.9792251586914,
-3.43726634979248,66.6117248535156,
5.58642673492432,54.2618446350098,
36.4681053161621,10.8544187545776,
44.8394355773926,-2.27449703216553,
15.4342870712280,15.8467359542847,
-21.5179119110107,14.4888086318970,
-33.4208984375000,-18.8911056518555,
-22.0453281402588,-41.5078430175781,
-5.46940422058106,-24.4585876464844,
3.24456453323364,3.75792598724365,
-1.78901863098145,3.36948633193970,
-17.7453861236572,-22.4794349670410,
-30.4525413513184,-42.3333930969238,
-26.5089130401611,-46.5897521972656,
-10.7810068130493,-43.7135925292969,
2.17316794395447,-25.9926471710205,
2.34905552864075,16.0562019348145,
-13.1884899139404,51.8427200317383,
-36.5549621582031,33.4872474670410,
-59.3617897033691,-26.4161224365234,
-62.7421607971191,-53.1288528442383,
-30.1581821441650,-11.7672348022461,
21.2822265625000,39.6434860229492,
42.4658241271973,27.8786315917969,
12.0112342834473,-28.1969089508057,
-28.3969573974609,-41.7893714904785,
-26.5958957672119,16.6796627044678,
2.60887956619263,75.8216094970703,
4.99997854232788,65.1810913085938,
-25.2647533416748,9.17235374450684,
-34.2339897155762,-18.3428840637207,
11.7370681762695,-1.29936170578003,
68.2285919189453,10.7835655212402,
70.1070632934570,-11.4950389862061,
20.1127490997314,-32.8267707824707,
-23.4878940582275,-16.6351203918457,
-28.4120292663574,14.5037975311279,
-11.7143459320068,18.4737606048584,
7.67842245101929,-3.80611586570740,
27.6941089630127,-9.63928604125977,
39.9076805114746,20.0945167541504,
18.6257553100586,47.1787681579590,
-29.6009559631348,33.2314453125000,
-50.1807823181152,-4.17571735382080,
-12.0329799652100,-19.0210514068604,
51.2686195373535,3.14695620536804,
72.7094116210938,33.4815826416016,
36.2375488281250,39.7379417419434,
-8.17308044433594,24.1461601257324,
-15.4559383392334,10.8905696868896,
3.76846623420715,9.20635604858398,
12.1431350708008,2.45399522781372,
-0.755950808525085,-19.0515975952148,
-18.4446678161621,-37.1590270996094,
-24.2377796173096,-32.3283729553223,
-15.4915075302124,-6.00938606262207,
1.35773050785065,16.6677188873291,
13.0689449310303,16.7275581359863,
6.27205324172974,5.11520338058472,
-22.9420433044434,3.76047897338867,
-53.3346366882324,10.8269720077515,
-55.1486129760742,-0.175188064575195,
-19.9735851287842,-32.1219596862793,
25.5088882446289,-49.3720970153809,
39.1414794921875,-20.7929801940918,
13.1914720535278,34.8883132934570,
-25.1185245513916,54.2133255004883,
-44.1225051879883,9.78859519958496,
-33.2127761840820,-53.1259994506836,
-11.5629014968872,-70.7483596801758,
-3.12985682487488,-34.9189071655273,
-16.2958965301514,4.94578075408936,
-37.2872352600098,13.0179443359375,
-46.9389801025391,0.543001174926758,
-36.3150215148926,-3.60552549362183,
-14.4049339294434,-2.17533659934998,
7.32256841659546,-17.3948230743408,
24.9304523468018,-40.0349807739258,
40.1436576843262,-35.2856941223145,
48.1445770263672,8.99812889099121,
34.5413818359375,54.0545921325684,
-0.772273659706116,56.3534317016602,
-36.4914665222168,15.8221635818481,
-51.2654533386231,-23.6681995391846,
-45.8206062316895,-31.8836097717285,
-35.4423103332520,-21.9176845550537,
-30.9843463897705,-15.7886819839478,
-26.7852611541748,-12.4357261657715,
-18.6430034637451,1.32275307178497,
-11.4729261398315,22.4148464202881,
-6.58150243759155,26.6200122833252,
4.75096368789673,2.60303330421448,
21.8446521759033,-27.6110267639160,
29.8447360992432,-37.5734977722168,
12.7891798019409,-25.8518104553223,
-16.7507324218750,-14.6085567474365,
-31.9927825927734,-16.7728614807129,
-23.7676277160645,-26.1831321716309,
-13.4629783630371,-28.9748458862305,
-17.5436840057373,-21.7964057922363,
-25.3409118652344,-9.47179031372070,
-19.3559169769287,7.04282760620117,
4.39094352722168,25.0092449188232,
24.1744174957275,36.5512847900391,
24.7746810913086,34.2876510620117,
10.1817684173584,22.7209091186523,
-2.09056782722473,9.77470874786377,
-1.45383894443512,-2.64695572853088,
8.88820362091065,-17.7726783752441,
17.5262565612793,-29.2615432739258,
16.6504058837891,-30.1246643066406,
9.99406909942627,-22.2568435668945,
9.15954399108887,-20.6712493896484,
16.6776561737061,-35.5602073669434,
17.6689186096191,-49.8052101135254,
-0.124305009841919,-43.1905403137207,
-31.3764610290527,-14.2047252655029,
-50.3171310424805,19.8799953460693,
-42.7161026000977,43.8790702819824,
-16.6010189056397,54.3049964904785,
7.61449575424194,53.7220001220703,
18.2995510101318,42.7155952453613,
15.7303485870361,29.9052391052246,
3.30816602706909,21.6548881530762,
-13.4750308990479,14.6014642715454,
-24.7102584838867,-3.61718964576721,
-15.7689609527588,-31.7340488433838,
8.67728424072266,-44.4627914428711,
28.4399375915527,-20.2733955383301,
24.3602180480957,24.6989288330078,
-4.40693473815918,50.4429855346680,
-40.6211547851563,43.7057571411133,
-60.8152427673340,24.1038532257080,
-51.6635513305664,14.5287990570068,
-18.9008045196533,16.5647754669189,
11.0814304351807,21.0608139038086,
11.4870901107788,25.1671657562256,
-16.2704696655273,28.8431091308594,
-34.3041534423828,19.3210773468018,
-9.17287158966065,-5.05002307891846,
34.3949508666992,-26.2362232208252,
39.1906738281250,-22.9162120819092,
-10.4042835235596,-6.39187526702881,
-60.0718040466309,-6.71410131454468,
-51.5711898803711,-26.3233184814453,
1.88028788566589,-33.3153724670410,
31.8886470794678,-4.95376777648926,
7.80677700042725,32.3653678894043,
-26.8172302246094,42.6995086669922,
-21.6154136657715,25.1967144012451,
9.40102767944336,4.39471054077148,
23.4069442749023,0.827125787734985,
16.2923030853272,8.27277565002441,
22.1627845764160,14.7009668350220,
45.5265312194824,17.4888420104980,
48.7880439758301,11.4360008239746,
12.8021945953369,-4.20072507858276,
-18.5391101837158,-18.3115005493164,
-3.25066661834717,-13.5956058502197,
33.5895347595215,15.0654602050781,
34.3906669616699,45.2097587585449,
-5.32344388961792,57.1405982971191,
-28.6717548370361,53.6021499633789,
-3.69144701957703,41.9423141479492,
26.0855331420898,19.3427886962891,
10.3449611663818,-12.5860376358032,
-32.2117919921875,-40.9524612426758,
-46.3334007263184,-47.9413261413574,
-22.1557235717773,-26.7823352813721,
-5.15534877777100,7.27663707733154,
-25.6423435211182,35.4445724487305,
-53.7578163146973,38.9189262390137,
-52.0872268676758,6.26904487609863,
-23.5038089752197,-46.8521728515625,
-4.59956216812134,-75.4360504150391,
-7.54377317428589,-46.2471733093262,
-12.5743751525879,14.5048198699951,
-11.5680437088013,40.7325897216797,
-13.6428747177124,9.75805473327637,
-19.6418228149414,-28.0699443817139,
-21.3517990112305,-19.4800529479980,
-11.5909070968628,26.4558773040772,
-1.98434090614319,46.4639358520508,
-5.44510555267334,13.8997001647949,
-17.3184432983398,-32.5678901672363,
-19.2519645690918,-46.9404106140137,
-0.377580642700195,-28.7346439361572,
32.5709342956543,-10.6694374084473,
57.1537857055664,-5.47488069534302,
49.3441734313965,-4.03987598419189,
-1.12282454967499,-0.550701916217804,
-59.4372406005859,-5.69640302658081,
-70.6627655029297,-20.4119739532471,
-18.5761432647705,-21.3939094543457,
46.4271888732910,-2.99976873397827,
58.1496925354004,12.6147766113281,
8.64320564270020,0.701940774917603,
-46.2312583923340,-29.6823825836182,
-53.9023857116699,-42.0130615234375,
-21.8371086120605,-13.4922199249268,
5.87696313858032,28.3236827850342,
5.94221830368042,38.7624893188477,
-11.0642156600952,12.3877143859863,
-31.5872726440430,-15.2621126174927,
-48.5835380554199,-9.92749881744385,
-52.1692924499512,19.2413692474365,
-30.5405387878418,32.3593444824219,
8.48472023010254,4.54449844360352,
30.0307407379150,-35.5000381469727,
16.5333919525147,-45.8366889953613,
-3.40720605850220,-23.3253383636475,
8.89410495758057,-6.86300325393677,
50.9149894714356,-12.1386651992798,
74.8327713012695,-10.6329660415649,
49.1010360717773,22.1392288208008,
2.31546115875244,60.5398635864258,
-19.9320659637451,53.6093864440918,
-15.0359401702881,2.23644137382507,
-13.7041397094727,-32.4360580444336,
-31.4946689605713,-16.1493759155273,
-46.8925476074219,9.04705524444580,
-38.6105041503906,-10.0629224777222,
-14.7543811798096,-59.0376091003418,
5.27578067779541,-77.0368576049805,
13.2802753448486,-50.0286331176758,
15.7053432464600,-27.5748214721680,
12.8872365951538,-42.2545166015625,
1.43572449684143,-52.8838653564453,
-8.91621971130371,-16.5342254638672,
-11.2796220779419,45.6332283020020,
-15.0590772628784,67.0620498657227,
-33.4717292785645,27.6702060699463,
-53.6767578125000,-22.0998878479004,
-55.7864570617676,-33.6485939025879,
-32.5689735412598,-14.2183399200439,
-1.07915735244751,1.35022163391113,
20.4794063568115,3.22500896453857,
27.2603588104248,4.08217763900757,
20.2507133483887,5.67772102355957,
-0.993671178817749,-2.09979414939880,
-24.3460350036621,-21.0603027343750,
-21.9401168823242,-43.5563468933106,
7.72812843322754,-59.2545852661133,
32.6989479064941,-66.4054260253906,
25.6400604248047,-58.9864921569824,
6.15242576599121,-28.2543125152588,
10.9866437911987,15.0550603866577,
37.8734092712402,39.0373840332031,
51.9556121826172,31.2441768646240,
37.2522926330566,17.4148311614990,
15.5949096679688,22.3525753021240,
5.69095516204834,39.6047477722168,
-3.52940368652344,42.8443145751953,
-28.5643711090088,23.5651245117188,
-47.7718505859375,5.84045743942261,
-31.8336830139160,2.07958650588989,
10.8419618606567,-0.245860248804092,
42.3845634460449,-8.52237701416016,
44.8526039123535,-4.80338907241821,
31.8554668426514,25.6679801940918,
13.9826879501343,56.3713912963867,
-7.83766269683838,48.8296318054199,
-23.4671173095703,3.09610319137573,
-17.8845634460449,-31.0281486511230,
6.48580789566040,-25.4797706604004,
15.1169643402100,-8.74182033538818,
-10.2072000503540,-15.2092618942261,
-38.5756111145020,-36.3524322509766,
-27.4388885498047,-28.7956008911133,
11.6289024353027,18.9997558593750,
32.3725090026856,64.2457199096680,
20.1611347198486,60.3396682739258,
11.5100135803223,17.7424621582031,
26.6085243225098,-16.5667610168457,
34.0930252075195,-12.4314527511597,
1.88467049598694,11.1593513488770,
-41.5981712341309,16.8359966278076,
-34.4500808715820,-7.89956665039063,
25.7420215606689,-30.9412841796875,
72.0742568969727,-13.7836942672730,
50.7077484130859,33.7039031982422,
-10.4905357360840,62.2064933776856,
-39.2605056762695,40.9856567382813,
-10.8584260940552,-2.99464702606201,
32.5240516662598,-18.8600883483887,
43.4140167236328,3.23197460174561,
22.2820587158203,22.9983043670654,
-8.07899665832520,7.35840034484863,
-32.2394180297852,-20.0075740814209,
-50.3534622192383,-23.0866012573242,
-57.9515914916992,-10.9540452957153,
-38.5250549316406,-16.4870414733887,
4.69177770614624,-44.2807197570801,
41.5625228881836,-55.5125923156738,
43.3685035705566,-29.6732788085938,
15.6787090301514,6.20448589324951,
-11.0868730545044,15.4051694869995,
-16.2857685089111,7.67606067657471,
-3.35564947128296,12.9038677215576,
-1.11393857002258,31.4991817474365,
-22.4243488311768,32.7630119323731,
-42.6115379333496,2.99613952636719,
-28.2518901824951,-22.6464366912842,
16.6779136657715,-10.0171165466309,
49.3846397399902,26.2613716125488,
32.0309066772461,44.4018135070801,
-17.3469963073730,26.8323764801025,
-40.2770423889160,-9.21292114257813,
-16.8344535827637,-39.7513427734375,
16.7205066680908,-52.8448944091797,
18.3751964569092,-51.4753608703613,
5.32667922973633,-42.6042861938477,
16.9152526855469,-36.9993705749512,
45.8013496398926,-41.9452781677246,
45.7939987182617,-45.4870071411133,
7.81643676757813,-24.8132839202881,
-17.4812564849854,16.0739536285400,
7.46629905700684,39.0600929260254,
43.9846763610840,19.2743206024170,
30.1286983489990,-20.4823722839355,
-26.7084751129150,-42.5007629394531,
-59.6395530700684,-41.2298240661621,
-30.2248649597168,-34.2797470092773,
24.8766746520996,-27.0598087310791,
50.1081809997559,-3.99286055564880,
41.0266151428223,29.6393547058105,
24.2527751922607,35.9158630371094,
8.95869445800781,1.04565644264221,
-9.23060417175293,-34.2612152099609,
-23.7536659240723,-27.3512020111084,
-15.7061052322388,4.11893510818481,
13.4157781600952,10.7984189987183,
37.4630279541016,-20.4428329467773,
35.3419952392578,-44.3827056884766,
14.9182567596436,-30.1273727416992,
-5.31834602355957,-5.09230375289917,
-19.0890598297119,-5.36413669586182,
-26.2910690307617,-19.9372978210449,
-21.2067527770996,-9.27865123748779,
-8.95867919921875,32.2814178466797,
-6.94901609420776,59.6423645019531,
-19.3808555603027,38.1504402160645,
-27.8523616790772,-8.87663173675537,
-9.19222640991211,-32.3242607116699,
27.6344356536865,-20.4579944610596,
44.7059097290039,-7.93856668472290,
25.6551017761230,-23.0270500183105,
-6.42368841171265,-50.4567222595215,
-17.0772438049316,-49.1478576660156,
-6.25766181945801,-7.20895576477051,
-0.311697781085968,34.7634696960449,
-8.60460758209229,28.3992328643799,
-11.2167787551880,-13.4681797027588,
9.39165210723877,-38.1176719665527,
33.3023910522461,-12.3321399688721,
27.3275775909424,30.8516941070557,
-5.39652538299561,34.1709671020508,
-25.9500923156738,-9.29092693328857,
-5.11260032653809,-48.0607948303223,
33.1588706970215,-39.2042160034180,
42.8310317993164,-3.67871189117432,
12.3978166580200,12.0521907806396,
-22.6388835906982,-3.27863407135010,
-30.6346359252930,-17.2893562316895,
-19.4561729431152,-9.62022590637207,
-14.9272127151489,-2.65002322196960,
-21.7692680358887,-27.1939888000488,
-18.0487422943115,-70.7963638305664,
6.65779399871826,-86.7726593017578,
27.9508323669434,-57.7339744567871,
17.5807838439941,-8.27651691436768,
-15.4884262084961,20.4765911102295,
-36.5951843261719,20.2283477783203,
-21.8218498229980,16.4674358367920,
12.7186450958252,25.7311820983887,
30.3713226318359,35.0680313110352,
18.4522895812988,24.4813098907471,
-1.17822825908661,-3.79708075523376,
-2.71181464195251,-29.6541061401367,
10.0109910964966,-36.1204948425293,
16.1048355102539,-26.0568981170654,
7.57834959030151,-12.3336534500122,
1.26852941513062,3.08715796470642,
13.9464874267578,30.3251571655273,
32.6407279968262,64.4223785400391,
23.4287414550781,85.2103347778320,
-21.3213481903076,75.9964599609375,
-68.9912338256836,36.1852416992188,
-76.5771255493164,-5.23091554641724,
-38.0111694335938,-26.5331764221191,
9.55338668823242,-26.2516269683838,
23.9323043823242,-18.8024787902832,
-0.531655192375183,-12.1754817962646,
-36.4415054321289,-5.74139499664307,
-50.3798217773438,-2.43343305587769,
-33.1484870910645,-9.09031105041504,
-2.90901207923889,-23.7504119873047,
15.8884773254395,-25.8418617248535,
12.9270410537720,6.28783988952637,
-0.910936713218689,57.4747657775879,
-12.5012063980103,80.7261962890625,
-20.1280651092529,45.4020500183106,
-29.1038627624512,-19.0047378540039,
-36.4409942626953,-61.0280799865723,
-28.1811275482178,-59.8615264892578,
-4.57267761230469,-47.1285972595215,
7.31921958923340,-49.8941535949707,
-8.80440139770508,-52.7644309997559,
-34.1601104736328,-29.2652206420898,
-35.1669197082520,16.4372844696045,
-5.93948745727539,49.5047035217285,
21.6465644836426,51.2223701477051,
16.6274776458740,38.1774635314941,
-7.86395120620728,25.9377231597900,
-23.8366336822510,11.0282211303711,
-23.2954158782959,-6.59605407714844,
-16.4188156127930,-10.8108243942261,
-7.85451698303223,6.39232254028320,
5.41882228851318,27.2833633422852,
12.2504138946533,30.1037197113037,
1.87737202644348,14.3595418930054,
-11.4228887557983,-7.12059926986694,
2.82882332801819,-25.3087482452393,
42.0811042785645,-39.5189094543457,
59.5677757263184,-33.6055145263672,
23.2469272613525,4.65862035751343,
-26.4046936035156,47.7355499267578,
-29.0846920013428,47.0980262756348,
17.6853828430176,4.22281265258789,
49.1456718444824,-26.5488033294678,
23.4921913146973,-13.5295734405518,
-22.6519241333008,9.54519939422607,
-33.9085884094238,-3.61069703102112,
-13.1892738342285,-38.8164176940918,
-3.23767948150635,-42.9201354980469,
-17.0538444519043,-12.1431255340576,
-21.5687484741211,3.23991799354553,
6.31704092025757,-20.0033397674561,
36.8923492431641,-35.5252990722656,
24.9048709869385,1.48128342628479,
-29.1749534606934,57.4028816223145,
-77.8523788452148,61.4335212707520,
-79.5057678222656,4.79160547256470,
-40.2164268493652,-50.1335487365723,
4.19445943832398,-51.0987205505371,
23.4133262634277,-18.0970859527588,
15.4376125335693,5.82769393920898,
3.81093144416809,10.7472333908081,
9.52586460113525,21.1177406311035,
22.7725429534912,44.2429161071777,
17.7063140869141,56.8791656494141,
-9.83946228027344,43.1468963623047,
-36.5181808471680,14.0849208831787,
-36.6789093017578,-6.67491102218628,
-13.4812355041504,-14.8253593444824,
3.61884498596191,-12.3412122726440,
3.07239580154419,4.18614435195923,
-3.81426906585693,33.7232093811035,
-5.08935832977295,60.9351119995117,
-3.95648908615112,67.9837570190430,
-2.13777518272400,51.7247886657715,
2.52614593505859,33.1098861694336,
12.9372901916504,26.7784881591797,
16.3527221679688,20.4780750274658,
7.20072841644287,1.78377127647400,
2.47150087356567,-19.3922176361084,
14.9097690582275,-18.6121654510498,
34.2923622131348,10.9474830627441,
31.6992321014404,42.5206146240234,
-0.510511875152588,49.9271736145020,
-42.5131187438965,29.9067440032959,
-68.6257781982422,5.29290485382080,
-69.1389160156250,-7.08071231842041,
-46.8033256530762,-7.92840528488159,
-12.3972835540771,-0.564985573291779,
12.5362272262573,12.6337566375732,
5.20355558395386,25.6849689483643,
-27.1975421905518,20.5000133514404,
-44.1898765563965,-0.155163526535034,
-15.8711395263672,-15.8853931427002,
32.1992225646973,-2.69483923912048,
47.7468528747559,34.1006317138672,
13.6053218841553,58.8541374206543,
-33.6444740295410,46.1783370971680,
-48.0274353027344,4.45230579376221,
-27.2220630645752,-31.7657794952393,
-5.16333055496216,-35.8253250122070,
-6.62332677841187,-11.3923978805542,
-23.6403598785400,18.7069473266602,
-38.1599235534668,31.0586891174316,
-37.9723739624023,24.4289054870605,
-22.5442352294922,21.4175739288330,
-2.89379668235779,39.0286178588867,
1.71903276443481,61.5781974792481,
-16.5248699188232,54.5547561645508,
-38.9097785949707,8.85122489929199,
-38.5067367553711,-49.8376770019531,
-16.8604316711426,-79.4154663085938,
-4.47816705703735,-62.5698928833008,
-18.5556793212891,-17.8279094696045,
-34.7840690612793,17.8955421447754,
-16.6995201110840,20.2280845642090,
20.1765861511230,-10.4157085418701,
25.0572280883789,-38.4272613525391,
-9.71717453002930,-26.7552928924561,
-38.1284065246582,20.7511291503906,
-22.4191322326660,54.4530410766602,
11.0688438415527,34.4106063842773,
15.2460660934448,-9.54253768920898,
-6.75525665283203,-16.0176048278809,
-10.7496633529663,24.7348861694336,
12.8505487442017,59.2503433227539,
23.8235893249512,49.9370536804199,
7.80615949630737,16.8485660552979,
-0.763953506946564,4.31796264648438,
26.6626300811768,17.9399394989014,
49.7251739501953,23.1170024871826,
21.9795475006104,11.6839761734009,
-30.2620391845703,-3.18460941314697,
-37.7542495727539,-16.8818073272705,
10.2916755676270,-35.0881195068359,
49.4626960754395,-42.3948478698731,
31.2837352752686,-12.4383678436279,
-8.77354907989502,38.9021949768066,
-13.9533233642578,54.8330116271973,
12.0720186233521,16.7365283966064,
14.9354486465454,-21.0971717834473,
-19.5583248138428,-7.34988021850586,
-56.2632446289063,32.7929344177246,
-65.7108688354492,33.6229896545410,
-59.5085296630859,-18.9828224182129,
-50.9253883361816,-63.4252395629883,
-29.1305122375488,-59.1132011413574,
10.2200260162354,-32.6899375915527,
42.6266822814941,-26.5820159912109,
42.9982261657715,-35.7537460327148,
21.8750820159912,-31.6339073181152,
14.1505517959595,-16.1998138427734,
31.9723281860352,-11.0023775100708,
46.8525657653809,-16.3373088836670,
42.6951866149902,-10.7191877365112,
34.0107688903809,6.54917430877686,
36.6189231872559,16.7820816040039,
46.8439178466797,9.90956687927246,
52.0060043334961,6.52614927291870,
44.6483345031738,21.2058029174805,
19.1965122222900,40.1294174194336,
-15.8137865066528,41.1863937377930,
-45.3858528137207,26.6019191741943,
-42.5865097045898,9.78282070159912,
-10.8042421340942,-11.7663316726685,
8.53113842010498,-34.7111740112305,
-16.4708843231201,-42.0842933654785,
-56.2981033325195,-23.6804485321045,
-48.3281822204590,-3.03810143470764,
11.1627521514893,-3.03303956985474,
58.4793434143066,-13.8734226226807,
44.1823577880859,2.42246580123901,
-1.03659534454346,48.7500915527344,
-17.9922847747803,85.5452804565430,
-4.12859678268433,81.3183593750000,
-14.1671009063721,50.6908607482910,
-64.4900207519531,24.6604213714600,
-98.1537933349609,4.17338848114014,
-66.8325042724609,-21.5670719146729,
-2.42382812500000,-34.5929107666016,
27.3103237152100,-16.3536396026611,
6.27826309204102,12.9263544082642,
-9.42088508605957,11.4028053283691,
15.2405452728271,-22.8247756958008,
49.7474327087402,-44.3455276489258,
50.2242965698242,-21.0412559509277,
24.3316287994385,25.5603637695313,
11.7598390579224,52.4005470275879,
20.6056747436523,48.2074279785156,
21.6995449066162,28.7976722717285,
-3.86420154571533,3.17649936676025,
-24.4562950134277,-23.3660163879395,
-10.5953149795532,-33.2308959960938,
18.8140201568604,-10.4054031372070,
19.9335746765137,24.4309196472168,
-15.6197071075439,30.1612434387207,
-57.0958442687988,1.34728169441223,
-66.6540451049805,-18.4432086944580,
-43.8341674804688,0.0331690311431885,
-11.7835674285889,35.4092063903809,
16.4611072540283,46.8182411193848,
37.9443168640137,25.2872714996338,
44.3745193481445,1.34642803668976,
24.4734134674072,0.0205167233943939,
-14.0826282501221,6.60711860656738,
-51.4024734497070,-2.03857135772705,
-65.2956237792969,-21.8189163208008,
-52.0475082397461,-30.7966060638428,
-22.8428211212158,-11.2408208847046,
5.06290912628174,24.8229789733887,
11.9231815338135,43.6803398132324,
-5.03915786743164,23.1060867309570,
-28.7180652618408,-23.5485630035400,
-33.4988250732422,-48.0140075683594,
-11.6916952133179,-24.4387321472168,
11.4554347991943,24.1711616516113,
12.3924140930176,46.0738258361816,
-3.89540386199951,18.5308570861816,
-7.39554309844971,-25.7649555206299,
15.9657173156738,-39.1428070068359,
40.4456710815430,-22.6519851684570,
35.5694656372070,-11.8666553497314,
1.28872644901276,-23.7482566833496,
-24.6493511199951,-35.6508216857910,
-7.09209823608398,-20.4939804077148,
40.1487121582031,9.09154033660889,
70.2001495361328,22.0439281463623,
50.2614669799805,15.3596200942993,
2.65454387664795,20.6844387054443,
-26.3161201477051,48.2152709960938,
-19.7768802642822,64.2501068115234,
-0.653835594654083,36.6960983276367,
4.37515926361084,-14.1409187316895,
0.0978554785251617,-31.1466865539551,
9.85796737670898,4.18315124511719,
30.2752590179443,43.3087005615234,
40.5710449218750,38.5715675354004,
37.3757400512695,4.06263446807861,
36.9088516235352,-8.92766380310059,
45.6009063720703,17.4957294464111,
44.1275939941406,42.6624488830566,
20.3229408264160,33.3347930908203,
-2.52097773551941,6.82243156433106,
0.403484821319580,2.49104118347168,
17.5434608459473,24.1432285308838,
16.4738044738770,38.6797142028809,
-5.42419052124023,27.0134601593018,
-15.0631847381592,4.85326147079468,
11.0969524383545,-7.19554424285889,
51.0042037963867,-6.06723594665527,
64.3732681274414,-0.886071681976318,
39.5153503417969,7.06734275817871,
-7.85463809967041,14.4071350097656,
-51.8342895507813,7.45337104797363,
-72.8378829956055,-20.9353637695313,
-58.9502029418945,-47.5358238220215,
-27.0925045013428,-43.7657661437988,
-11.5415315628052,-16.2413024902344,
-31.3797206878662,-0.892996609210968,
-54.1006355285645,-15.0429811477661,
-38.3864173889160,-35.8070602416992,
15.5952091217041,-30.5822525024414,
51.3857002258301,-1.32413482666016,
34.1535415649414,23.9320678710938,
-3.64419889450073,23.9599514007568,
-8.26638603210449,12.6272048950195,
21.9534969329834,13.0351982116699,
45.1005706787109,27.6767578125000,
38.9900856018066,35.3965911865234,
23.2120018005371,19.5610599517822,
24.6105842590332,-14.3981304168701,
34.7042121887207,-33.6243476867676,
33.2460365295410,-12.9531478881836,
24.8316688537598,32.5593948364258,
20.6664676666260,62.9698143005371,
8.17725658416748,63.1795234680176,
-33.5199737548828,47.1367607116699,
-86.5707321166992,27.9209022521973,
-99.0872573852539,-0.579429149627686,
-49.8678970336914,-42.0746917724609,
11.2432518005371,-65.6321868896484,
21.2518424987793,-36.6512451171875,
-15.8613777160645,18.3254127502441,
-42.0232124328613,29.5741939544678,
-23.0501785278320,-24.8026733398438,
16.5342044830322,-82.4873504638672,
33.5018043518066,-72.9102935791016,
27.4582252502441,-11.6644134521484,
27.2866554260254,25.3609752655029,
44.9322547912598,2.86429524421692,
57.7726135253906,-29.7772636413574,
47.8900756835938,-21.2207832336426,
25.2221069335938,7.60667181015015,
10.0647869110107,1.39829277992249,
4.33339977264404,-43.8253402709961,
-4.49808216094971,-71.7024612426758,
-17.0767192840576,-43.8975715637207,
-21.7726573944092,9.58846282958984,
-3.74895215034485,30.7779769897461,
22.7117385864258,9.29981231689453,
31.5077419281006,-15.9135990142822,
16.4274692535400,-22.5915813446045,
-2.13941812515259,-29.3835048675537,
-0.995589315891266,-51.1445922851563,
14.2173862457275,-66.7347793579102,
15.4795417785645,-43.7757949829102,
-6.75701951980591,1.45999586582184,
-29.1940937042236,12.8622636795044,
-26.9672660827637,-27.1788978576660,
-6.99042081832886,-63.5444793701172,
9.46778392791748,-41.1820869445801,
10.6778478622437,19.5754547119141,
9.35716342926025,46.6786842346191,
16.3328151702881,14.1342411041260,
23.9019298553467,-32.4826431274414,
22.1328105926514,-38.6178512573242,
10.5940923690796,-17.8761615753174,
-0.734993934631348,-14.9981355667114,
-3.24230504035950,-31.9394931793213,
0.509265959262848,-28.5937900543213,
2.03819966316223,9.52454280853272,
-10.1149606704712,40.3861694335938,
-32.7474441528320,29.1267299652100,
-42.8587303161621,-8.61360836029053,
-20.5607566833496,-26.9583568572998,
22.2262744903564,-16.3878211975098,
46.7598457336426,-10.8816318511963,
27.7126750946045,-27.0336208343506,
-11.3675012588501,-39.4650115966797,
-24.6960144042969,-22.5202407836914,
-0.170328378677368,10.4305553436279,
31.2204074859619,26.2264862060547,
33.0482025146484,16.2978382110596,
0.623302936553955,6.01322221755981,
-38.6235389709473,14.6063842773438,
-57.1790542602539,23.6790866851807,
-50.6389579772949,5.21549463272095,
-29.2173442840576,-31.3897418975830,
-5.20183849334717,-46.2081947326660,
9.31045722961426,-19.8167610168457,
5.85161209106445,23.2116851806641,
-9.16276073455811,46.2126998901367,
-18.5228939056397,45.6219711303711,
-4.32795715332031,42.5646743774414,
25.6827507019043,39.2862968444824,
40.3057022094727,19.5426769256592,
24.5826473236084,-16.6666908264160,
4.28517436981201,-32.5014495849609,
14.7257204055786,-6.85583019256592,
44.3715858459473,27.8998336791992,
48.4514312744141,23.1614151000977,
11.4902133941650,-18.7061138153076,
-20.9422473907471,-44.6137619018555,
-9.43184280395508,-27.3704071044922,
22.7921752929688,2.38013863563538,
20.1616420745850,6.87003898620606,
-16.6615772247314,-4.51248741149902,
-36.3817901611328,-4.67391729354858,
-17.5590934753418,5.97712135314941,
-1.77458000183105,-1.89365053176880,
-18.3599414825439,-32.2396926879883,
-33.1265296936035,-48.8711013793945,
-2.32025337219238,-30.4610939025879,
50.2249145507813,4.98685789108276,
58.3298530578613,28.7116985321045,
13.5935726165771,35.0663642883301,
-27.7997303009033,30.9094448089600,
-27.1998329162598,13.3941516876221,
-12.3950843811035,-12.7462949752808,
-24.1312999725342,-23.6369190216064,
-53.3463859558106,-4.68894100189209,
-59.0079078674316,16.3969364166260,
-37.1053123474121,3.01707530021668,
-21.7799415588379,-42.1670379638672,
-27.4157810211182,-67.4482421875000,
-34.0700683593750,-42.1361236572266,
-23.1535320281982,2.35931634902954,
-0.340327024459839,15.8665819168091,
18.3412151336670,-7.78828620910645,
26.7010021209717,-28.4487953186035,
24.8547058105469,-21.2477378845215,
12.7982606887817,3.74085950851440,
0.424340546131134,20.5501594543457,
2.30339789390564,22.2267570495605,
22.8925514221191,17.2179832458496,
35.1896705627441,17.7550220489502,
13.0411615371704,25.8334751129150,
-23.8376522064209,37.4775352478027,
-31.5128936767578,44.9699134826660,
0.376791477203369,44.5265846252441,
32.9933547973633,33.9844589233398,
29.4728202819824,18.0507335662842,
4.70009040832520,-0.244354113936424,
-5.60318756103516,-22.7359352111816,
8.84652423858643,-39.7342300415039,
24.3694286346436,-37.4549674987793,
26.9964790344238,-24.5465908050537,
29.5044136047363,-23.6351909637451,
42.8946914672852,-33.6098060607910,
50.1588211059570,-23.0006141662598,
33.5162239074707,26.0048217773438,
6.80443191528320,79.6778717041016,
-3.06148576736450,83.9758605957031,
6.24821662902832,39.9127464294434,
10.9633769989014,8.94492626190186,
-3.54217362403870,28.2203865051270,
-31.9119720458984,57.7382049560547,
-53.4120864868164,44.0266189575195,
-54.1552619934082,0.373792529106140,
-33.6809387207031,-10.9158430099487,
-4.56175184249878,21.5381431579590,
5.76431608200073,43.6645355224609,
-18.3524589538574,17.1883201599121,
-55.1891288757324,-16.6236610412598,
-59.5121002197266,-6.83433151245117,
-24.2536277770996,30.8359737396240,
10.1021642684937,34.0087585449219,
9.34173679351807,-10.4282274246216,
-5.58185386657715,-45.9523773193359,
-2.40336084365845,-28.2663822174072,
9.93913841247559,15.5330390930176,
-5.61755275726318,30.4056568145752,
-49.0551872253418,12.4824237823486,
-71.3802108764648,-6.75626850128174,
-40.7692070007324,-9.85804748535156,
8.24182510375977,-8.46029090881348,
27.2608699798584,-16.9452171325684,
19.4172248840332,-32.2983741760254,
19.1904354095459,-42.7737159729004,
30.4427623748779,-42.7159233093262,
27.5065193176270,-26.9080638885498,
6.38106060028076,4.48077964782715,
-1.53225505352020,32.5707664489746,
12.3380517959595,30.2019996643066,
27.2907924652100,4.58159923553467,
26.3145885467529,-3.42356300354004,
21.7405319213867,15.8953790664673,
26.8273677825928,23.7600269317627,
25.9431762695313,-2.70735836029053,
-1.83879971504211,-29.2602462768555,
-32.8220367431641,-7.10265874862671,
-30.4026947021484,49.2998199462891,
-0.222095608711243,70.5083312988281,
16.8963127136230,27.2541351318359,
9.50231456756592,-27.2476749420166,
-0.381575465202332,-40.5994949340820,
-7.15461587905884,-29.6156768798828,
-29.2450981140137,-31.5947589874268,
-57.8775672912598,-36.1772613525391,
-56.7339859008789,-7.54492092132568,
-13.9001674652100,36.7497825622559,
23.0487995147705,40.5952339172363,
12.7354869842529,-4.19760894775391,
-13.3765077590942,-38.1340789794922,
6.48242378234863,-19.5193939208984,
60.6828994750977,13.3320512771606,
76.9151458740234,7.33680534362793,
31.3886318206787,-19.4207038879395,
-17.1997718811035,-8.69765949249268,
-22.7594928741455,38.6148796081543,
-10.6119155883789,60.0033569335938,
-15.9711685180664,27.5145587921143,
-19.0700092315674,-10.1751985549927,
14.9973201751709,-8.99016094207764,
60.6980857849121,7.68819427490234,
61.2828750610352,-8.04803085327148,
17.9326725006104,-46.2893524169922,
-8.60369586944580,-54.6446723937988,
9.20892047882080,-16.1448993682861,
27.8648471832275,27.4273433685303,
8.03907394409180,37.5840606689453,
-19.6249732971191,31.0502147674561,
-12.1218433380127,32.8710479736328,
12.3028135299683,30.2517604827881,
8.76789188385010,4.66014337539673,
-19.5666065216064,-26.7361011505127,
-32.9350852966309,-26.7371807098389,
-11.3299570083618,5.83350086212158,
16.6038074493408,33.3952636718750,
22.4525852203369,33.3174209594727,
17.7538547515869,17.8684921264648,
21.6922569274902,6.85099029541016,
32.0963401794434,-0.895011067390442,
39.0697860717773,-11.0753393173218,
47.2121315002441,-8.30164909362793,
52.8516273498535,21.0510158538818,
31.6064243316650,50.7153587341309,
-18.2623825073242,42.8602294921875,
-54.8044509887695,-0.567888200283051,
-37.8944664001465,-34.2172164916992,
8.83664703369141,-23.9629039764404,
22.7440681457520,11.2609939575195,
-16.0622348785400,29.0410575866699,
-53.6488265991211,8.37906455993652,
-36.2797470092773,-24.3887367248535,
15.6751003265381,-31.0410594940186,
37.9209632873535,-3.71278476715088,
13.6269693374634,30.7125129699707,
-19.2573852539063,41.2160186767578,
-25.4907531738281,22.6105003356934,
-22.1937618255615,-0.565328836441040,
-35.2438507080078,-4.87642574310303,
-55.4789543151856,0.114431500434875,
-52.7739143371582,-10.3827629089355,
-28.4303722381592,-33.4499130249023,
-8.75618076324463,-37.6392211914063,
-7.44113922119141,-16.5929031372070,
-7.70612335205078,-2.01771473884583,
7.81654167175293,-22.2121772766113,
20.0898532867432,-56.3716163635254,
9.15402126312256,-57.5195236206055,
-11.5052623748779,-21.6995754241943,
-4.48556566238403,6.91832256317139,
38.1766548156738,-1.39601469039917,
79.0842514038086,-19.1768760681152,
79.1981811523438,-9.93603515625000,
38.2698860168457,19.8777961730957,
-5.44310283660889,31.1198291778564,
-18.7696380615234,9.58980560302734,
-0.496249437332153,-12.7705125808716,
26.0391998291016,-8.84232330322266,
33.5805740356445,15.7322139739990,
5.63239097595215,34.9310340881348,
-42.9028472900391,26.5763206481934,
-70.9459686279297,-9.96929359436035,
-47.3392028808594,-52.0806808471680,
10.6560220718384,-68.3643569946289,
50.5964202880859,-41.7003326416016,
35.6671867370606,8.05042648315430,
-14.6088781356812,42.0897674560547,
-50.5832214355469,36.5858459472656,
-48.1726760864258,14.1925306320190,
-21.2599372863770,-4.21713638305664,
6.13624572753906,-25.3592510223389,
24.3465480804443,-59.8629951477051,
29.0193386077881,-79.6055297851563,
20.6977920532227,-46.0289077758789,
11.1508798599243,23.9083080291748,
13.4568433761597,67.5697479248047,
22.0822620391846,50.2966308593750,
14.1468839645386,5.89422988891602,
-11.4841480255127,-11.3460721969605,
-24.0266532897949,-2.95935368537903,
-2.24123144149780,-5.28910303115845,
34.8777542114258,-17.3182067871094,
41.5034217834473,-1.54907178878784,
11.8075008392334,50.1525611877441,
-16.7939224243164,89.6924972534180,
-19.8647956848145,82.1363067626953,
-8.94511032104492,45.1560249328613,
-0.132459282875061,11.3347587585449,
6.70869207382202,-15.5403337478638,
16.9891204833984,-47.0476493835449,
19.8909301757813,-57.6696548461914,
9.13080787658691,-21.0669574737549,
2.70121002197266,36.5826492309570,
13.3003578186035,51.5292243957520,
21.6609630584717,9.94382190704346,
2.30392718315125,-27.2244224548340,
-31.8123722076416,-15.8562717437744,
-34.3444137573242,7.84203863143921,
5.64597558975220,-4.43326187133789,
41.8658027648926,-30.8532657623291,
33.7857551574707,-12.1002092361450,
-0.0114340782165527,49.0706253051758,
-15.7554235458374,75.9282455444336,
-2.60995793342590,26.9676494598389,
15.0010881423950,-46.6592330932617,
12.8046026229858,-67.5086364746094,
-8.88406372070313,-33.7751693725586,
-35.9138412475586,-3.56300973892212,
-53.2057914733887,-8.79115104675293,
-45.0488662719727,-22.3212680816650,
-5.01380634307861,-21.9655666351318,
39.4530143737793,-23.0444355010986,
49.9968566894531,-35.7715721130371,
21.7293968200684,-38.6223297119141,
-5.93527412414551,-8.77355384826660,
-2.65652489662170,33.8528938293457,
14.4841527938843,45.8719253540039,
18.3098125457764,14.5121850967407,
14.7315645217896,-21.0018043518066,
21.5535697937012,-17.8314189910889,
34.5564308166504,18.1608428955078,
24.9320087432861,46.8095054626465,
-12.3560533523560,43.2962112426758,
-37.4645233154297,12.0230283737183,
-17.5902862548828,-19.2746887207031,
23.1351833343506,-23.8058662414551,
43.9414024353027,-3.71172547340393,
35.1315383911133,11.5254459381104,
19.6775836944580,7.90748214721680,
10.3424816131592,5.31962633132935,
-2.03736996650696,27.5541267395020,
-16.7387714385986,64.7732696533203,
-21.3946800231934,77.5297470092773,
-19.2344150543213,53.3025550842285,
-31.5463771820068,27.8753166198730,
-59.0476531982422,34.7859382629395,
-64.1308746337891,47.9434509277344,
-19.1754646301270,23.9657783508301,
34.8670272827148,-18.9384727478027,
33.2041969299316,-26.4456310272217,
-23.4209041595459,3.64802956581116,
-64.1054458618164,14.9857959747314,
-39.8286247253418,-24.2023506164551,
14.0402431488037,-56.5321502685547,
36.1953849792481,-19.8527450561523,
15.6274032592773,55.6111640930176,
-9.75615596771240,88.9944610595703,
-17.7228889465332,59.6695709228516,
-19.4987239837647,28.2312221527100,
-22.8544979095459,28.8217391967773,
-13.6264991760254,22.5464363098145,
6.81240749359131,-24.9492969512939,
8.58961105346680,-63.3736877441406,
-15.7312974929810,-37.0116271972656,
-32.7449913024902,26.8956775665283,
-8.11166572570801,42.7002067565918,
34.0366249084473,-11.3801097869873,
49.0393981933594,-68.6682891845703,
28.9631500244141,-67.5623245239258,
1.06823062896729,-22.6785011291504,
-12.6606788635254,17.0132980346680,
-18.1630268096924,34.5627975463867,
-20.7702789306641,44.0972938537598,
-6.32448387145996,39.0882186889648,
26.3885002136230,11.6526832580566,
45.0329475402832,-8.90652656555176,
25.1113662719727,5.84694766998291,
-18.0173339843750,34.7634315490723,
-49.0927162170410,28.3212223052979,
-50.7366218566895,-19.3721313476563,
-28.3862857818604,-55.6620407104492,
9.52180194854736,-42.8249053955078,
44.0080490112305,-5.70424222946167,
44.8279457092285,9.63240432739258,
4.31892204284668,1.90598368644714,
-42.1291084289551,-0.772432625293732,
-45.9452819824219,0.574609994888306,
-7.51479530334473,-20.8108348846436,
16.2638740539551,-52.7195816040039,
-6.84231090545654,-54.1016540527344,
-40.9405555725098,-18.8633594512939,
-37.8588752746582,3.38160324096680,
0.738304138183594,-20.8137416839600,
33.4375190734863,-58.9770469665527,
43.7257270812988,-55.2529830932617,
44.7017135620117,-9.02207660675049,
39.9007835388184,27.4794273376465,
19.0120964050293,21.0405597686768,
-13.4079446792603,-5.40794134140015,
-19.8479881286621,-13.2806053161621,
14.0758161544800,-0.909968852996826,
46.9367637634277,15.1288576126099,
32.2688369750977,24.5657482147217,
-17.3269367218018,26.1548175811768,
-41.0416831970215,15.7759418487549,
-7.84331226348877,-4.70641756057739,
43.8351974487305,-18.6288757324219,
62.4712295532227,-15.2226486206055,
42.3248291015625,2.96503782272339,
10.9127016067505,16.8587722778320,
-10.4113044738770,12.4787425994873,
-26.4773368835449,-5.91894006729126,
-43.2219276428223,-21.9451007843018,
-50.0345840454102,-26.6066379547119,
-41.2420616149902,-12.1886329650879,
-25.8726348876953,18.1356697082520,
-19.1224536895752,38.2534751892090,
-19.4359111785889,30.1979064941406,
-11.6782236099243,11.0181274414063,
5.49177026748657,8.51230430603027,
20.2237968444824,22.9756393432617,
21.8819141387939,17.8652896881104,
4.72172117233276,-22.6414985656738,
-20.1507530212402,-57.8546066284180,
-33.7347335815430,-37.7607994079590,
-29.2069072723389,16.7507476806641,
-16.2503414154053,33.7763595581055,
-9.93493270874023,-10.7196445465088,
-9.59701538085938,-50.5771408081055,
-1.77070975303650,-21.2463436126709,
10.2547922134399,47.2620506286621,
3.48574066162109,70.3035049438477,
-33.5921821594238,22.8504447937012,
-66.1827850341797,-23.4619636535645,
-53.7559509277344,-5.43796157836914,
-9.08615684509277,47.3830299377441,
11.3509998321533,65.4144973754883,
-15.1196098327637,37.8045883178711,
-46.7791938781738,19.4377384185791,
-41.2140541076660,39.8287086486816,
-12.2617254257202,64.1215820312500,
-4.55718994140625,50.3682022094727,
-22.2332935333252,18.7820320129395,
-30.0865173339844,9.69357109069824,
-13.2678165435791,20.1688709259033,
0.736525654792786,13.1496953964233,
-7.51663637161255,-21.7850818634033,
-14.9310827255249,-48.1329956054688,
2.65426874160767,-40.1295928955078,
31.3433284759522,-22.3675251007080,
38.3801612854004,-35.0301094055176,
21.3177814483643,-66.6705627441406,
5.15638637542725,-73.4458312988281,
-2.34204363822937,-39.2697792053223,
-12.3531808853149,1.45093894004822,
-26.2012538909912,10.9965496063232,
-29.2688865661621,-17.5760955810547,
-12.7116718292236,-53.8914756774902,
6.00533580780029,-68.4480361938477,
9.86880588531494,-50.1784400939941,
6.07281684875488,-11.1773719787598,
11.8124132156372,27.3275604248047,
25.6646595001221,45.3805770874023,
34.6904182434082,38.4304504394531,
36.4356040954590,24.9455928802490,
33.3739242553711,20.1681613922119,
15.2118787765503,20.8450794219971,
-22.7387123107910,19.5527534484863,
-60.4329986572266,12.7014350891113,
-70.8435516357422,2.49523305892944,
-48.9618682861328,-14.5417871475220,
-28.0596694946289,-32.2855987548828,
-34.9034423828125,-39.1632194519043,
-55.6474456787109,-27.2003116607666,
-60.9650421142578,-12.1057357788086,
-44.9128456115723,-20.0486850738525,
-24.0442314147949,-42.7949180603027,
-5.80477046966553,-40.6605911254883,
15.1929111480713,1.12317085266113,
27.3866558074951,49.0261497497559,
8.46081256866455,55.4674301147461,
-33.4358329772949,22.3353385925293,
-50.0030097961426,-11.0614452362061,
-9.13709831237793,-19.7300834655762,
54.8523597717285,-14.7028589248657,
75.9221343994141,-11.2960729598999,
36.0817565917969,-1.53841781616211,
-13.6579551696777,20.7118911743164,
-19.7383365631104,36.6234321594238,
7.73535966873169,18.5395278930664,
23.4615097045898,-24.8696556091309,
5.49299907684326,-55.0224876403809,
-22.8156909942627,-46.3325004577637,
-34.8531303405762,-12.1983375549316,
-27.4126853942871,16.8385028839111,
-17.8110046386719,25.8155593872070,
-18.5161800384522,16.6925601959229,
-28.5791530609131,1.13709223270416,
-37.0968780517578,-11.0255889892578,
-33.8201370239258,-23.0279731750488,
-13.3455162048340,-39.1380081176758,
19.3441371917725,-55.3244705200195,
42.0149955749512,-51.6997070312500,
42.2418098449707,-9.10968589782715,
29.5409336090088,55.1180534362793,
16.2245731353760,91.3579864501953,
6.84375810623169,65.6364440917969,
1.44264638423920,4.98032283782959,
1.09533715248108,-30.5747718811035,
2.47484779357910,-23.9713001251221,
-2.30636405944824,-13.4193725585938,
-18.0403461456299,-26.7326049804688,
-26.2041015625000,-45.0284919738770,
-6.62041378021240,-32.2430076599121,
26.7488098144531,6.44916343688965,
30.0837039947510,31.2318286895752,
-12.1294116973877,24.3606281280518,
-58.3940887451172,6.58026266098023,
-61.7783546447754,-5.01854896545410,
-31.5797290802002,-21.9310607910156,
-9.28285884857178,-41.6573791503906,
-6.66633367538452,-38.1634140014648,
-3.20599555969238,0.877261221408844,
11.5016622543335,40.1446723937988,
12.5194244384766,33.9532928466797,
-13.4757452011108,-0.331747770309448,
-41.6615142822266,-11.7802009582520,
-44.8728446960449,12.5194425582886,
-36.4765739440918,30.0037956237793,
-39.4248161315918,8.06127452850342,
-39.1538810729981,-20.4198188781738,
-8.39534568786621,-11.1431293487549,
35.3069267272949,18.7194843292236,
40.8477859497070,17.6636543273926,
1.32360100746155,-18.0130481719971,
-31.8006076812744,-42.5791511535645,
-18.7840080261230,-22.9149169921875,
20.0637989044189,16.7088394165039,
37.4601211547852,35.2671127319336,
27.2054786682129,28.8577976226807,
14.1165266036987,15.7253789901733,
8.05840396881104,2.54153037071228,
-3.36562061309814,-12.4753217697144,
-21.0195159912109,-14.9906711578369,
-23.2628822326660,9.57715892791748,
-5.19173431396484,37.9940109252930,
7.61518812179565,27.2488536834717,
4.00318002700806,-19.6379547119141,
-3.29103302955627,-44.5319099426270,
3.52828526496887,-8.22153663635254,
17.6892738342285,49.8733139038086,
23.8959960937500,62.4796066284180,
15.8113775253296,23.7403030395508,
-1.46483898162842,-10.7771692276001,
-19.2664108276367,-2.94909715652466,
-27.4483451843262,16.9507217407227,
-13.8126802444458,7.91512870788574,
18.3823432922363,-13.5991210937500,
37.0271949768066,-6.09978437423706,
18.4281349182129,33.0580596923828,
-14.0481595993042,53.4974822998047,
-16.1242923736572,29.5961933135986,
22.8023891448975,-1.60658490657806,
59.0314025878906,2.76758241653442,
51.9475593566895,34.1651840209961,
12.2156152725220,41.2558174133301,
-17.7933101654053,3.84094905853272,
-18.1022624969482,-39.4305763244629,
-7.36180400848389,-44.2618293762207,
-7.03237533569336,-18.4106178283691,
-9.19503593444824,-1.15941321849823,
1.92813992500305,0.193081334233284,
16.1507244110107,14.4372177124023,
7.15172863006592,53.4685935974121,
-27.2496528625488,80.6384887695313,
-53.2559356689453,50.6535148620606,
-37.7866477966309,-21.4024047851563,
7.34074687957764,-60.0201606750488,
40.4216995239258,-19.2471332550049,
35.4604110717773,55.1032409667969,
6.20508241653442,86.7241210937500,
-15.2908535003662,57.5758323669434,
-16.1638851165772,16.9411163330078,
-5.04724836349487,3.82467412948608,
5.63849878311157,-5.97498703002930,
5.76554870605469,-44.0120773315430,
-4.53649187088013,-80.4953689575195,
-13.7870292663574,-59.2569808959961,
-4.52098035812378,7.53527927398682,
20.5252342224121,43.6029357910156,
39.2311935424805,12.3202800750732,
32.2392005920410,-34.5981903076172,
7.35298585891724,-33.0182991027832,
-6.90774297714233,0.953099787235260,
-1.55376744270325,-1.66233348846436,
6.32336425781250,-46.8146018981934,
10.4159431457520,-67.8159942626953,
20.8307571411133,-26.1388854980469,
36.8979377746582,37.1774826049805,
40.3468437194824,57.8919448852539,
23.1588745117188,34.7243309020996,
3.12501788139343,22.4126739501953,
-4.17140007019043,43.8729438781738,
-12.8631620407105,64.4485168457031,
-41.1009826660156,43.9184455871582,
-64.1948623657227,-8.40529251098633,
-37.0229721069336,-57.0321922302246,
32.4564018249512,-67.8352050781250,
76.1631851196289,-32.3728256225586,
51.9687843322754,19.9394855499268,
0.654906749725342,43.9583129882813,
-13.3926143646240,23.8988647460938,
11.6475000381470,-6.44243240356445,
28.5092926025391,0.369956731796265,
16.9669742584229,42.6601600646973,
7.49519062042236,68.0537719726563,
18.3136119842529,42.5939826965332,
21.0884857177734,3.47417426109314,
-8.26653385162354,0.0784718692302704,
-40.1006393432617,14.1667785644531,
-28.3188285827637,-3.54787635803223,
13.7810211181641,-47.2471618652344,
29.7362823486328,-58.2526588439941,
0.837424039840698,-14.5365781784058,
-32.2568244934082,31.0919837951660,
-35.6415100097656,27.3524246215820,
-23.3984947204590,-1.94782876968384,
-23.6346263885498,-5.23109197616577,
-35.1747283935547,18.1404190063477,
-35.1914558410645,19.5803298950195,
-18.1254158020020,-15.2807426452637,
1.42763066291809,-43.7693824768066,
16.8452816009522,-37.3242797851563,
31.7881317138672,-16.1689224243164,
35.4133796691895,-10.4575567245483,
12.6658697128296,-11.6929216384888,
-16.3076133728027,-7.92771863937378,
-12.6206007003784,-10.4501581192017,
25.5059719085693,-23.8887901306152,
51.1838417053223,-24.5122280120850,
30.5150203704834,9.02607345581055,
-14.2369384765625,44.0445213317871,
-40.7997093200684,23.4751567840576,
-36.9767608642578,-46.4571075439453,
-23.9244766235352,-85.0022735595703,
-15.1685733795166,-44.5335884094238,
-3.97763538360596,24.2285614013672,
9.58637714385986,44.5919494628906,
12.4012002944946,10.3142004013062,
8.86141014099121,-24.4533786773682,
19.1204357147217,-29.0508975982666,
43.0311088562012,-21.7602863311768,
55.0306549072266,-16.1225719451904,
38.6259269714356,8.67032718658447,
9.36500740051270,60.9746017456055,
-15.5001077651978,95.0301742553711,
-37.8675918579102,70.8820724487305,
-53.3666572570801,14.2566013336182,
-43.9849128723145,-9.45554828643799,
0.451535224914551,11.2088851928711,
50.0288543701172,23.2810363769531,
59.2222671508789,-6.11327791213989,
27.9018363952637,-40.1396827697754,
-3.40889382362366,-33.6515502929688,
-10.4015989303589,6.17798995971680,
-10.0061931610107,29.8003826141357,
-18.3980751037598,16.0385208129883,
-22.9029407501221,-8.06412124633789,
-11.3104419708252,-18.1151504516602,
0.892352759838104,-25.3435802459717,
-2.27102756500244,-44.0680313110352,
-4.72458934783936,-62.1629905700684,
11.0293588638306,-60.2133827209473,
33.6453247070313,-42.7776947021484,
30.4271774291992,-28.2925453186035,
1.32767486572266,-21.2825202941895,
-16.6908073425293,-18.1639385223389,
-1.92025232315063,-13.1295185089111,
19.0420589447022,-10.2966842651367,
16.5000209808350,-12.3192462921143,
-1.61233234405518,-16.0358657836914,
-12.3286323547363,-19.4350738525391,
-13.6569890975952,-25.6788272857666,
-17.9757270812988,-29.0903644561768,
-18.4201011657715,-21.2278614044189,
-3.10960841178894,-13.4800662994385,
14.7417898178101,-19.0982780456543,
5.68849182128906,-28.1872310638428,
-28.7742938995361,-15.7275800704956,
-47.5491180419922,19.2968883514404,
-22.3723583221436,36.3787651062012,
17.3195915222168,7.09958887100220,
23.3784389495850,-42.1679916381836,
-12.4682979583740,-55.9534797668457,
-52.4332008361816,-24.5790748596191,
-62.7677650451660,3.85975098609924,
-38.8888931274414,-3.40688896179199,
4.85984373092651,-18.9536075592041,
45.8398437500000,-0.444292545318604,
55.4689025878906,39.9526557922363,
21.3465385437012,53.5353050231934,
-35.0716857910156,21.4342765808105,
-66.6197814941406,-12.9752988815308,
-50.0844497680664,-11.9793100357056,
-14.6867218017578,11.4867115020752,
-3.35036587715149,18.7909870147705,
-20.5840911865234,1.90994608402252,
-37.7792968750000,-12.1693792343140,
-35.3092041015625,-4.91214752197266,
-26.1907825469971,6.78179311752319,
-20.7087612152100,3.09155678749084,
-13.6674613952637,-8.55159473419190,
-4.42833280563355,-9.52786827087402,
-4.79157733917236,0.513097524642944,
-27.1379890441895,-1.94040238857269,
-49.4176406860352,-30.5116653442383,
-36.5949592590332,-68.5943222045898,
10.5519447326660,-79.8641433715820,
53.8011703491211,-46.0096740722656,
60.4562492370606,4.21473026275635,
40.9432754516602,26.9565429687500,
27.2838706970215,9.37577342987061,
28.7268848419189,-16.7984199523926,
32.4944534301758,-16.9137935638428,
30.3994331359863,9.65402984619141,
30.2310314178467,33.2522048950195,
31.2978343963623,36.3206291198731,
15.4197521209717,27.3055152893066,
-20.3885135650635,13.7699375152588,
-43.8369178771973,-12.6420469284058,
-25.8812751770020,-40.5705604553223,
12.7874279022217,-36.6955451965332,
24.2010955810547,3.13358402252197,
-1.76474118232727,36.7598266601563,
-21.4004688262939,27.9826889038086,
-4.46535587310791,-2.71746635437012,
22.4656963348389,0.124127864837646,
20.1274242401123,32.0029716491699,
-6.62617206573486,33.4077873229981,
-15.5021276473999,-18.1088695526123,
1.47744798660278,-59.0051727294922,
9.27207565307617,-30.9031162261963,
-14.0131731033325,25.7439708709717,
-37.7203102111816,22.3467235565186,
-30.0371456146240,-46.5199851989746,
-0.310748517513275,-84.3730850219727,
13.6255159378052,-28.4919223785400,
2.89487195014954,58.6630897521973,
-7.43331289291382,73.3578491210938,
-0.457064867019653,7.47663068771362,
15.2223300933838,-50.3802070617676,
22.5092639923096,-43.8674163818359,
17.9921360015869,-10.2928428649902,
8.27569484710693,-13.9411239624023,
-2.40893220901489,-47.2368202209473,
-14.8761901855469,-53.9360847473145,
-22.0371723175049,-17.6626205444336,
-19.0993518829346,15.3020334243774,
-14.9055423736572,7.93531990051270,
-20.5575847625732,-19.5936889648438,
-36.9679603576660,-26.8465766906738,
-49.7952575683594,-11.3129549026489,
-36.7017097473145,2.39819979667664,
8.68070888519287,4.85584831237793,
54.6842308044434,14.6954298019409,
58.0027008056641,42.5026245117188,
12.6071481704712,63.9053421020508,
-28.5592155456543,56.7177047729492,
-12.7911071777344,32.2293548583984,
44.0046463012695,13.8631114959717,
70.6598739624023,10.9763031005859,
33.0559959411621,12.9704198837280,
-24.7065086364746,14.2078828811646,
-36.7936477661133,18.6409492492676,
-4.92289972305298,23.1070499420166,
15.5853738784790,7.73115491867065,
1.44171404838562,-32.8503532409668,
-18.3253936767578,-65.7299957275391,
-14.0245008468628,-61.3322181701660,
3.38153266906738,-23.1761722564697,
11.5390548706055,14.0461168289185,
12.9509840011597,17.4001445770264,
22.3767395019531,-12.0929956436157,
25.7041873931885,-46.4098663330078,
9.53046607971191,-52.7957458496094,
-8.16859340667725,-25.9341144561768,
6.19410419464111,12.4472246170044,
48.3276443481445,25.0036067962647,
67.8805236816406,5.73165035247803,
34.1793403625488,-5.42928457260132,
-12.4562339782715,24.2839946746826,
-15.6666021347046,67.6153945922852,
20.4747467041016,61.2329063415527,
43.4170875549316,-9.86147689819336,
22.1246719360352,-77.1092910766602,
-21.5760154724121,-70.1258392333984,
-39.4671936035156,-6.34015178680420,
-16.3942832946777,39.2991638183594,
23.5797939300537,27.6162796020508,
49.7116127014160,-2.34856009483337,
43.2219047546387,1.59269082546234,
10.0356626510620,32.3409233093262,
-22.7700691223145,39.6606216430664,
-27.9460716247559,4.60496711730957,
-8.06032943725586,-41.7569160461426,
3.24496912956238,-59.2027244567871,
-11.2060718536377,-37.4231796264648,
-19.8591403961182,3.35784125328064,
4.28954744338989,34.6447792053223,
36.2374992370606,41.3793678283691,
23.8847827911377,29.1062049865723,
-39.5816802978516,22.1679229736328,
-89.4575195312500,22.8942489624023,
-66.5798797607422,12.4234495162964,
3.47915935516357,-16.6012248992920,
47.8984680175781,-39.5330123901367,
38.9539337158203,-16.0460700988770,
7.14015483856201,47.5413932800293,
-14.4429426193237,90.8251953125000,
-24.5886287689209,69.5008773803711,
-27.5335941314697,11.3794307708740,
-10.8276882171631,-28.4601688385010,
20.6221771240234,-27.6309661865234,
32.6747932434082,-5.39851665496826,
-0.968341886997223,15.3325462341309,
-46.4964752197266,29.8009395599365,
-49.4337310791016,26.8169479370117,
-9.97804069519043,-4.86238622665405,
18.1569824218750,-44.4703788757324,
6.24553966522217,-52.5479202270508,
-13.2443046569824,-15.2487001419067,
-0.916551947593689,27.8128852844238,
19.0224666595459,35.4321594238281,
7.13313674926758,15.7065582275391,
-28.6641540527344,10.1230764389038,
-42.4814300537109,28.7493228912354,
-21.0575523376465,44.5628776550293,
-9.75876808166504,40.5690116882324,
-37.6777839660645,21.7231025695801,
-69.8244628906250,-0.0473346188664436,
-55.3541450500488,-18.2364139556885,
-3.36896657943726,-23.7968006134033,
24.9732055664063,-6.99308490753174,
4.76658439636231,21.7527160644531,
-23.2825450897217,29.5894947052002,
-16.3477077484131,5.47373771667481,
22.5408458709717,-19.1254844665527,
51.6301689147949,-14.3256397247314,
48.7502212524414,3.03265213966370,
26.5914402008057,-8.92504882812500,
7.70451116561890,-49.1012687683106,
-3.12634992599487,-67.2748870849609,
-10.3910989761353,-40.9600753784180,
-15.3694610595703,-1.82010078430176,
-13.5475387573242,9.50278091430664,
1.22091126441956,-2.25945544242859,
24.7827453613281,0.877136707305908,
41.9511566162109,24.9909515380859,
27.8093395233154,37.3095245361328,
-11.6752099990845,15.2294864654541,
-39.1724815368652,-20.9703407287598,
-21.8693695068359,-37.6604118347168,
29.9295272827148,-27.8020858764648,
69.2234725952148,-12.3463163375855,
63.7854003906250,-6.09248733520508,
32.4527206420898,-11.5419397354126,
14.7439994812012,-26.8586959838867,
20.5133514404297,-47.6652488708496,
32.2355918884277,-58.5535850524902,
31.9117908477783,-45.4757575988770,
18.1292324066162,-14.0669612884521,
-5.94130325317383,13.4900083541870,
-35.4784851074219,21.2480831146240,
-54.8876991271973,16.8726692199707,
-44.9275627136231,16.3932571411133,
-9.52771472930908,22.1311111450195,
18.3949527740479,27.4495449066162,
14.2689332962036,29.1837673187256,
-11.0459508895874,25.8233318328857,
-26.9367942810059,7.65787792205811,
-17.5995216369629,-27.7820358276367,
0.527679085731506,-64.5544586181641,
6.02891063690186,-77.3220825195313,
3.36999106407166,-59.0360221862793,
-0.264884918928146,-31.2886085510254,
-1.09886848926544,-20.5710659027100,
-0.672888994216919,-24.1919498443604,
0.949254512786865,-28.9341335296631,
-0.560918688774109,-24.5069484710693,
-7.54650831222534,-18.1201343536377,
-17.7740707397461,-15.2234582901001,
-15.1439781188965,-17.6762123107910,
1.02359318733215,-29.1162948608398,
8.57430171966553,-45.6653976440430,
-12.1491928100586,-46.7206344604492,
-38.0956459045410,-20.7313652038574,
-22.1000232696533,14.5977010726929,
33.0072822570801,20.8398571014404,
67.3583908081055,-9.81964683532715,
38.4319229125977,-38.6794204711914,
-18.3230419158936,-26.7533645629883,
-34.8453025817871,22.1546497344971,
-3.45687842369080,61.7556533813477,
18.2059364318848,68.8155975341797,
-8.02065563201904,51.7020606994629,
-47.7766685485840,21.2365722656250,
-50.8455505371094,-15.3394088745117,
-21.7217826843262,-39.2752609252930,
-4.07147789001465,-30.1236495971680,
-10.6024770736694,7.11635780334473,
-6.98465633392334,35.7203407287598,
24.2934494018555,29.4457073211670,
56.5713500976563,10.0418128967285,
58.5426750183106,6.39252185821533,
33.3148994445801,11.1628522872925,
7.10017013549805,-0.732109785079956,
-1.79194223880768,-17.7368507385254,
6.87291717529297,-1.10615420341492,
18.0191307067871,42.6075096130371,
24.3633441925049,51.1133270263672,
20.1605415344238,-5.34563541412354,
11.8250560760498,-67.4880523681641,
13.7262973785400,-62.2692756652832,
20.2707729339600,5.73504590988159,
8.32880210876465,51.7248268127441,
-28.6291160583496,28.5629634857178,
-52.6065979003906,-19.6534786224365,
-27.5817432403564,-30.0054378509522,
20.6449699401855,-3.77961206436157,
35.9139633178711,10.2784204483032,
7.79860019683838,1.20231330394745,
-12.7355718612671,-1.62933015823364,
11.8982801437378,18.1535034179688,
45.3973617553711,40.0475502014160,
29.6826477050781,42.2152214050293,
-32.3214454650879,30.4164829254150,
-74.7244796752930,16.1395912170410,
-53.4031791687012,-7.55019569396973,
6.39132690429688,-41.3868789672852,
51.2712249755859,-58.5439491271973,
56.4757766723633,-34.1561279296875,
27.8310279846191,12.4597482681274,
-11.7661266326904,34.2691040039063,
-38.3989143371582,28.0397739410400,
-39.0756912231445,27.4232711791992,
-29.0707817077637,44.6929244995117,
-31.1225357055664,46.5946998596191,
-40.2913589477539,10.3244743347168,
-30.7184028625488,-30.8596305847168,
5.74999380111694,-25.9690647125244,
38.2325172424316,15.2749519348145,
35.0897979736328,34.8323097229004,
15.7001609802246,9.86857223510742,
21.9888954162598,-16.6697635650635,
45.3195571899414,-8.01306724548340,
39.0984992980957,14.5918216705322,
-3.95382642745972,13.2360830307007,
-38.2093544006348,-3.91962099075317,
-31.9990730285645,-2.23137116432190,
-9.35083484649658,21.8155994415283,
-6.35036420822144,34.6032791137695,
-8.22600460052490,21.4780788421631,
13.6913166046143,10.9240865707397,
41.4386520385742,24.2039699554443,
24.0663509368897,42.9980087280273,
-35.5734405517578,32.3051567077637,
-69.5143508911133,-1.61954832077026,
-35.2171707153320,-23.4624042510986,
20.3258094787598,-14.2590608596802,
28.5973472595215,14.4462337493896,
-10.5926532745361,44.4220199584961,
-41.1418457031250,58.4636268615723,
-34.0288314819336,41.4988441467285,
-15.3195190429688,-6.38483142852783,
-12.0941143035889,-59.5775032043457,
-14.8826065063477,-78.8130722045898,
-6.20830726623535,-51.1752929687500,
4.83267879486084,-5.82069396972656,
-1.16130065917969,24.6063003540039,
-11.4895439147949,35.0954513549805,
-2.08642292022705,38.0545425415039,
20.8579082489014,37.1404151916504,
19.4693565368652,28.6744155883789,
-15.8098573684692,22.3856678009033,
-50.1960639953613,25.1949806213379,
-51.8666114807129,23.8131561279297,
-23.0411148071289,5.29708862304688,
9.16360473632813,-17.9333972930908,
26.7596740722656,-19.4150791168213,
32.1400375366211,7.87032794952393,
32.2820053100586,32.9279212951660,
23.0311717987061,28.6763381958008,
12.1477222442627,1.72828149795532,
10.2318201065063,-24.6765842437744,
15.9227390289307,-38.0867843627930,
23.7238254547119,-39.4201812744141,
31.3273735046387,-21.1645717620850,
39.0748138427734,12.3858032226563,
35.6485519409180,30.7319755554199,
12.4935760498047,5.71311855316162,
-13.1381721496582,-39.7103195190430,
-13.6982250213623,-45.3774261474609,
8.13938045501709,7.62613630294800,
15.7594461441040,65.0998001098633,
-13.0126953125000,62.1466064453125,
-39.5262031555176,8.39573764801025,
-14.4931707382202,-28.4674434661865,
45.3090667724609,-10.5135593414307,
71.6028671264648,27.4490890502930,
25.1813869476318,32.7528800964356,
-47.7351760864258,7.63719272613525,
-76.6218032836914,-10.3965673446655,
-50.7934799194336,-3.61025738716126,
-14.7180986404419,7.08384275436401,
-2.59220862388611,-4.06951045989990,
-4.14151144027710,-28.3187561035156,
2.48150539398193,-44.0680236816406,
12.2617607116699,-43.2515220642090,
5.06736946105957,-41.6096343994141,
-14.3020429611206,-51.0902366638184,
-19.3489742279053,-54.0618972778320,
-0.112409710884094,-30.5205345153809,
18.7155303955078,13.6353759765625,
7.63909912109375,49.1238975524902,
-29.3713455200195,42.5251007080078,
-57.1560859680176,-1.12958920001984,
-42.2214469909668,-41.9837684631348,
7.89427280426025,-46.1563835144043,
51.7584037780762,-18.2901134490967,
52.0135116577148,13.6165838241577,
12.7733802795410,32.7563629150391,
-27.9455528259277,42.6758918762207,
-33.3384017944336,48.7131462097168,
-4.67691516876221,39.1914978027344,
25.9749927520752,2.25178670883179,
28.5682296752930,-41.4474983215332,
8.14391422271729,-55.2869796752930,
-6.24791336059570,-21.7938861846924,
-1.80717968940735,31.9289016723633,
2.93277883529663,59.7563514709473,
-13.3698482513428,40.9065933227539,
-41.5003356933594,-3.70902609825134,
-41.5069770812988,-35.4443359375000,
5.40735149383545,-38.0508041381836,
62.1306686401367,-19.3856315612793,
72.9030151367188,2.20252370834351,
25.4380798339844,18.1243019104004,
-30.6917743682861,28.6297264099121,
-38.0525512695313,29.5949573516846,
3.74767684936523,12.3850126266480,
39.8765487670898,-16.9559211730957,
28.2580280303955,-31.0899181365967,
-12.0430049896240,-10.7865810394287,
-28.1712265014648,30.3428230285645,
0.341256767511368,56.4758567810059,
42.4400138854981,43.8805389404297,
53.5325393676758,14.9056434631348,
27.1377182006836,9.15985393524170,
0.245900273323059,30.6106719970703,
-1.47448468208313,48.0219230651856,
6.99275875091553,35.3092994689941,
-4.97516536712647,-0.840509474277496,
-31.5295047760010,-30.3789672851563,
-29.7415657043457,-39.1193161010742,
15.4371194839478,-34.6473846435547,
66.8628921508789,-22.4604167938232,
67.2491912841797,1.29206728935242,
17.4654731750488,27.4880714416504,
-24.2029380798340,27.1598548889160,
-15.2679405212402,-5.99425601959229,
19.6679706573486,-37.2171592712402,
26.0295391082764,-26.9235267639160,
-11.2127447128296,12.7589092254639,
-50.5909309387207,23.4871692657471,
-49.5076713562012,-20.0849475860596,
-10.8515262603760,-69.0814056396484,
33.0846176147461,-65.9193420410156,
52.7703399658203,-22.2132549285889,
40.4890747070313,2.19275617599487,
9.00458145141602,-17.2017688751221,
-22.9192333221436,-35.3320350646973,
-41.4252090454102,-12.5893802642822,
-44.8595199584961,21.7466659545898,
-41.5346527099609,17.9618968963623,
-32.2536201477051,-19.0053558349609,
-17.8864784240723,-34.1336898803711,
-2.86662173271179,-4.02794075012207,
-3.96726799011230,25.6631679534912,
-20.7233867645264,7.15898323059082,
-26.8871974945068,-47.2187728881836,
-10.2097511291504,-76.8079528808594,
7.29812860488892,-52.4613647460938,
-0.134490936994553,-5.07082176208496,
-21.4961357116699,22.2388439178467,
-18.9778366088867,19.3952941894531,
16.5148639678955,2.95926904678345,
42.0024490356445,-2.97299861907959,
21.1200714111328,6.35259914398193,
-29.0118522644043,17.0057868957520,
-60.7481994628906,11.9225549697876,
-59.0810661315918,-6.12904262542725,
-45.2987174987793,-21.3183631896973,
-30.3504104614258,-27.1183242797852,
-5.72690820693970,-29.5608234405518,
26.8177051544189,-42.0122413635254,
40.0159835815430,-51.0712318420410,
22.3428955078125,-31.6839828491211,
4.08639574050903,10.8349189758301,
15.8844795227051,34.4297676086426,
41.5192642211914,19.9871692657471,
38.1632881164551,-8.02639770507813,
2.98505377769470,-13.2439966201782,
-20.0615787506104,3.12590837478638,
-3.49183320999146,14.8276958465576,
18.4389915466309,17.4196376800537,
5.02376127243042,27.2508335113525,
-28.8571796417236,38.2409782409668,
-40.0531044006348,16.5960826873779,
-16.4247398376465,-41.7412452697754,
12.6578178405762,-87.8122024536133,
19.3355579376221,-76.2512435913086,
13.5836544036865,-29.3959045410156,
9.73003387451172,-6.59545183181763,
6.40892791748047,-20.8684844970703,
-2.10963082313538,-33.8436927795410,
-7.46479892730713,-20.7311286926270,
-5.41543865203857,-0.453907936811447,
-13.9308414459229,1.46543192863464,
-41.3392562866211,-10.5600194931030,
-56.8299636840820,-23.2469387054443,
-34.4103507995606,-36.8783149719238,
1.87222015857697,-55.4967231750488,
5.68178510665894,-60.9403800964356,
-27.6793422698975,-35.5578689575195,
-50.6126480102539,-3.61624765396118,
-28.5957965850830,-1.58720159530640,
11.7708740234375,-22.6033916473389,
25.6630992889404,-17.8843784332275,
13.6211919784546,22.8005504608154,
0.845016121864319,51.4972419738770,
-11.5988454818726,35.6313018798828,
-33.9477043151856,-4.10374069213867,
-46.2664566040039,-28.9448490142822,
-22.3047790527344,-35.8614997863770,
18.1009654998779,-45.3609733581543,
25.7784652709961,-54.9575233459473,
-4.85190057754517,-39.5116653442383,
-21.0639114379883,-7.10218524932861,
5.63304901123047,5.43213462829590,
34.4789848327637,-4.15225458145142,
12.2311925888062,-6.03166723251343,
-34.7074165344238,3.53566288948059,
-39.0134239196777,-11.7619524002075,
2.83380866050720,-56.4185676574707,
25.8462982177734,-70.7154159545898,
4.70761394500732,-17.2392368316650,
-14.7853136062622,49.3244590759277,
4.83842086791992,51.9821357727051,
30.2630786895752,2.84841322898865,
15.6033735275269,-9.66385555267334,
-15.1658229827881,44.3483505249023,
-10.6719274520874,84.7118453979492,
20.9922809600830,48.4245605468750,
18.2021293640137,-22.6510486602783,
-36.4696502685547,-41.2718238830566,
-79.3240051269531,-7.26383209228516,
-61.0077819824219,8.91792678833008,
-17.9142875671387,-24.8582477569580,
-9.13640880584717,-64.9667587280273,
-27.4539089202881,-68.8067398071289,
-20.1803474426270,-46.2893218994141,
21.5044689178467,-28.5627021789551,
52.8601570129395,-12.3744010925293,
39.2952079772949,14.4071865081787,
0.980945825576782,37.9472961425781,
-21.9804210662842,24.0137100219727,
-22.4649753570557,-22.7725868225098,
-12.1566486358643,-63.8225326538086,
4.05358934402466,-73.3641128540039,
23.7019729614258,-57.2147521972656,
31.0230731964111,-29.0057334899902,
12.9228267669678,-5.03534936904907,
-9.30178070068359,2.52018141746521,
-4.40096426010132,-7.72553396224976,
22.7695903778076,-16.0298175811768,
41.7698783874512,0.727855324745178,
35.1385192871094,36.9515991210938,
20.8295898437500,58.7772865295410,
21.8043899536133,44.7038116455078,
27.2180290222168,23.0572700500488,
10.2419157028198,24.6228446960449,
-32.6052398681641,40.8641433715820,
-68.4347381591797,34.7016372680664,
-66.4779739379883,1.28595483303070,
-26.3207950592041,-23.9079113006592,
22.2744941711426,-16.1972656250000,
48.6678047180176,13.5137929916382,
39.1934394836426,33.2316398620606,
10.0569286346436,34.8594703674316,
-6.59529733657837,32.0799026489258,
1.76050436496735,31.8214035034180,
18.6929664611816,29.0811271667480,
16.8719425201416,26.0821971893311,
-8.24802780151367,32.7833023071289,
-39.9484672546387,44.8168907165527,
-54.4925727844238,44.1799545288086,
-48.6032600402832,25.4621543884277,
-27.6794242858887,12.7918481826782,
-1.94487428665161,23.1005935668945,
13.9821701049805,38.7085456848145,
3.30628395080566,25.1632061004639,
-31.1761493682861,-11.0035114288330,
-57.1435813903809,-25.0471801757813,
-47.1570892333984,4.45678520202637,
-9.07997512817383,41.1799278259277,
23.7269821166992,37.6297607421875,
36.6325912475586,2.87701630592346,
39.8068733215332,-13.4368162155151,
37.0431671142578,11.5547485351563,
15.4943923950195,39.2158088684082,
-26.8508739471436,34.3270339965820,
-62.2342567443848,11.8641157150269,
-61.2780113220215,7.28267145156860,
-31.5973854064941,19.8934822082520,
-8.71570682525635,16.3077583312988,
-3.72902870178223,-14.9842863082886,
2.97937512397766,-36.1681251525879,
21.1465682983398,-15.1171302795410,
35.4755859375000,29.3309516906738,
26.9843692779541,46.8797264099121,
3.70842719078064,23.0377082824707,
-13.0361480712891,-8.96564674377441,
-17.1845798492432,-7.56778287887573,
-17.1746520996094,29.5147953033447,
-16.6187095642090,54.2143440246582,
-7.50888729095459,28.7878265380859,
0.0585557594895363,-30.4340209960938,
-8.14526557922363,-67.8264923095703,
-29.6455383300781,-50.8498420715332,
-38.1619987487793,-2.62088537216187,
-22.5965194702148,20.6650543212891,
-13.0631484985352,2.50195479393005,
-36.6666908264160,-23.0001277923584,
-75.4894256591797,-23.4062442779541,
-77.7430801391602,-10.9954891204834,
-26.6550064086914,-16.2818717956543,
31.8257923126221,-31.9510974884033,
47.4302444458008,-20.5075759887695,
27.0335712432861,25.4762649536133,
17.2768363952637,60.9775314331055,
39.1111717224121,47.5923194885254,
61.8852424621582,5.22612380981445,
55.8109016418457,-11.1273965835571,
31.6798591613770,17.8504905700684,
17.2846755981445,56.2157821655273,
19.1674594879150,55.9949836730957,
20.1389904022217,14.7341585159302,
12.8264074325562,-23.4789237976074,
8.16817855834961,-24.1755104064941,
13.6282176971436,9.19165802001953,
15.0696086883545,38.6548461914063,
2.61739730834961,28.0901260375977,
-15.9367656707764,-15.7137832641602,
-20.1153488159180,-42.5402183532715,
-4.40727424621582,-19.1586055755615,
26.6749858856201,27.8986797332764,
55.0059585571289,38.8833312988281,
57.0006179809570,-0.121128559112549,
24.8445701599121,-33.8073539733887,
-17.1176986694336,-7.56511878967285,
-34.5262336730957,47.7291374206543,
-14.0391883850098,51.6854591369629,
15.6405744552612,-6.04704761505127,
24.4014377593994,-46.6217269897461,
17.9335842132568,-12.9203643798828,
22.5021800994873,49.6091537475586,
36.5033111572266,58.0662918090820,
36.0384750366211,8.92488670349121,
17.3597202301025,-19.4735050201416,
6.19387578964233,12.7351160049438,
7.37067222595215,51.4719963073731,
-2.37423086166382,37.9202041625977,
-30.0538501739502,-5.08978939056397,
-45.6173019409180,-17.5330295562744,
-18.4953765869141,5.26607847213745,
24.1478271484375,8.87271881103516,
32.1321372985840,-28.8549957275391,
3.33600926399231,-64.9407043457031,
-16.0296993255615,-59.1488800048828,
-2.21361875534058,-29.2865142822266,
13.8521709442139,-8.49404716491699,
3.29071593284607,1.03539311885834,
-15.9364728927612,17.6041011810303,
-16.8048000335693,38.5822296142578,
-12.3858041763306,39.2789306640625,
-31.2376842498779,14.6453456878662,
-54.4315567016602,-4.74070167541504,
-39.0627746582031,-1.00502598285675,
18.5992202758789,8.06438541412354,
62.4651679992676,5.31568527221680,
45.1355628967285,-2.79172945022583,
-10.0380640029907,-5.95977258682251,
-40.0563392639160,-0.677882671356201,
-24.0082626342773,11.4310569763184,
6.62968730926514,25.4014415740967,
17.5805950164795,32.1878814697266,
2.29208898544312,21.0253505706787,
-23.4806766510010,-4.29022216796875,
-31.9781475067139,-13.4721851348877,
-8.76106739044190,8.87135505676270,
31.7127628326416,35.9815788269043,
47.1870918273926,31.1879272460938,
12.2261581420898,6.82022094726563,
-38.0433425903320,8.41809368133545,
-42.9397850036621,39.8882675170898,
7.67133808135986,52.0737953186035,
50.4412536621094,14.9339170455933,
29.1599388122559,-28.5270671844482,
-27.7981586456299,-21.9989814758301,
-45.5333938598633,27.9281940460205,
-12.3127441406250,57.7601547241211,
14.9763669967651,37.4914245605469,
-9.53082847595215,3.26043343544006,
-59.1057586669922,-7.62193918228149,
-77.0966567993164,-6.75602102279663,
-44.4336242675781,-21.8556156158447,
5.21446180343628,-43.6482315063477,
35.5192146301270,-37.8996543884277,
34.4708976745606,-4.20938491821289,
2.85005879402161,21.0281276702881,
-42.1323127746582,18.6059989929199,
-69.5760574340820,-1.52141904830933,
-57.0849952697754,-18.6237564086914,
-22.9409503936768,-32.0650634765625,
-8.66147327423096,-45.6594886779785,
-23.1561298370361,-50.4000663757324,
-30.4051113128662,-34.5219688415527,
-13.2743225097656,-7.69302988052368,
-0.176752254366875,6.84474706649780,
-26.5299797058105,0.754386603832245,
-68.1373367309570,-19.1892757415772,
-63.2117271423340,-38.3541526794434,
3.87836837768555,-43.3750991821289,
70.8211975097656,-24.4356174468994,
80.1800460815430,6.16259956359863,
44.4513092041016,14.9619560241699,
17.0222930908203,-16.2023010253906,
16.7841854095459,-61.5713500976563,
15.9618835449219,-73.7935333251953,
-5.89255619049072,-37.6344909667969,
-25.8214893341064,11.0344371795654,
-24.0646915435791,28.1368255615234,
-10.7833757400513,13.5801773071289,
-13.0630865097046,-4.76206016540527,
-27.4083271026611,-8.91723918914795,
-31.5437049865723,-2.39764237403870,
-16.1534576416016,13.8905153274536,
1.13036417961121,33.6653366088867,
3.88158631324768,44.3733863830566,
1.54700493812561,37.8733177185059,
-2.85631847381592,24.9447917938232,
-12.9567108154297,22.4545974731445,
-25.7944774627686,20.7536582946777,
-29.5456199645996,-6.10637807846069,
-11.1454696655273,-50.3408203125000,
19.9017791748047,-61.8075218200684,
40.0791397094727,-13.3199005126953,
37.1824188232422,48.6571998596191,
24.2291660308838,53.6176452636719,
23.2179260253906,3.94559812545776,
38.9254226684570,-24.5978107452393,
57.4047012329102,9.15850925445557,
50.5231704711914,60.1800231933594,
2.09479904174805,60.1589317321777,
-59.4066848754883,16.2366809844971,
-81.0393600463867,-7.94458913803101,
-44.6998443603516,12.9206485748291,
3.98269653320313,36.8216934204102,
11.8883476257324,24.2042598724365,
-19.6356906890869,-0.901028633117676,
-41.8150749206543,3.61271309852600,
-30.2323303222656,28.5226650238037,
-13.5776033401489,27.8787097930908,
-19.4468727111816,-11.1515293121338,
-21.6559333801270,-49.7789726257324,
10.3486995697021,-56.1157493591309,
50.5245056152344,-41.5031433105469,
44.8897056579590,-32.2518081665039,
-4.28115797042847,-35.0432090759277,
-34.5844078063965,-37.5663375854492,
-14.1680202484131,-32.4649810791016,
11.4239311218262,-26.3745365142822,
-11.4267292022705,-18.9712543487549,
-55.0501174926758,-9.75177574157715,
-54.1743469238281,-7.36449718475342,
2.68566560745239,-17.3859176635742,
45.0015792846680,-25.2261886596680,
20.7790451049805,-14.6275529861450,
-33.2075691223145,3.50857734680176,
-46.6741218566895,7.30721759796143,
-8.79189109802246,-9.01955699920654,
34.2018356323242,-27.1201038360596,
47.2732734680176,-28.8901672363281,
39.7578926086426,-14.8022127151489,
32.8526458740234,3.90572261810303,
28.9422454833984,25.2484416961670,
22.0794563293457,40.5060005187988,
14.1031799316406,35.1590881347656,
3.70591402053833,10.6217451095581,
-17.5448970794678,-4.23583412170410,
-46.1351356506348,4.37267875671387,
-57.2558479309082,7.35565185546875,
-31.4103279113770,-24.1107330322266,
5.59466648101807,-69.4843597412109,
21.2541503906250,-81.0139846801758,
20.4266166687012,-55.0081405639648,
27.4216346740723,-31.4887733459473,
41.1419944763184,-35.2521362304688,
34.4401702880859,-36.9127960205078,
1.56253397464752,-7.26158142089844,
-23.6446590423584,27.2513675689697,
-6.98784685134888,20.6774177551270,
31.2357158660889,-10.5892219543457,
49.4665451049805,-15.8066473007202,
37.4763832092285,14.6371603012085,
15.2438058853149,32.5281066894531,
-10.7435369491577,11.9336118698120,
-39.2901458740234,-13.4222354888916,
-55.1745605468750,-9.51152801513672,
-36.3125038146973,0.469884783029556,
0.0727952718734741,-22.8961238861084,
18.0782566070557,-61.3933906555176,
10.2755298614502,-61.6401176452637,
14.8897027969360,-14.2007808685303,
48.2673187255859,21.6520748138428,
66.6009750366211,14.6616983413696,
31.7327117919922,1.63113296031952,
-24.7182407379150,25.3868999481201,
-32.1348152160645,64.7467498779297,
13.7356729507446,69.7607803344727,
40.2812576293945,45.1277847290039,
4.98237991333008,34.2969131469727,
-48.2752685546875,49.7854995727539,
-57.6593780517578,54.7123756408691,
-25.9183197021484,24.0849628448486,
-10.6359491348267,-9.59031009674072,
-37.5938835144043,-10.0616903305054,
-74.7923126220703,6.86690998077393,
-76.7595214843750,-1.54341816902161,
-40.9597091674805,-34.2897071838379,
4.18109512329102,-46.5035896301270,
32.7845764160156,-17.0351581573486,
33.6963043212891,23.6143817901611,
12.1405057907105,34.0611534118652,
-11.0068225860596,6.16582393646240,
-6.11264801025391,-33.6610260009766,
21.2407493591309,-57.2069511413574,
37.5433311462402,-50.6542892456055,
22.2579936981201,-22.8273239135742,
-3.69104480743408,13.4337320327759,
-9.10742950439453,39.4501647949219,
3.76280856132507,46.5597343444824,
3.11755275726318,42.4705924987793,
-19.1520271301270,36.1260643005371,
-34.7309913635254,28.2694797515869,
-24.6949996948242,23.4506454467773,
-11.9189434051514,30.7948760986328,
-12.3835439682007,41.6033096313477,
-9.28884315490723,34.5599746704102,
21.2843418121338,13.8228578567505,
58.4448471069336,8.16342735290527,
51.1798782348633,34.1487998962402,
-4.01277923583984,59.6677055358887,
-50.4758644104004,35.5413208007813,
-41.8645095825195,-25.6331882476807,
-1.90483343601227,-53.9275283813477,
14.9513864517212,-17.5608940124512,
-0.992176711559296,33.0950660705566,
-9.43707370758057,28.4370574951172,
7.52277803421021,-16.5703182220459,
20.2964820861816,-28.9060802459717,
1.34795558452606,16.0231056213379,
-30.3957118988037,53.0095596313477,
-37.2223739624023,23.8991165161133,
-12.5252332687378,-41.0296783447266,
12.8260421752930,-62.4760513305664,
18.4020252227783,-20.9354324340820,
7.92317581176758,23.5274505615234,
-7.36025667190552,15.3381090164185,
-20.1320972442627,-29.8840866088867,
-28.5733394622803,-54.2211837768555,
-21.2896251678467,-33.7089080810547,
-1.39237022399902,3.56863617897034,
7.50241279602051,28.3015747070313,
-6.08387470245361,36.9124603271484,
-25.6180095672607,41.6867332458496,
-25.6731929779053,47.5050506591797,
-2.97075867652893,45.0671348571777,
19.4546527862549,28.0917968750000,
13.0109577178955,5.44479846954346,
-22.2458381652832,-7.65845537185669,
-52.2521858215332,-13.8914375305176,
-44.7217559814453,-22.2531719207764,
0.985440254211426,-37.8481750488281,
44.8478889465332,-49.1936302185059,
39.6697616577148,-30.9153575897217,
-13.8719072341919,19.7131900787354,
-58.8764114379883,61.2449684143066,
-47.3675117492676,48.0635108947754,
0.814372062683106,-10.9974231719971,
23.2530269622803,-58.6335220336914,
-0.781584501266480,-46.9068679809570,
-22.4968986511230,3.54434967041016,
-2.08946561813355,34.6761627197266,
35.5403327941895,30.1845893859863,
35.8524246215820,24.3677387237549,
-7.06651973724365,45.4247741699219,
-39.6663894653320,64.1984100341797,
-24.0613174438477,45.3911209106445,
8.06074428558350,6.85869359970093,
10.2578973770142,-4.38661766052246,
-14.2168426513672,15.4599037170410,
-25.2060546875000,26.6299686431885,
-1.81837654113770,6.65269422531128,
36.5121955871582,-13.5650196075439,
61.3338508605957,-0.277708530426025,
51.7114562988281,27.2091007232666,
4.84289407730103,31.2571220397949,
-55.7097167968750,11.0458354949951,
-81.7584304809570,-3.80373334884644,
-45.1300201416016,-9.11264991760254,
11.9138088226318,-27.2894115447998,
18.0001144409180,-52.4137191772461,
-33.3287811279297,-46.5123405456543,
-67.2063217163086,-6.53262710571289,
-26.1453208923340,18.8790893554688,
41.2477340698242,-0.0504510402679443,
51.2044258117676,-27.3034553527832,
5.68957996368408,-9.15103244781494,
-15.3063287734985,38.6498489379883,
20.0006237030029,51.8117790222168,
49.5665550231934,12.9385404586792,
12.0580482482910,-23.8742427825928,
-63.0602149963379,-19.0153102874756,
-85.9484558105469,-1.52687156200409,
-29.3965873718262,-11.9845237731934,
46.6123657226563,-34.3954315185547,
70.1707916259766,-32.9161376953125,
29.5614147186279,-13.2851915359497,
-32.6321716308594,-11.2162170410156,
-64.5815887451172,-30.1232738494873,
-44.9874114990234,-31.9302043914795,
4.63156366348267,-0.614615678787231,
24.8396339416504,28.4906826019287,
-9.09918594360352,23.6186370849609,
-47.3839607238770,3.29884815216064,
-26.6588935852051,-1.92108678817749,
46.2525520324707,2.64291357994080,
95.3600616455078,1.62884712219238,
67.0818862915039,9.81633472442627,
0.424278497695923,41.4491271972656,
-30.5311870574951,68.5837707519531,
-15.4431152343750,52.0150032043457,
-8.35664367675781,3.35899424552918,
-29.4742317199707,-16.9402160644531,
-51.9583168029785,11.3978023529053,
-58.4301376342773,33.5830688476563,
-61.7168884277344,-0.364551305770874,
-67.3072357177734,-52.2017440795898,
-46.1654548645020,-50.1777763366699,
7.71780776977539,0.127034664154053,
42.5375938415527,28.6629829406738,
14.2742424011230,4.57423686981201,
-48.1036720275879,-25.4377899169922,
-72.9616622924805,-17.7979564666748,
-44.0363082885742,2.93753671646118,
-19.5627670288086,-7.76694059371948,
-38.4251785278320,-40.3595161437988,
-58.9957847595215,-47.8122215270996,
-35.8077888488770,-22.3733596801758,
11.9221572875977,1.57960641384125,
32.2089424133301,-0.250880241394043,
12.4000787734985,-6.17386627197266,
-14.9166460037231,1.38267111778259,
-25.5199794769287,4.06091499328613,
-24.9739418029785,-15.3304595947266,
-14.4659423828125,-38.9687881469727,
18.0747871398926,-42.9519424438477,
59.1281356811523,-27.3261299133301,
62.6565628051758,-10.5228700637817,
9.90793037414551,-2.16755867004395,
-47.2103309631348,1.77950835227966,
-44.8830604553223,7.81443309783936,
5.81410169601440,15.3769178390503,
35.9684486389160,25.5618133544922,
7.97187089920044,39.2837028503418,
-42.0057563781738,43.3045272827148,
-63.1459884643555,26.8381366729736,
-49.6563835144043,7.10041570663452,
-36.3923301696777,9.25691986083984,
-42.3743019104004,24.5930347442627,
-51.7537269592285,20.5657501220703,
-51.8434829711914,-14.0401134490967,
-50.7690887451172,-45.0165596008301,
-50.3564720153809,-46.5398674011231,
-41.2390670776367,-32.6240348815918,
-16.6931247711182,-31.4803504943848,
10.8452806472778,-39.0661468505859,
28.3957405090332,-24.5066509246826,
34.0422744750977,19.0434360504150,
29.3496303558350,53.8876647949219,
13.6966314315796,51.7849235534668,
-9.92716407775879,26.7971858978272,
-30.3274555206299,4.69479131698608,
-34.9527816772461,-7.29196262359619,
-30.5740108489990,-19.3940620422363,
-33.3679885864258,-31.4920692443848,
-32.3355979919434,-40.7728004455566,
-7.49210166931152,-55.4895324707031,
32.5218162536621,-74.3054962158203,
49.6423683166504,-71.4801635742188,
28.3457641601563,-26.2031497955322,
-5.99806833267212,33.0627098083496,
-19.8429870605469,45.7831764221191,
-11.6937799453735,-5.86113643646240,
-3.87619900703430,-65.2339935302734,
5.05203866958618,-64.5231094360352,
29.2249908447266,-9.58906459808350,
50.5589179992676,36.4524726867676,
33.6287307739258,38.3643302917481,
-14.5213356018066,7.81279468536377,
-34.8758621215820,-19.0171356201172,
3.92762088775635,-21.6037845611572,
49.8767356872559,-1.49676775932312,
38.1825523376465,28.9954223632813,
-16.0966606140137,45.3208999633789,
-37.1525955200195,33.0493087768555,
1.59091401100159,6.97088003158569,
37.1800880432129,4.59916353225708,
12.5246229171753,26.9097385406494,
-47.2599563598633,34.2304420471191,
-69.8825683593750,-0.902631759643555,
-38.3980255126953,-32.5812911987305,
0.648930788040161,-4.54759025573731,
9.56220436096191,60.1879997253418,
-1.73436617851257,86.4555435180664,
-6.45793294906616,37.0401229858398,
-1.66755998134613,-34.3622016906738,
10.8137531280518,-54.1176338195801,
29.2217063903809,-19.5865192413330,
46.0718154907227,17.2341175079346,
41.8642311096191,28.9847297668457,
6.37647485733032,27.6532325744629,
-38.2634506225586,25.3746051788330,
-57.8973770141602,15.0436353683472,
-47.4429168701172,3.10475325584412,
-28.9470977783203,16.1531696319580,
-13.9571723937988,51.9941825866699,
0.915872097015381,63.5121803283691,
9.90536117553711,19.1443004608154,
9.03884792327881,-49.6270828247070,
7.51217460632324,-77.5069885253906,
25.4171657562256,-47.0907859802246,
56.4703369140625,-4.93431472778320,
68.2328033447266,2.96861386299133,
47.8165016174316,-16.5538406372070,
23.5279846191406,-27.2473506927490,
30.6607093811035,-17.5902996063232,
53.6104469299316,2.20358753204346,
51.8794174194336,23.6910934448242,
17.2310104370117,40.1490402221680,
-10.1446084976196,40.3907546997070,
-0.446153044700623,17.8968715667725,
22.7517871856689,-6.14678287506104,
25.9741783142090,-0.0302776694297791,
2.79848003387451,35.9202308654785,
-23.4957351684570,62.1662254333496,
-37.5664634704590,41.5963211059570,
-38.3809509277344,-15.8920869827271,
-21.7248649597168,-63.4952316284180,
13.8399095535278,-74.6627502441406,
54.9244384765625,-52.1227302551270,
74.5519332885742,-14.4764347076416,
59.3895835876465,19.3336238861084,
30.8191566467285,32.8826293945313,
12.7545318603516,26.4842319488525,
9.89733409881592,13.2371168136597,
15.5167417526245,7.95414113998413,
28.2515907287598,11.7458648681641,
42.2829055786133,9.45347499847412,
44.6583480834961,3.94277715682983,
32.0474052429199,14.8785209655762,
14.8621139526367,40.3549804687500,
-1.29740476608276,45.7119102478027,
-21.1716442108154,10.3598213195801,
-50.8304901123047,-28.5891075134277,
-70.1804656982422,-22.4354362487793,
-52.9894714355469,14.9003391265869,
-10.2911024093628,20.8654670715332,
12.0688276290894,-28.8652305603027,
-6.21953821182251,-70.4201278686523,
-30.8549537658691,-42.6669502258301,
-29.7856979370117,25.5160751342773,
-10.7401180267334,48.7464561462402,
1.09752869606018,2.51328325271606,
8.51966667175293,-43.0291213989258,
28.1501522064209,-25.1176471710205,
43.3120117187500,29.3036918640137,
16.5947933197022,52.0934677124023,
-40.1509857177734,26.0508594512939,
-64.8919296264648,-9.47779273986816,
-24.3497581481934,-17.4728832244873,
32.3153800964356,-5.49992227554321,
34.3308105468750,4.46234416961670,
-14.2806634902954,2.58639287948608,
-42.0208702087402,-9.77432441711426,
-19.0390548706055,-31.2771739959717,
14.5204124450684,-48.7853546142578,
10.8027572631836,-41.1685676574707,
-22.1027622222900,-8.33731365203857,
-40.6267166137695,16.1293392181397,
-23.8095092773438,16.5101165771484,
5.77843284606934,16.1829566955566,
19.0513858795166,33.0848464965820,
8.95492935180664,43.2443695068359,
-8.60957241058350,13.8657484054565,
-9.42651081085205,-39.2886924743652,
14.1275215148926,-57.0593605041504,
44.8130035400391,-16.9630279541016,
46.9410095214844,25.4646244049072,
4.31888771057129,17.5335636138916,
-43.7432746887207,-17.9946498870850,
-52.1052131652832,-25.9472675323486,
-22.4436416625977,1.29180324077606,
6.03300714492798,14.0784091949463,
6.91764354705811,-15.3546028137207,
-7.42971992492676,-41.5004730224609,
-8.94575595855713,-21.9817161560059,
8.48079109191895,22.6234054565430,
28.7369480133057,40.0859680175781,
40.6441802978516,21.4519138336182,
35.9857673645020,8.62810230255127,
7.79217433929443,25.3408660888672,
-31.2689838409424,35.9207496643066,
-44.5715446472168,3.96569204330444,
-12.2261543273926,-41.4214897155762,
33.8285560607910,-37.7240562438965,
41.4723930358887,24.1752815246582,
3.73464465141296,80.1425476074219,
-25.2772884368897,62.9749107360840,
-3.94098043441772,-19.9546527862549,
39.9990158081055,-88.5934066772461,
44.5122947692871,-76.1828613281250,
1.21797871589661,-8.19653320312500,
-35.0148811340332,34.2881469726563,
-22.7670612335205,7.22426605224609,
10.0002574920654,-47.4928588867188,
17.0008869171143,-56.4282073974609,
2.00536394119263,-6.61438417434692,
1.84253025054932,42.4796791076660,
23.6683082580566,36.5984191894531,
27.0499134063721,-4.35085391998291,
-6.94693660736084,-26.2121658325195,
-35.2773361206055,-18.1626834869385,
-13.7033882141113,-10.2844791412354,
35.5997734069824,-11.0143728256226,
52.4417648315430,3.16016101837158,
20.6857872009277,42.7607803344727,
-16.9579181671143,74.0645446777344,
-26.6530818939209,65.9335327148438,
-21.6162414550781,36.6513023376465,
-24.8918819427490,16.3663921356201,
-25.0719871520996,1.38516366481781,
-7.39738082885742,-31.3679428100586,
10.8974885940552,-66.1548309326172,
4.30667304992676,-59.2330818176270,
-15.3826818466187,-8.06166648864746,
-13.7807874679565,31.7850914001465,
11.1413335800171,25.3180580139160,
18.9727268218994,1.89222252368927,
-6.69890785217285,4.24002695083618,
-27.3744640350342,19.2991485595703,
-8.27128028869629,6.42411994934082,
27.7249469757080,-26.9573993682861,
30.3228626251221,-31.8021812438965,
-17.5078315734863,6.61608886718750,
-71.6987152099609,34.7028694152832,
-79.1436538696289,7.30472135543823,
-33.3371734619141,-40.3830299377441,
20.5958843231201,-44.0839576721191,
33.6002731323242,-0.116452753543854,
-2.01301765441895,27.6691093444824,
-45.6634292602539,1.15824794769287,
-46.4444541931152,-37.7513847351074,
0.539086818695068,-32.5775184631348,
45.5319862365723,15.8384494781494,
38.4606971740723,51.2458190917969,
-8.54495811462402,35.8430252075195,
-37.9372787475586,-8.71928596496582,
-21.1704978942871,-40.7285537719727,
14.8536520004272,-50.3235054016113,
31.4958419799805,-53.9902458190918,
25.6407184600830,-54.8256378173828,
24.9228935241699,-41.8387756347656,
40.0530319213867,-10.1149187088013,
46.0908164978027,23.3355808258057,
29.9294872283936,32.0166549682617,
2.78028225898743,9.99863910675049,
-13.9747447967529,-15.8046388626099,
-14.1601181030273,-17.1899986267090,
-3.82883310317993,3.04530572891235,
10.4183263778687,18.5046920776367,
24.4825935363770,13.8211927413940,
22.8024215698242,0.811300694942474,
-1.67135882377625,5.70478010177612,
-27.6569633483887,27.0584449768066,
-25.6436405181885,27.7217674255371,
3.33986330032349,-5.88566923141480,
27.8572139739990,-40.3661079406738,
14.5530872344971,-37.3434944152832,
-22.1999778747559,-5.45751190185547,
-45.5954780578613,12.7730684280396,
-38.7937469482422,-0.943095266819000,
-20.2675209045410,-13.7447729110718,
-13.8044471740723,4.97103929519653,
-25.0348758697510,26.7265243530273,
-38.8689422607422,8.30001926422119,
-35.5020446777344,-42.6463546752930,
-7.96148061752319,-71.7551956176758,
31.3779640197754,-54.9695701599121,
55.7330780029297,-31.0827655792236,
49.2880973815918,-42.0857315063477,
29.2088184356689,-66.4098434448242,
31.9642429351807,-52.8314590454102,
63.8003654479981,-1.34493494033813,
89.1152725219727,33.5285224914551,
69.1623153686523,15.8580827713013,
15.5148992538452,-21.8777847290039,
-22.1206378936768,-23.9798469543457,
-22.1746425628662,15.4434719085693,
-4.72972631454468,51.2271308898926,
0.386892884969711,49.8501014709473,
-6.72440528869629,27.1812229156494,
-8.86604404449463,15.5868606567383,
-3.75962901115418,17.7688560485840,
-2.82030701637268,13.1512861251831,
-5.10542726516724,-12.1275758743286,
3.50430440902710,-46.5725860595703,
25.7911491394043,-54.8065872192383,
45.3768234252930,-24.8237762451172,
47.4816436767578,25.4204730987549,
35.6863670349121,54.4015579223633,
16.8227825164795,42.7251167297363,
-5.18884658813477,5.67910671234131,
-27.5725593566895,-20.6856594085693,
-33.2420272827148,-23.2987518310547,
-16.3531284332275,-19.6176376342773,
8.83024978637695,-19.0236968994141,
20.4376697540283,-7.77090597152710,
20.9673900604248,20.6009769439697,
26.4345912933350,41.9060897827148,
35.7484054565430,23.0487937927246,
26.3832855224609,-25.2925243377686,
-7.46172237396240,-49.1652259826660,
-35.2164688110352,-16.3952598571777,
-21.8235263824463,41.7244529724121,
19.6822643280029,67.1146316528320,
39.3091583251953,45.4728088378906,
14.2462863922119,14.9582843780518,
-28.7616691589355,11.9980459213257,
-41.7132301330566,29.0598144531250,
-16.7918643951416,30.5444316864014,
7.45704174041748,6.50444030761719,
-0.277896881103516,-17.8081417083740,
-28.4813365936279,-19.2715053558350,
-37.9751091003418,-4.15793704986572,
-16.3464469909668,2.61948704719543,
9.34628868103027,-13.3053388595581,
4.14025592803955,-34.0361328125000,
-26.4858551025391,-34.8431015014648,
-47.5479278564453,-12.1359519958496,
-35.1859855651856,14.9447364807129,
-13.3338041305542,25.1451072692871,
-17.4307689666748,11.3216991424561,
-44.9926223754883,-12.6346683502197,
-57.0357513427734,-28.0340118408203,
-28.6465778350830,-27.5603542327881,
20.2287387847900,-11.3055000305176,
48.1026535034180,12.7321052551270,
40.8148651123047,34.1594238281250,
24.8997249603272,36.1397781372070,
21.6496868133545,10.8077554702759,
25.9054794311523,-36.0562171936035,
23.1371974945068,-72.5088119506836,
17.0119857788086,-68.6730575561523,
24.9075241088867,-26.7773933410645,
48.1544952392578,14.7552928924561,
62.4356307983398,18.5378208160400,
46.5456199645996,-13.7491569519043,
12.0931491851807,-42.2142829895020,
-15.7817707061768,-37.4943885803223,
-21.1687164306641,-9.84360980987549,
-10.8659162521362,10.9655227661133,
-0.378482401371002,8.64523983001709,
6.17681789398193,-6.87189722061157,
16.2316589355469,-22.0025329589844,
26.8737926483154,-35.8628425598145,
32.4516487121582,-48.7199974060059,
27.6649303436279,-54.9281921386719,
15.7124872207642,-46.4229354858398,
9.25314998626709,-22.2920646667480,
13.1331777572632,4.43368148803711,
15.9734792709351,21.8638038635254,
2.42282915115356,15.1383428573608,
-25.2424736022949,-8.28179168701172,
-36.9958457946777,-22.8654174804688,
-8.32366275787354,-12.3925638198853,
45.1907615661621,13.8618335723877,
73.4424133300781,25.7459278106689,
48.7458038330078,4.70826721191406,
6.37867927551270,-23.2980308532715,
5.62954521179199,-25.8153057098389,
50.8708305358887,-4.29535675048828,
86.4223098754883,15.7599802017212,
65.7485046386719,21.5912094116211,
8.56275653839111,22.6505508422852,
-29.0975589752197,15.6255970001221,
-24.6389961242676,-17.7277317047119,
-2.35231399536133,-64.9542388916016,
6.16663408279419,-74.0734863281250,
-1.36383819580078,-13.5034523010254,
-14.9487085342407,63.3532714843750,
-31.9987220764160,72.3575134277344,
-40.9542655944824,2.92973232269287,
-26.3146114349365,-65.5822601318359,
5.79441165924072,-58.9538192749023,
20.0805530548096,0.278109550476074,
-6.72291183471680,37.0049133300781,
-44.2960472106934,21.5103778839111,
-48.6753692626953,-17.0928783416748,
-15.9066429138184,-43.9273109436035,
13.6439609527588,-49.7992401123047,
21.7842578887939,-39.5296478271484,
28.7857074737549,-14.5345325469971,
52.4029769897461,19.0689163208008,
55.7918052673340,43.3526496887207,
10.9125919342041,49.7928733825684,
-48.0855903625488,40.4519882202148,
-59.4187355041504,17.5147533416748,
-18.9945583343506,-23.9134941101074,
15.4242897033691,-64.7585067749023,
5.51620244979858,-62.2304229736328,
-17.0197849273682,-8.19867610931397,
-12.1989622116089,43.0286178588867,
4.97525119781494,43.4495468139648,
-5.52955055236816,9.65311622619629,
-36.0874748229981,-5.27777814865112,
-41.4335136413574,12.7946186065674,
-15.4165477752686,25.4963665008545,
-8.33368206024170,6.53328561782837,
-42.3357772827148,-18.7013397216797,
-73.6946945190430,-18.3184528350830,
-55.3094367980957,-2.77511477470398,
-9.95658779144287,-2.63223242759705,
10.1763715744019,-16.1909847259522,
-6.21298027038574,-25.7981681823730,
-19.3386859893799,-28.9543151855469,
-3.82560205459595,-37.1974067687988,
12.0388736724854,-38.9195632934570,
1.02586698532105,-15.0146112442017,
-20.3290882110596,20.9834022521973,
-27.1417713165283,41.2898330688477,
-24.7059955596924,41.2060661315918,
-26.1888103485107,39.7597160339356,
-22.4973430633545,42.4778099060059,
-1.44607329368591,24.2844944000244,
21.9341106414795,-21.3304519653320,
30.3701477050781,-52.7983398437500,
33.4203033447266,-36.2097167968750,
55.3851585388184,1.93645298480988,
81.6165542602539,15.8233270645142,
65.9775161743164,10.3284368515015,
4.94718742370606,25.8709945678711,
-39.3222999572754,58.5889968872070,
-21.8662757873535,58.4535903930664,
21.7342777252197,8.59586906433106,
30.0829696655273,-39.9235992431641,
1.67666554450989,-33.0700492858887,
-13.5007572174072,14.6967287063599,
1.75709080696106,47.1134033203125,
12.1865100860596,43.8757095336914,
-3.12602066993713,35.5753898620606,
-11.4995756149292,41.8726196289063,
16.2895259857178,46.2286872863770,
48.5056304931641,30.3537654876709,
34.8304748535156,4.98053073883057,
-12.8479633331299,-14.0890207290649,
-32.4829216003418,-29.3834991455078,
-2.43846106529236,-35.6192245483398,
31.1895999908447,-18.6893196105957,
22.0144138336182,24.6267013549805,
-14.1680793762207,61.7014427185059,
-32.8515472412109,59.9401283264160,
-20.4722137451172,25.7459259033203,
2.05423808097839,-3.93980932235718,
15.0998029708862,-13.2412176132202,
23.4890861511230,-23.3947544097900,
28.8063392639160,-47.2585563659668,
21.2314872741699,-59.5098915100098,
-0.515958428382874,-43.5611953735352,
-15.9126806259155,-12.5462884902954,
-6.46184492111206,2.04626798629761,
16.6147041320801,3.04953169822693,
26.0477390289307,16.5849475860596,
11.5679149627686,48.0376625061035,
-14.1464853286743,67.6875381469727,
-28.0204963684082,50.5676727294922,
-16.8156032562256,10.9231948852539,
9.13891029357910,-16.7515354156494,
30.1546726226807,-21.3306274414063,
38.0199699401856,-14.4570655822754,
40.3995361328125,2.76557970046997,
41.9982757568359,34.7366027832031,
33.1991462707520,69.2572631835938,
6.91881370544434,71.7962112426758,
-20.8938293457031,26.4666862487793,
-22.1061935424805,-32.9813194274902,
6.48806524276733,-58.1331596374512,
28.2473793029785,-35.1287918090820,
16.9681148529053,3.79420995712280,
-7.01839065551758,24.2949390411377,
-9.37905788421631,24.5599117279053,
7.31788301467896,14.4169540405273,
10.5808734893799,-3.03738880157471,
-7.69007205963135,-27.6430225372314,
-12.0444631576538,-41.1954383850098,
17.7879848480225,-26.7410926818848,
46.0906944274902,10.3829851150513,
27.8679656982422,36.7014617919922,
-25.9317207336426,32.7708740234375,
-49.3089256286621,10.6754837036133,
-15.8160562515259,-1.67262828350067,
28.6842861175537,11.6710634231567,
26.4641132354736,32.1206436157227,
-15.9468383789063,35.7393684387207,
-39.3650016784668,15.1743431091309,
-16.4981346130371,-20.5451202392578,
20.8503456115723,-45.0570564270020,
28.1184692382813,-43.8686599731445,
4.41264343261719,-25.7727661132813,
-19.6681060791016,-8.69666194915772,
-24.2379798889160,-4.16980218887329,
-15.7300252914429,-14.5733728408813,
-0.640548467636108,-35.4106712341309,
23.4213047027588,-55.2970924377441,
46.3530273437500,-53.0400238037109,
47.3252067565918,-14.7172393798828,
18.8051013946533,38.3503036499023,
-14.9121532440186,50.7702178955078,
-26.6962795257568,-4.73169660568237,
-10.2128810882568,-79.1713027954102,
19.6491508483887,-94.3231735229492,
45.1812744140625,-38.4034118652344,
57.0199241638184,19.4847354888916,
52.2581214904785,16.6513309478760,
32.7114067077637,-22.6258468627930,
17.7238540649414,-28.4302253723145,
22.4057331085205,15.1699810028076,
33.9523658752441,58.7138977050781,
22.3723030090332,55.5389251708984,
-17.6992454528809,24.0141868591309,
-57.4067230224609,6.85397195816040,
-68.7315521240234,6.76236343383789,
-49.8783760070801,0.980296850204468,
-21.7010498046875,-16.3252162933350,
-2.40843963623047,-22.6560745239258,
5.27091693878174,-8.03445625305176,
-0.242398768663406,2.43151760101318,
-15.8743648529053,-12.3660087585449,
-21.4532051086426,-41.6787796020508,
-2.78867506980896,-63.1754302978516,
25.3145885467529,-61.4437179565430,
36.1977653503418,-38.8050079345703,
24.9981422424316,-4.28689718246460,
19.0595188140869,30.1681270599365,
29.4125251770020,47.0271759033203,
26.6645984649658,32.0580711364746,
-15.7363491058350,-4.27404832839966,
-71.5759048461914,-29.3569316864014,
-82.4472274780273,-26.5924186706543,
-30.4735679626465,-5.51537942886353,
29.7169494628906,15.0207958221436,
36.9043045043945,22.0976657867432,
-6.23893451690674,14.3240928649902,
-45.1334533691406,3.02544140815735,
-42.3028297424316,-5.56798934936523,
-16.1144390106201,-13.9156789779663,
-0.305746495723724,-27.4294281005859,
-4.00530385971069,-40.6812248229981,
-9.58884429931641,-37.2105827331543,
-1.91232252120972,-6.28419780731201,
14.7057256698608,25.3286685943604,
29.3521900177002,19.7654457092285,
35.7804794311523,-22.4011783599854,
33.4336090087891,-51.5953598022461,
28.5248107910156,-25.4406852722168,
25.9488410949707,28.3197078704834,
28.1768684387207,44.1948204040527,
28.1627025604248,-0.764840602874756,
22.9489898681641,-54.0410346984863,
24.5122909545898,-54.4983253479004,
42.7371292114258,-9.39901351928711,
64.5665512084961,26.5753135681152,
61.3470191955566,19.9198417663574,
22.2232131958008,-2.47886419296265,
-22.9728584289551,-3.18648338317871,
-32.4430541992188,14.8355560302734,
0.945099771022797,23.2628345489502,
40.4110794067383,8.87271022796631,
44.9104804992676,-7.37923431396484,
11.4322566986084,-9.26021099090576,
-25.9197692871094,-4.51264572143555,
-31.7095031738281,-10.3405437469482,
-6.90247774124146,-23.1662044525147,
18.9936809539795,-26.0125465393066,
19.3122158050537,-9.15782642364502,
-1.86868369579315,19.0873069763184,
-14.3734540939331,45.1097183227539,
-2.65357732772827,59.8260726928711,
18.1506538391113,55.9279670715332,
23.2112445831299,33.5753402709961,
12.2455759048462,6.81021022796631,
-3.59715747833252,-1.80584180355072,
-12.5409240722656,13.4399662017822,
-16.6636829376221,31.9966602325439,
-17.2415714263916,35.9389457702637,
-9.68691730499268,31.5097007751465,
1.32743930816650,38.3920173645020,
0.420204460620880,49.9998397827148,
-13.5604848861694,36.3584976196289,
-17.3605613708496,-8.47301673889160,
0.946089625358582,-45.2388191223145,
20.9173316955566,-33.7129631042481,
14.4865226745605,14.2082462310791,
-12.2204236984253,45.0548782348633,
-18.5836601257324,23.7052001953125,
14.0959033966064,-24.5727653503418,
52.0829315185547,-47.8775444030762,
56.6486206054688,-21.8587608337402,
31.9746017456055,25.4822483062744,
15.8234815597534,54.1222877502441,
25.2152976989746,46.8267784118652,
36.8851890563965,19.8377647399902,
30.1054725646973,2.09877681732178,
20.7185649871826,4.52025651931763,
34.2648811340332,10.3349704742432,
57.5625038146973,3.61466836929321,
51.5419044494629,-8.18547916412354,
1.08978939056396,-2.55783700942993,
-53.9281234741211,20.6456909179688,
-60.6698913574219,31.8734264373779,
-11.0366592407227,9.66819763183594,
45.2801399230957,-22.7437419891357,
54.3709220886231,-20.1011905670166,
16.1755104064941,18.3036155700684,
-24.3203678131104,44.6039733886719,
-29.6946563720703,23.5204753875732,
-5.77188444137573,-25.1002922058105,
7.64575386047363,-50.6740341186523,
-6.17442512512207,-34.5358276367188,
-24.2236919403076,-9.94816493988037,
-13.8006114959717,-4.29683208465576,
20.7062854766846,-6.68329381942749,
46.2884674072266,5.89439201354981,
40.2458114624023,28.8439865112305,
17.9965515136719,30.9062137603760,
5.65201330184937,5.03351736068726,
8.42527770996094,-17.4236488342285,
3.96582889556885,-4.52874660491943,
-18.3667011260986,28.4738769531250,
-39.1408691406250,37.8278465270996,
-34.5951919555664,10.1636133193970,
-1.86134886741638,-19.3481807708740,
28.3929367065430,-15.7967233657837,
24.9840126037598,10.3222913742065,
-7.93495178222656,19.8308944702148,
-37.5805587768555,-1.00497555732727,
-40.3305549621582,-19.9064331054688,
-22.9802284240723,-7.62842226028442,
-7.92628955841064,25.3033962249756,
-3.82186865806580,47.5364837646484,
-2.65045404434204,47.7749557495117,
2.62304162979126,38.7887687683106,
7.92369937896729,25.2558135986328,
12.2529649734497,5.20457077026367,
22.5556735992432,-12.6068887710571,
35.8821487426758,-7.45408821105957,
34.6388702392578,19.6580009460449,
13.4332447052002,31.1829528808594,
-6.03633117675781,-0.826158285140991,
-0.847218215465546,-48.3414764404297,
19.4914741516113,-55.7673873901367,
29.1211814880371,-12.0887031555176,
22.4849567413330,32.0973052978516,
16.8792591094971,33.8978424072266,
15.4040508270264,8.11091232299805,
3.48615169525147,-6.17258167266846,
-19.0204582214355,-6.00482749938965,
-21.9695453643799,-19.3066177368164,
9.71663570404053,-44.1368103027344,
45.2201004028320,-43.9767303466797,
42.0455360412598,-3.78749537467957,
6.85293769836426,32.0792274475098,
-11.6550540924072,18.9759311676025,
7.04779863357544,-24.4519519805908,
29.0893211364746,-38.8939247131348,
18.1810989379883,-9.40307331085205,
-21.0166091918945,13.9382028579712,
-50.5008697509766,-6.93076848983765,
-43.9954795837402,-40.3616333007813,
-8.64081192016602,-33.4973754882813,
25.3837642669678,14.7942285537720,
36.0268745422363,50.1546707153320,
23.0743198394775,35.4519462585449,
8.05319499969482,-3.58756470680237,
12.6613073348999,-20.6288890838623,
29.6982994079590,-7.87358331680298,
27.6675395965576,9.26701164245606,
-6.40840196609497,10.8135576248169,
-39.7953300476074,1.57055771350861,
-30.1578330993652,-6.46603250503540,
10.4905681610107,-9.19047069549561,
34.6533737182617,-4.93778848648071,
21.9707698822022,1.66383588314056,
-0.00399762392044067,6.20706081390381,
1.97959983348846,3.11612033843994,
17.0416870117188,-7.95686864852905,
13.5171089172363,-14.1226224899292,
-11.2069931030273,-10.3039894104004,
-30.7538833618164,-7.98518848419189,
-30.3738269805908,-7.97451305389404,
-19.3463954925537,1.75430214405060,
-11.3371419906616,18.4287490844727,
-3.57337331771851,25.9437770843506,
1.52838170528412,8.33552837371826,
-7.69703435897827,-19.4975528717041,
-30.0352191925049,-32.4090728759766,
-40.9441184997559,-30.5942592620850,
-25.9296684265137,-34.9887466430664,
3.99017906188965,-40.3060455322266,
28.3294143676758,-14.1940135955811,
38.8321914672852,46.3227119445801,
41.1950836181641,82.3966827392578,
37.4483833312988,42.8654441833496,
24.2133865356445,-36.3477401733398,
11.8944530487061,-64.2620620727539,
11.9485015869141,-7.69814920425415,
12.8653383255005,64.5076217651367,
-7.34587764739990,67.0767364501953,
-34.3165321350098,2.97005939483643,
-32.5606956481934,-55.3597869873047,
2.46685004234314,-60.7164726257324,
24.0488491058350,-31.0984973907471,
-5.06119537353516,-9.79027175903320,
-53.4001426696777,-7.79043245315552,
-57.5231742858887,-11.3474903106689,
-14.3592033386230,-15.5483388900757,
16.8163852691650,-22.8347587585449,
-6.80218601226807,-24.5136051177979,
-48.6490364074707,-9.95371723175049,
-52.1438865661621,10.9552183151245,
-18.4047718048096,20.0087833404541,
-3.52179598808289,2.24098658561707,
-29.8604316711426,-26.9053726196289,
-57.2460632324219,-33.7054939270020,
-42.0722274780273,-11.2168121337891,
2.84178018569946,12.8417081832886,
28.5945758819580,7.75300025939941,
13.9671707153320,-23.0972194671631,
-9.60963821411133,-42.8723526000977,
-7.08265304565430,-21.9369945526123,
18.4765110015869,12.8175926208496,
38.9168548583984,10.8854713439941,
35.4695358276367,-32.2597999572754,
18.2417182922363,-58.0682868957520,
5.08135318756104,-20.7899780273438,
9.72550964355469,48.5290298461914,
25.0438194274902,75.5151672363281,
25.2235984802246,37.5568199157715,
1.94305324554443,-15.9528694152832,
-25.0113182067871,-35.0865135192871,
-20.3384151458740,-28.5894203186035,
19.6185588836670,-37.8456344604492,
51.4318885803223,-57.8076858520508,
30.8989772796631,-50.6417884826660,
-22.2984066009522,-10.2772197723389,
-47.0650482177734,22.1990242004395,
-17.7194213867188,13.9296970367432,
29.2771644592285,-14.9512901306152,
45.5662231445313,-18.0491905212402,
32.0278739929199,9.80573081970215,
18.2470741271973,36.2683105468750,
11.7376537322998,42.2412796020508,
-8.85355186462402,37.2731971740723,
-43.3077926635742,27.9574546813965,
-57.1497993469238,2.95196175575256,
-27.9298191070557,-47.4714355468750,
18.9861907958984,-89.3817825317383,
33.1010322570801,-78.7953948974609,
4.91411304473877,-21.1402778625488,
-25.5983963012695,32.0512275695801,
-18.6943893432617,40.5783576965332,
15.3711185455322,19.8613376617432,
35.5083961486816,11.3681812286377,
17.5015697479248,26.8357162475586,
-21.6165027618408,40.3730659484863,
-39.0803794860840,28.6844501495361,
-23.8952713012695,5.72039747238159,
-4.99889230728149,-1.14629185199738,
-8.63365840911865,13.5616569519043,
-25.8484935760498,36.2346305847168,
-21.8540916442871,49.7035217285156,
9.61566543579102,43.1214485168457,
43.0416259765625,16.1101551055908,
49.6915817260742,-12.8069648742676,
39.5159263610840,-15.7909965515137,
34.4015693664551,13.6392078399658,
27.8517761230469,50.9178886413574,
-0.0620892047882080,52.7906494140625,
-37.9212989807129,10.5927181243896,
-44.0534553527832,-38.2595329284668,
-3.65484499931335,-62.2205047607422,
43.0654907226563,-58.9003829956055,
49.5091400146484,-37.7369766235352,
19.2583560943604,-3.29149866104126,
-9.08443355560303,29.1399059295654,
-20.0756721496582,33.8403091430664,
-31.0245094299316,6.67652130126953,
-48.9155464172363,-14.4741048812866,
-55.7021903991699,6.43966007232666,
-38.8217315673828,42.0582046508789,
-16.6189823150635,32.2841072082520,
-8.40036392211914,-19.7403964996338,
-1.99246549606323,-43.7847709655762,
12.6872138977051,-2.66051244735718,
16.8182220458984,45.7954940795898,
-9.71371078491211,30.9148941040039,
-43.6170997619629,-22.4130115509033,
-40.0049781799316,-35.5971183776856,
0.299743533134460,6.45140171051025,
27.7182178497314,40.6038475036621,
11.1774168014526,19.1935348510742,
-24.2748336791992,-13.8446664810181,
-34.4699363708496,-6.30262088775635,
-21.4113864898682,19.8266868591309,
-16.0985488891602,9.30375671386719,
-22.4156684875488,-39.5570983886719,
-16.5057621002197,-67.3436737060547,
3.39573359489441,-46.4272956848145,
11.9834957122803,-12.0807113647461,
-4.85016584396362,-2.22535657882690,
-26.1828098297119,-5.84819602966309,
-24.8664207458496,-3.17474508285522,
-2.47141981124878,0.956092000007629,
20.3889904022217,-10.2443342208862,
30.6195640563965,-22.9439582824707,
28.0140552520752,-5.17165184020996,
13.2862062454224,39.7139396667481,
-10.4008522033691,65.7949600219727,
-24.4956588745117,40.8346481323242,
-14.9682321548462,-12.4742717742920,
5.55390787124634,-47.8578224182129,
7.36991167068481,-49.7965850830078,
-14.0024023056030,-36.3819618225098,
-29.3351325988770,-29.5184116363525,
-16.4594421386719,-36.5128746032715,
10.6531801223755,-46.9003601074219,
20.3179950714111,-55.4971199035645,
5.31729936599731,-61.0608139038086,
-6.19166612625122,-58.5428657531738,
9.84255599975586,-39.7693939208984,
40.2299118041992,-5.15947055816650,
55.4375991821289,27.3004302978516,
48.3530044555664,34.4528083801270,
38.2405853271484,15.5389633178711,
42.6433029174805,-5.65032434463501,
52.4268302917481,-4.36383676528931,
46.4358291625977,22.4519214630127,
19.9184303283691,41.3544998168945,
-12.7655029296875,31.2238769531250,
-29.6348457336426,4.91024398803711,
-24.5928859710693,-13.8459653854370,
-5.41992092132568,-14.4553594589233,
14.9633522033691,-8.32905864715576,
21.8616390228272,-0.495346188545227,
13.2660179138184,11.2421483993530,
1.46871232986450,19.7591495513916,
-1.11557185649872,8.25064182281494,
0.605951428413391,-21.9950733184814,
-2.03318309783936,-35.5185737609863,
-7.12099170684814,-6.89186191558838,
-7.90272474288940,30.1746330261230,
-0.783177316188812,16.9259662628174,
4.17024612426758,-44.7954902648926,
8.24242305755615,-85.7779083251953,
24.1723384857178,-53.9925765991211,
48.0394325256348,15.5541934967041,
47.4324150085449,48.3578987121582,
6.86644268035889,34.1347656250000,
-42.0785408020020,24.5127010345459,
-52.7074012756348,46.8358879089356,
-26.3229656219482,63.5198287963867,
-12.6747903823853,44.3606758117676,
-34.1466560363770,20.8803749084473,
-54.9166450500488,30.7746906280518,
-34.4506950378418,47.8709144592285,
17.4151115417480,19.5620689392090,
55.5229301452637,-43.4264869689941,
58.1516838073731,-63.8735275268555,
47.4574012756348,-8.11620807647705,
49.9539794921875,55.7313728332520,
58.4311904907227,51.5049324035645,
52.3425140380859,-5.94213390350342,
20.5117206573486,-41.5879783630371,
-21.7412586212158,-22.9682369232178,
-45.3120536804199,0.905463755130768,
-30.6479549407959,-8.79009532928467,
11.6414337158203,-25.8035488128662,
38.1816177368164,-11.1810312271118,
15.7097244262695,16.2464656829834,
-30.3784923553467,10.6993665695190,
-44.8182334899902,-30.9704723358154,
-8.14590454101563,-51.2975463867188,
35.6990852355957,-15.4364452362061,
27.1714763641357,45.5337409973145,
-30.8330421447754,67.8475723266602,
-76.7926864624023,32.7620468139648,
-64.7959365844727,-15.0654067993164,
-6.62250518798828,-33.1127433776856,
46.1109733581543,-18.5620822906494,
59.7832489013672,5.62939071655273,
36.1033935546875,22.4843730926514,
3.51320314407349,32.4827156066895,
-10.1313638687134,39.4529113769531,
5.16559982299805,39.5992507934570,
38.7673912048340,30.8758926391602,
61.3411407470703,25.8411216735840,
51.5026550292969,39.1636734008789,
14.7916049957275,61.3864822387695,
-20.9241962432861,61.5222702026367,
-34.4810295104981,25.3326568603516,
-28.8909912109375,-25.3572711944580,
-15.7297286987305,-52.5231513977051,
7.93473672866821,-38.3217353820801,
46.8656349182129,-7.70451164245606,
80.7703552246094,15.4441070556641,
81.8316574096680,27.2515392303467,
44.2318878173828,32.0343399047852,
6.80881214141846,21.5435886383057,
6.02200078964233,-8.89590549468994,
25.3234767913818,-38.1773338317871,
22.1371192932129,-32.7959175109863,
-7.70924568176270,-0.432767152786255,
-24.5468864440918,14.5886306762695,
-2.10996198654175,-9.12687206268311,
29.8682994842529,-36.1380233764648,
30.6120967864990,-15.7977228164673,
6.25347995758057,41.1393508911133,
-8.99817085266113,80.2547683715820,
-4.79939699172974,69.3874435424805,
-10.0517053604126,35.2663345336914,
-36.8835716247559,21.1229763031006,
-56.4377288818359,25.4717636108398,
-45.4793891906738,18.8326206207275,
-17.3042945861816,-7.41422176361084,
0.776290059089661,-37.1754837036133,
10.1538600921631,-49.8249855041504,
24.8825225830078,-43.4203262329102,
36.6315460205078,-25.1760711669922,
23.6897640228272,-0.0653518140316010,
-7.89927101135254,20.6776371002197,
-31.0557308197022,31.0084762573242,
-32.4305839538574,32.2633361816406,
-32.7875022888184,27.2709846496582,
-41.4549293518066,15.7897558212280,
-34.9586372375488,-5.38731098175049,
1.30617833137512,-24.4674625396729,
34.9471702575684,-14.9338693618774,
26.5868167877197,25.0933227539063,
-11.0120449066162,62.8126716613770,
-24.0928783416748,62.9052200317383,
9.36939907073975,29.3512973785400,
52.0402870178223,-4.08054161071777,
56.3398742675781,-8.98652267456055,
26.6696872711182,16.9444370269775,
-2.53722524642944,48.3242950439453,
-21.0790805816650,59.1374931335449,
-41.4954566955566,35.6696205139160,
-65.9220657348633,-9.29100418090820,
-68.9597778320313,-38.6968803405762,
-40.5177650451660,-28.5826721191406,
-10.8208847045898,-1.55215322971344,
-7.62525177001953,0.585967659950256,
-17.0347080230713,-25.8182258605957,
-7.35243034362793,-41.1970520019531,
23.9174118041992,-17.9352626800537,
42.3920364379883,14.2634477615356,
21.0216655731201,9.21595668792725,
-17.0115184783936,-22.0283126831055,
-28.4440422058105,-26.6097049713135,
-7.10016298294067,18.7352848052979,
8.54934692382813,63.9542007446289,
-10.9787511825562,48.2055625915527,
-49.2944717407227,-17.7453193664551,
-57.7907829284668,-63.6876754760742,
-11.4904518127441,-47.7100639343262,
55.8580551147461,-2.44693946838379,
83.3938217163086,12.8375053405762,
50.3809280395508,-13.6123113632202,
-4.07670879364014,-39.9272766113281,
-24.2448596954346,-30.4283485412598,
-1.62093472480774,0.497344732284546,
25.9316387176514,23.3718624114990,
27.4770030975342,24.8218212127686,
12.1194829940796,15.5305671691895,
8.10777282714844,0.733289837837219,
16.6685428619385,-21.2105636596680,
22.0352249145508,-39.3535842895508,
19.4200477600098,-33.1833076477051,
21.1214065551758,-1.87304449081421,
30.2139091491699,24.7454814910889,
28.7567367553711,30.5964355468750,
1.26091051101685,27.4979152679443,
-41.8827552795410,34.5196418762207,
-67.9607696533203,39.2888793945313,
-61.8025970458984,11.7116260528564,
-29.4323062896729,-41.9475135803223,
2.70855069160461,-76.8884506225586,
14.5493288040161,-66.0921783447266,
13.1451244354248,-32.7777481079102,
18.1450443267822,-13.3575668334961,
34.5356941223145,-12.2054252624512,
44.4663581848145,-4.93138217926025,
25.6495780944824,14.1461887359619,
-10.2270164489746,19.5893707275391,
-30.0143356323242,-3.06044912338257,
-20.2258472442627,-34.0426254272461,
-4.59231710433960,-47.5278053283691,
-5.52898883819580,-43.5335006713867,
-7.45684623718262,-33.5654678344727,
16.5592193603516,-24.5909099578857,
50.6538276672363,-14.1704730987549,
54.3168525695801,-5.11207008361816,
15.5418338775635,6.47902488708496e-05,
-27.7315483093262,12.8812103271484,
-35.1113052368164,34.1007537841797,
-8.13722229003906,43.7075576782227,
22.8885383605957,14.3368864059448,
37.7392311096191,-33.5019645690918,
38.3571548461914,-46.1703147888184,
25.4197368621826,-2.90318632125855,
2.85003590583801,48.6879730224609,
-12.8964900970459,49.6878013610840,
-0.0546975135803223,9.69138431549072,
29.7950344085693,-5.66012954711914,
38.3896598815918,32.9466361999512,
6.57025909423828,83.0859222412109,
-38.8194198608398,85.2618026733398,
-56.4267349243164,36.1752166748047,
-41.9771995544434,-13.3108501434326,
-28.5908470153809,-25.1770744323730,
-30.0551643371582,-15.4071693420410,
-24.4829692840576,-20.6471424102783,
3.59559464454651,-40.2246322631836,
28.2928428649902,-39.8447380065918,
22.0230846405029,-5.35818958282471,
0.521850526332855,31.9660987854004,
7.33986377716064,28.7459907531738,
45.7150459289551,-13.3918838500977,
63.3061904907227,-35.4364166259766,
25.7835617065430,-0.548223257064819,
-24.3811912536621,46.7528305053711,
-24.8754673004150,36.0916099548340,
12.5967388153076,-30.4432353973389,
22.1137657165527,-77.2203903198242,
-18.3958892822266,-53.9087142944336,
-46.9866142272949,-3.91175961494446,
-12.5877637863159,-2.32591700553894,
41.4773864746094,-43.7448768615723,
38.4606933593750,-58.1223182678223,
-21.0357532501221,-14.1737051010132,
-62.6809043884277,28.6460208892822,
-49.9143104553223,15.9159259796143,
-24.1004734039307,-29.4218959808350,
-30.9125633239746,-45.4663581848145,
-46.1322517395020,-24.9020195007324,
-24.8627910614014,-13.2838287353516,
21.3082542419434,-30.9620456695557,
32.8466339111328,-44.4579429626465,
-2.95120859146118,-21.9011363983154,
-37.3424797058106,17.5575866699219,
-32.9188041687012,39.4983520507813,
-8.82696342468262,40.1706047058106,
-6.15037727355957,32.5971908569336,
-28.8997535705566,11.0392332077026,
-39.7440032958984,-35.6711044311523,
-14.7892093658447,-83.5966949462891,
23.7788677215576,-85.5087356567383,
38.5522918701172,-42.4926795959473,
24.7690773010254,-7.72154664993286,
8.72040843963623,-20.1635704040527,
16.2362461090088,-44.2461738586426,
40.0956153869629,-24.6110801696777,
46.3518180847168,33.8152542114258,
18.8242568969727,69.1086730957031,
-11.3352766036987,49.6969451904297,
-10.3642730712891,15.2706699371338,
14.8591346740723,15.7887411117554,
24.7690925598145,35.2201614379883,
1.46779942512512,20.3749008178711,
-26.8819217681885,-33.5020904541016,
-28.3171157836914,-73.4509429931641,
-11.2110185623169,-58.9278907775879,
-10.7557659149170,-20.9663486480713,
-30.7423305511475,-17.6452941894531,
-31.7986164093018,-57.2812957763672,
7.58994054794312,-87.7679290771484,
56.2590522766113,-60.5656700134277,
63.0992698669434,3.44932150840759,
16.7007846832275,42.9404525756836,
-44.2645530700684,34.2935867309570,
-73.2756881713867,5.26831245422363,
-56.8813285827637,-1.74212586879730,
-9.17706775665283,18.9352054595947,
40.4536247253418,30.1298084259033,
63.2707405090332,12.6056442260742,
39.4373245239258,-10.2965850830078,
-17.8550643920898,-9.89179897308350,
-61.0592994689941,4.34131240844727,
-51.3319511413574,1.05552268028259,
-4.40129137039185,-18.7718982696533,
24.9097919464111,-18.5172863006592,
9.89433479309082,18.5459136962891,
-20.4514350891113,51.8323974609375,
-27.3264179229736,23.9521636962891,
-14.9551000595093,-47.1196174621582,
-7.41837072372437,-83.9991226196289,
-5.49753332138062,-46.4413833618164,
14.4030704498291,18.8189468383789,
52.6736106872559,36.9813461303711,
67.5620956420898,1.97530770301819,
40.1416816711426,-30.6351432800293,
5.91571521759033,-22.3378887176514,
3.22104501724243,5.09595394134522,
21.6900043487549,20.8202724456787,
21.7825222015381,20.1494197845459,
-3.99008464813232,11.7560367584229,
-23.4221267700195,-9.96176242828369,
-15.4333152770996,-48.6523704528809,
5.70460987091064,-79.0010528564453,
20.7408847808838,-67.3125152587891,
25.3385944366455,-16.8970966339111,
16.6407566070557,28.1761512756348,
-15.6439428329468,36.5858535766602,
-49.7523994445801,20.9449367523193,
-40.4959335327148,6.16609430313110,
20.0490303039551,13.5986309051514,
70.6376724243164,38.4677505493164,
45.4343338012695,58.0793991088867,
-27.3749618530273,49.3023185729981,
-61.4466285705566,7.70616149902344,
-21.9045124053955,-40.4184379577637,
27.0073909759522,-53.0929450988770,
15.3996734619141,-25.0587940216064,
-41.4787826538086,4.45714139938355,
-67.6414260864258,0.308876037597656,
-38.6662368774414,-19.3575229644775,
-4.54384231567383,-15.5871295928955,
-14.8552742004395,7.06388235092163,
-49.7227821350098,3.36891841888428,
-57.5423965454102,-41.7647552490234,
-21.2492389678955,-83.9174804687500,
25.3199729919434,-71.0571823120117,
44.2883377075195,-17.1659164428711,
32.1644134521484,16.5681076049805,
14.3285942077637,0.435446977615356,
15.3631887435913,-28.9179077148438,
26.7834815979004,-31.8974246978760,
25.1722793579102,-6.17798709869385,
3.65926694869995,20.7088871002197,
-26.8419589996338,36.9283828735352,
-43.3514328002930,48.4440917968750,
-43.8702049255371,44.2095451354981,
-44.9747390747070,11.2103147506714,
-57.2699089050293,-35.9372749328613,
-61.2586860656738,-54.7864913940430,
-42.1187171936035,-28.0027656555176,
-10.6055393218994,9.75407981872559,
12.1195306777954,17.2199802398682,
21.5594902038574,-0.523165166378021,
30.8521308898926,3.07683539390564,
38.0105667114258,37.0715179443359,
23.9924030303955,64.9830780029297,
-11.1476049423218,54.4237060546875,
-34.6796302795410,16.4878845214844,
-17.4789905548096,-14.2643890380859,
25.2531871795654,-16.1435966491699,
54.6797599792481,1.10750973224640,
53.8584671020508,21.1061687469482,
45.1536750793457,34.3185119628906,
43.9313735961914,30.9692344665527,
40.7695236206055,11.8702192306519,
28.5944938659668,-7.38544893264771,
15.1019954681396,-13.7097692489624,
9.57674598693848,-21.4606952667236,
1.03292965888977,-43.3384513854981,
-16.9139022827148,-55.2891044616699,
-32.1930961608887,-30.6763896942139,
-27.8260021209717,12.3252687454224,
-14.4964456558228,18.1176605224609,
-9.02564334869385,-25.4151954650879,
-4.46912193298340,-64.8182525634766,
20.4034328460693,-44.5216941833496,
55.2513656616211,6.66935253143311,
53.2499465942383,23.0555706024170,
0.933177709579468,3.09102773666382,
-48.6707916259766,2.01366662979126,
-48.4513893127441,30.5611972808838,
-9.20263004302979,31.8508777618408,
17.0479507446289,-21.7636547088623,
11.7825136184692,-68.4990463256836,
2.60949254035950,-43.6884498596191,
14.0224313735962,25.4562053680420,
27.4483718872070,55.7425689697266,
27.4508094787598,31.8227424621582,
22.2062644958496,12.7130556106567,
18.0803470611572,34.9598999023438,
-2.91409683227539,56.9385108947754,
-35.1444587707520,33.1757469177246,
-35.3653564453125,-12.4133749008179,
14.8928928375244,-30.6816043853760,
61.4472389221191,-23.6433048248291,
34.0361557006836,-21.7176265716553,
-42.0196037292481,-22.7779903411865,
-68.2119903564453,-5.35153770446777,
-6.84698581695557,20.3508892059326,
55.1584472656250,19.3074760437012,
24.3737907409668,-12.0499849319458,
-64.7375717163086,-39.2031517028809,
-99.2214889526367,-37.5881423950195,
-49.9880828857422,-23.1414680480957,
-2.49409580230713,-19.9120235443115,
-18.6014499664307,-17.5949325561523,
-52.5740013122559,0.822746157646179,
-30.2565574645996,21.0459823608398,
31.6190013885498,23.7756919860840,
56.8585624694824,20.0197219848633,
25.2719135284424,24.5324230194092,
-3.99298644065857,32.8605651855469,
12.0860013961792,32.8419342041016,
38.6692581176758,31.6741428375244,
23.8214263916016,38.3965034484863,
-18.8617362976074,37.8294754028320,
-39.5101852416992,10.7721252441406,
-26.9206962585449,-26.1166801452637,
-6.06387138366699,-31.7841873168945,
4.77434110641480,-4.90045213699341,
9.08675384521484,3.56821012496948,
13.8615741729736,-34.7973251342773,
15.6605710983276,-74.4461593627930,
16.1710262298584,-57.5886230468750,
23.1736106872559,-0.221464157104492,
30.1589679718018,37.5694808959961,
17.0359687805176,37.3210296630859,
-12.1440258026123,33.7718048095703,
-23.5289249420166,51.5919494628906,
-7.67679834365845,64.8680648803711,
2.71127915382385,45.4413871765137,
-14.9502143859863,13.9006404876709,
-29.3961868286133,7.21920394897461,
-5.06966400146484,21.6754531860352,
40.3261833190918,25.2997188568115,
46.2438507080078,8.89118957519531,
-4.07697677612305,-2.87692666053772,
-53.2047576904297,-0.265596032142639,
-49.2609901428223,-6.77278995513916,
-6.88391256332398,-30.3171234130859,
19.0544548034668,-42.3409080505371,
14.0216112136841,-18.0528068542480,
2.26866626739502,22.1350116729736,
-1.07503688335419,32.6416969299316,
-7.59117317199707,-4.04818487167358,
-17.2584686279297,-54.1751365661621,
-4.61182498931885,-72.3203811645508,
38.6554565429688,-44.7744750976563,
76.7068405151367,1.99316060543060,
68.6805038452148,36.1592864990234,
17.3251686096191,36.2219848632813,
-26.9572162628174,9.80494976043701,
-27.0183200836182,-12.7475967407227,
6.89535093307495,-8.66635799407959,
41.0034408569336,15.1117181777954,
56.5711593627930,33.5514755249023,
55.5609474182129,37.6386070251465,
42.9751091003418,38.3982009887695,
24.7234725952148,39.8369369506836,
2.27762222290039,25.8738498687744,
-18.8784904479980,-9.27378940582275,
-24.2081794738770,-38.6536674499512,
-4.09473705291748,-27.6439990997314,
35.4260520935059,17.4618721008301,
65.1888275146484,46.6218643188477,
51.0621528625488,32.7745552062988,
-5.28828430175781,-3.01902484893799,
-58.4293785095215,-14.0220794677734,
-58.8822708129883,11.7396202087402,
-14.5685377120972,41.1633453369141,
25.0622558593750,43.4151763916016,
29.1035404205322,22.7684516906738,
17.4437980651855,6.57047224044800,
20.6591243743897,15.1801090240479,
29.1282730102539,38.2963829040527,
9.05644130706787,46.3794441223145,
-39.4259681701660,25.0485210418701,
-65.3008422851563,-8.42647933959961,
-34.1904144287109,-31.1291713714600,
21.1253376007080,-37.9943389892578,
42.9028778076172,-40.0754165649414,
16.9265384674072,-43.9748153686523,
-16.7529697418213,-35.4832687377930,
-17.1309509277344,-3.88046431541443,
0.783516883850098,28.1753139495850,
4.32895040512085,37.2568893432617,
-9.67903041839600,29.6834392547607,
-21.2243881225586,31.0695381164551,
-17.0699386596680,40.5308341979981,
-8.47014904022217,29.7794284820557,
-2.61835622787476,-9.69881629943848,
10.7741832733154,-38.2734375000000,
30.3603668212891,-19.2812652587891,
32.6814613342285,25.5431709289551,
-0.805503726005554,39.3675231933594,
-39.7184791564941,3.81011605262756,
-37.3442115783691,-35.5679168701172,
14.6053447723389,-27.1790561676025,
64.9281768798828,20.9120178222656,
64.1472244262695,59.2070159912109,
23.2862434387207,51.2187156677246,
-7.21820449829102,11.4497766494751,
-0.783142447471619,-24.4287605285645,
18.3865280151367,-32.7666244506836,
22.2072410583496,-16.1522712707520,
13.2090320587158,4.02214670181274,
7.26903343200684,12.8317441940308,
4.43469333648682,6.92098474502564,
-10.3717231750488,-1.20313453674316,
-37.4356155395508,-4.14807033538818,
-52.0441207885742,-2.37299442291260,
-37.5900726318359,-3.09414601325989,
-16.3702278137207,-4.21621799468994,
-18.2113456726074,-3.62084245681763,
-37.4892044067383,-5.32437705993652,
-33.1314430236816,-16.4394588470459,
11.5007305145264,-30.5872745513916,
61.9067306518555,-28.5782241821289,
60.7159118652344,1.42599630355835,
8.48797798156738,46.3011550903320,
-33.3040847778320,67.0445098876953,
-18.5611248016357,37.8975143432617,
23.9820327758789,-17.2568473815918,
30.4804058074951,-49.1633758544922,
-10.7187700271606,-36.9622802734375,
-45.3909912109375,-14.5469532012939,
-30.8875789642334,-29.7394676208496,
10.0289354324341,-72.9025497436523,
35.6798324584961,-88.9019165039063,
40.2629547119141,-51.0316123962402,
50.2514266967773,-0.396707564592361,
67.6709213256836,12.9824199676514,
65.0803298950195,-5.22835493087769,
35.6778831481934,-15.8874282836914,
6.35288858413696,-9.28603076934815,
-3.44998240470886,-10.7982711791992,
-9.36872005462647,-24.0114345550537,
-28.3095893859863,-18.7569561004639,
-42.8089904785156,16.0683135986328,
-30.3548755645752,39.4237098693848,
-5.35409832000732,13.6771278381348,
7.59187698364258,-37.3082885742188,
13.0623579025269,-57.9567871093750,
30.6585617065430,-38.0417137145996,
55.7294044494629,-16.9929103851318,
57.3785591125488,-18.2765140533447,
28.7157764434814,-20.3262233734131,
2.66158366203308,-6.64494323730469,
2.59834718704224,14.0763559341431,
8.04718875885010,27.5862083435059,
-9.21655941009522,39.8066940307617,
-32.5626564025879,51.5524406433106,
-38.9130630493164,44.1178321838379,
-34.5287170410156,5.33720064163208,
-40.8105125427246,-32.6037178039551,
-47.7791519165039,-26.4487037658691,
-28.9242935180664,10.9024610519409,
6.64951848983765,22.4760761260986,
18.2721843719482,-9.53471565246582,
-9.68263435363770,-40.3699760437012,
-39.9975585937500,-36.5725631713867,
-41.7851486206055,-23.0399417877197,
-33.2035827636719,-32.3518638610840,
-42.8161468505859,-51.6463699340820,
-54.2529563903809,-45.1784515380859,
-26.0021171569824,-23.3710136413574,
28.7829704284668,-25.3287925720215,
59.0298995971680,-49.0456542968750,
43.5844917297363,-42.5076141357422,
20.2702903747559,10.4407510757446,
21.0369529724121,53.8235931396484,
33.5746574401856,32.9723052978516,
23.9966220855713,-21.5835914611816,
-5.25025558471680,-42.5056076049805,
-24.0958042144775,-19.7510242462158,
-14.9562940597534,-0.615792453289032,
8.82619285583496,-13.3838834762573,
29.9235324859619,-27.9003124237061,
39.7184448242188,-12.7481756210327,
28.5616130828857,17.6378936767578,
-9.00798702239990,29.0548572540283,
-49.1844558715820,20.4574317932129,
-63.6534614562988,13.2609338760376,
-52.3218193054199,9.87117862701416,
-42.2578277587891,-2.97636795043945,
-47.3020668029785,-18.5889205932617,
-49.1660194396973,-8.60572338104248,
-28.5499286651611,22.3870258331299,
0.393224149942398,36.6292877197266,
11.7573108673096,12.3577699661255,
3.26255273818970,-26.6257400512695,
-1.02370691299438,-35.8138542175293,
6.83139657974243,-5.49330711364746,
8.06522464752197,28.9353656768799,
-2.86858129501343,32.9502716064453,
-7.20896053314209,9.01283740997315,
12.4383897781372,-16.5948448181152,
41.0053901672363,-21.7666225433350,
49.5467987060547,-4.70078945159912,
27.5836448669434,14.5019636154175,
-7.65680456161499,7.93825721740723,
-34.2733612060547,-24.6678771972656,
-40.9476165771484,-51.5942611694336,
-23.7973136901855,-41.3525009155273,
8.00898742675781,-2.77577614784241,
32.9729995727539,25.3673877716064,
23.1964359283447,21.6690692901611,
-15.5911636352539,6.23297119140625,
-49.0313491821289,6.69433021545410,
-48.2747802734375,16.1755638122559,
-21.2744617462158,7.52708339691162,
3.83538341522217,-18.5980758666992,
19.2337436676025,-33.3617935180664,
37.2583923339844,-20.1736888885498,
58.1298675537109,-2.08910465240479,
61.0166511535645,-6.84204912185669,
32.6240768432617,-27.9716548919678,
-3.74849033355713,-33.8566360473633,
-14.2004566192627,-14.3960886001587,
-3.36869335174561,8.34103679656982,
-7.40610456466675,4.92649126052856,
-41.8396072387695,-22.2125663757324,
-76.8676300048828,-37.5428504943848,
-74.2547760009766,-20.1992244720459,
-32.0935478210449,10.4129972457886,
14.6650714874268,16.5301704406738,
33.7295875549316,-12.2074298858643,
23.6646537780762,-40.5971908569336,
4.28223848342896,-24.7028408050537,
-5.86906003952026,31.0867004394531,
3.84988594055176,68.5059356689453,
25.4671363830566,46.4111595153809,
38.4500350952148,-3.09901762008667,
30.0133686065674,-13.6026506423950,
12.7256917953491,30.6718215942383,
17.1618919372559,72.7799377441406,
40.0449295043945,54.6509056091309,
42.4037475585938,-4.55304241180420,
3.44139099121094,-37.2640838623047,
-43.3859405517578,-22.9090137481689,
-46.2434730529785,-2.60719394683838,
4.55807685852051,-11.7252635955811,
53.7403602600098,-26.7961959838867,
54.5207023620606,-16.5520401000977,
18.8801174163818,1.08251202106476,
-3.37991809844971,-16.4776859283447,
15.0277976989746,-65.3967437744141,
51.9334678649902,-83.8325424194336,
63.3469314575195,-42.6151046752930,
31.3076610565186,7.75149202346802,
-19.7574634552002,8.18535232543945,
-41.5289649963379,-28.1273517608643,
-11.3050327301025,-38.7453956604004,
36.8527832031250,0.352348387241364,
48.8474464416504,45.6666336059570,
9.55236625671387,58.7148857116699,
-35.5886573791504,56.6547431945801,
-40.9667243957520,66.0346832275391,
-13.7768621444702,69.0145187377930,
-2.52617430686951,30.3687000274658,
-17.6959266662598,-36.6497383117676,
-20.1256999969482,-73.4862060546875,
16.1377868652344,-52.3854255676270,
64.3936233520508,-12.8960103988647,
79.3295288085938,-2.34344387054443,
59.6701202392578,-13.2771558761597,
39.4139480590820,-3.49222111701965,
36.2776145935059,31.8664608001709,
28.5790576934814,55.4365768432617,
-4.90436077117920,43.7108001708984,
-47.4742088317871,10.9737415313721,
-68.1131591796875,-10.6516151428223,
-58.4828987121582,-6.95821380615234,
-42.3423767089844,7.57304763793945,
-38.4273185729981,18.2518825531006,
-42.3215675354004,20.2103481292725,
-42.2593574523926,17.0211315155029,
-29.7996215820313,10.7703571319580,
-9.68815612792969,7.45525550842285,
2.77719664573669,6.75746631622314,
-7.07923460006714,2.24229979515076,
-31.2122840881348,-2.11889982223511,
-38.2000885009766,-5.08870315551758,
-8.61013031005859,-16.6501426696777,
41.1180076599121,-45.8906669616699,
59.9008941650391,-75.0119476318359,
30.7241325378418,-68.3887252807617,
-9.34918117523193,-21.8899822235107,
-13.5385761260986,22.2022361755371,
11.3879661560059,16.0129699707031,
19.9592781066895,-26.0451984405518,
-2.99076199531555,-42.3652076721191,
-23.3880233764648,-8.91934108734131,
-15.8082761764526,29.1994876861572,
2.75887274742126,23.5355281829834,
-1.12285137176514,-9.02531147003174,
-19.4473724365234,-18.8243179321289,
-21.8874778747559,6.54750204086304,
-5.91325569152832,33.8472290039063,
-2.55368685722351,39.9197616577148,
-24.7432785034180,33.0329627990723,
-47.1974792480469,24.3790645599365,
-40.8248100280762,4.69830656051636,
-15.6559228897095,-28.7086067199707,
0.396708786487579,-42.8984985351563,
5.44114971160889,-17.6158542633057,
8.79008293151856,19.9386329650879,
9.04247856140137,26.3281536102295,
-0.929095745086670,1.49487352371216,
-20.3262634277344,-11.4551734924316,
-32.0993728637695,1.32177054882050,
-27.7788200378418,12.7681522369385,
-19.1617603302002,5.46916723251343,
-13.4272680282593,1.21939373016357,
0.168469369411469,20.2373504638672,
25.6186237335205,39.3828735351563,
46.7416038513184,26.2828178405762,
54.0874137878418,-6.51128911972046,
51.7472000122070,-10.0790414810181,
38.7784309387207,24.6051616668701,
5.95729970932007,48.5877456665039,
-36.0639724731445,25.3657379150391,
-46.1025886535645,-23.7179374694824,
-0.313135147094727,-56.5587310791016,
60.4444503784180,-58.9329528808594,
66.0042343139648,-44.5842056274414,
12.0917224884033,-27.8841609954834,
-28.3444461822510,-15.7354812622070,
-4.58286952972412,-10.9546928405762,
37.2328109741211,-7.86004829406738,
27.5099945068359,7.67460346221924,
-26.4362678527832,36.7185440063477,
-49.9920539855957,49.8627777099609,
-10.2717361450195,24.4627494812012,
39.1641883850098,-8.37692546844482,
41.6983528137207,6.24605941772461,
3.79611587524414,58.5125465393066,
-23.5585365295410,76.2872848510742,
-28.5374851226807,23.0417175292969,
-32.2453651428223,-47.0240249633789,
-39.3910789489746,-59.3435325622559,
-29.8237972259522,-16.7042827606201,
-1.27185606956482,14.4042530059814,
12.6869249343872,4.77331256866455,
-5.24648809432983,-7.18363523483276,
-30.8724231719971,9.79889774322510,
-32.5657386779785,26.7113590240479,
-9.96685028076172,5.54166936874390,
17.2571506500244,-30.7185420989990,
36.8847122192383,-28.5231113433838,
50.3562431335449,19.6841506958008,
53.4465904235840,58.6805725097656,
31.8683986663818,52.7508621215820,
-5.36529493331909,25.6209793090820,
-27.3868618011475,18.1553897857666,
-21.9247798919678,35.6104621887207,
-6.05366754531860,45.1662483215332,
1.64817309379578,22.9602928161621,
4.99555683135986,-13.5600280761719,
10.6458406448364,-30.1414813995361,
12.0829439163208,-17.8009490966797,
4.06668949127197,10.1041297912598,
-1.16781890392303,28.8579597473145,
9.54016685485840,24.7927246093750,
24.3165264129639,16.9074668884277,
16.5410118103027,27.4458312988281,
-15.2255468368530,46.3373947143555,
-38.8861579895020,33.0460777282715,
-34.4043655395508,-20.1345844268799,
-14.8839979171753,-62.1505126953125,
-7.50731849670410,-36.8070678710938,
-12.5960321426392,40.6450691223145,
-20.3983573913574,85.0330352783203,
-31.7740287780762,50.9635696411133,
-46.8188247680664,-4.78744840621948,
-55.1094512939453,-3.56438064575195,
-42.7889556884766,44.4136695861816,
-16.5873870849609,55.8917808532715,
2.38357949256897,-2.33949184417725,
7.50211381912231,-70.3270492553711,
14.2733745574951,-76.9281387329102,
25.7991085052490,-39.5772972106934,
27.5760326385498,-22.3730373382568,
16.6935749053955,-38.9466400146484,
13.8201951980591,-41.4728775024414,
29.0281581878662,-7.66131973266602,
39.0731124877930,23.6077823638916,
21.7900600433350,13.9259443283081,
-5.79850721359253,-16.4533843994141,
-3.72240328788757,-13.8029603958130,
27.8510494232178,27.9703483581543,
44.9371299743652,59.4782066345215,
20.0134849548340,52.8820571899414,
-13.3022127151489,31.1888217926025,
-6.19494962692261,28.4798183441162,
36.9729347229004,43.9550361633301,
61.3568763732910,47.2012710571289,
33.4873504638672,21.3753147125244,
-15.4386930465698,-4.83468103408814,
-28.4871807098389,-6.82583427429199,
0.938253164291382,3.24475479125977,
30.9650154113770,-4.26679849624634,
23.7126159667969,-29.6221408843994,
-10.7143945693970,-40.8341026306152,
-35.3336753845215,-13.4625997543335,
-30.2189903259277,25.9958038330078,
-14.0032806396484,29.8186492919922,
-5.98431587219238,-2.63700246810913,
-5.34734869003296,-21.3686637878418,
-6.69518995285034,8.82094287872315,
-16.4967803955078,54.6057510375977,
-38.7660942077637,56.9186325073242,
-55.8655357360840,3.06993412971497,
-38.8937110900879,-48.9353294372559,
12.5905275344849,-44.5488433837891,
58.0433235168457,5.81384420394898,
54.5068283081055,44.1687278747559,
10.8197116851807,31.4465026855469,
-22.2426223754883,-13.5950889587402,
-7.32241344451904,-42.0935211181641,
38.2568054199219,-29.9953918457031,
59.3604202270508,8.43045902252197,
26.3078498840332,40.6452560424805,
-31.6387653350830,46.2330741882324,
-64.2047805786133,31.8126678466797,
-47.9190940856934,14.0917167663574,
-7.09789800643921,2.77699422836304,
17.8231105804443,-7.11850929260254,
15.5814037322998,-20.9370002746582,
0.916744709014893,-29.1293411254883,
-8.78329658508301,-13.5022659301758,
-13.7220020294189,23.0627250671387,
-20.8224449157715,50.9048576354981,
-22.6103782653809,36.6954689025879,
-10.1699838638306,-13.6909704208374,
11.8361148834229,-49.0504188537598,
20.2562732696533,-29.9293174743652,
1.96713781356812,25.9703330993652,
-29.1439838409424,64.0157089233398,
-42.4586753845215,49.8940544128418,
-25.1019153594971,13.0303554534912,
11.7835731506348,4.52080154418945,
32.0521087646484,26.4599990844727,
11.8417053222656,42.7130088806152,
-32.9379043579102,31.8886413574219,
-63.8534774780273,13.8710641860962,
-57.2970352172852,10.3337163925171,
-28.9942092895508,7.59165668487549,
-14.1712007522583,-6.50997829437256,
-18.1745758056641,-16.4414443969727,
-13.6742877960205,0.414132773876190,
13.4665870666504,25.9181232452393,
34.5129280090332,16.0209140777588,
25.0383262634277,-30.8560218811035,
10.5714673995972,-61.7822799682617,
28.8885078430176,-35.1634941101074,
71.0748367309570,19.7042388916016,
86.9953689575195,44.4366264343262,
52.2185440063477,28.4918975830078,
6.17285060882568,2.52680516242981,
-5.66904449462891,-9.08630371093750,
2.54636693000793,-2.21920108795166,
-5.53772544860840,21.4174365997314,
-25.2108078002930,54.8384780883789,
-24.2407779693604,72.5767517089844,
-3.96842336654663,47.7154960632324,
-7.40126323699951,-3.24817419052124,
-38.6209182739258,-26.4161643981934,
-44.0590934753418,-7.48229837417603,
3.24062395095825,11.4659852981567,
52.0844650268555,-5.76243400573731,
38.1277923583984,-31.5833568572998,
-17.5487174987793,-20.5314846038818,
-34.3874015808106,8.17381572723389,
12.6284523010254,4.69429874420166,
59.3697967529297,-25.5689163208008,
40.7630653381348,-24.8398990631104,
-14.9264106750488,29.6721401214600,
-41.7235031127930,81.4784927368164,
-21.4905490875244,67.7472381591797,
9.71271038055420,9.43292999267578,
21.1498947143555,-18.3073635101318,
14.5505981445313,12.2454957962036,
-2.28002476692200,61.8686218261719,
-25.5210800170898,77.2381973266602,
-47.3809852600098,50.8444786071777,
-50.2987594604492,5.21041822433472,
-36.1996002197266,-34.1015434265137,
-26.8374786376953,-42.5489845275879,
-30.2691555023193,-11.8560819625855,
-20.9662399291992,28.9760608673096,
12.6122894287109,33.3836326599121,
40.1828193664551,-9.21898174285889,
33.0244064331055,-57.5463066101074,
13.4129629135132,-64.5966720581055,
16.1382350921631,-31.6628017425537,
36.2855415344238,-3.66464400291443,
38.7523117065430,-12.7092065811157,
14.0443458557129,-39.1650581359863,
2.70844292640686,-50.3430633544922,
29.5455722808838,-35.5097122192383,
54.5419273376465,-6.58858919143677,
34.0937957763672,16.4102554321289,
-8.76041030883789,13.7857875823975,
-18.6758728027344,-5.47817897796631,
7.35810279846191,-13.3779354095459,
26.0390987396240,7.86151790618897,
17.5931339263916,32.6977615356445,
14.5473365783691,27.1097698211670,
30.1575775146484,-4.35182905197144,
31.4068412780762,-18.4219360351563,
-1.11330270767212,8.28414916992188,
-29.6735420227051,41.1156730651856,
-6.93170452117920,36.9947395324707,
37.4885635375977,15.4433498382568,
33.8925323486328,21.9436092376709,
-19.2730293273926,46.6260032653809,
-45.8637161254883,32.8144760131836,
-12.5693655014038,-27.2734794616699,
24.6217060089111,-67.3744354248047,
12.1099309921265,-39.6947135925293,
-25.9916763305664,8.52954483032227,
-41.2091598510742,5.27878093719482,
-36.6447601318359,-43.2698745727539,
-42.3211822509766,-60.8517951965332,
-45.2902679443359,-18.0501022338867,
-5.97216129302979,28.2628269195557,
52.5310516357422,27.2776851654053,
58.1049842834473,4.53811168670654,
1.88586640357971,4.57047557830811,
-36.9612731933594,15.5976505279541,
-7.32894134521484,0.467898488044739,
33.5193748474121,-31.2911682128906,
18.4893646240234,-40.9587936401367,
-21.6282119750977,-24.5322380065918,
-11.4011278152466,-18.3481292724609,
42.1309852600098,-26.6095542907715,
60.5561370849609,-6.52269601821899,
14.5812692642212,50.3795471191406,
-30.1521911621094,86.6892242431641,
-12.2450580596924,47.9345359802246,
29.9684982299805,-26.5296878814697,
30.1682262420654,-50.1945762634277,
-13.0695953369141,-11.2301225662231,
-45.8600807189941,22.8625545501709,
-46.2262535095215,6.07037353515625,
-37.4177551269531,-27.6435585021973,
-26.4558486938477,-24.9703884124756,
1.41610693931580,5.88112449645996,
43.8445892333984,16.5360126495361,
69.0466995239258,-5.39919185638428,
58.2374534606934,-18.7257556915283,
32.5323295593262,8.75436210632324,
18.5426368713379,52.9516143798828,
9.36123657226563,71.1110763549805,
-15.2590160369873,51.6540794372559,
-48.2219429016113,16.9835872650147,
-57.5571250915527,-8.86697578430176,
-35.2427902221680,-19.5398521423340,
-9.41333866119385,-17.6708755493164,
-0.200171798467636,-12.8039360046387,
1.43138766288757,-8.87494754791260,
11.6124076843262,-5.38207054138184,
26.5559024810791,0.545357644557953,
27.0447502136230,10.3596105575562,
8.72592830657959,18.4279022216797,
-7.52203989028931,17.2576141357422,
2.56211709976196,10.1864156723022,
31.7024631500244,6.91551113128662,
42.0039634704590,8.00247764587402,
16.2366333007813,5.57819938659668,
-21.8303928375244,-5.90159320831299,
-29.0254211425781,-17.5004272460938,
4.15201568603516,-17.8063774108887,
36.1781005859375,-5.50651645660400,
24.2074413299561,8.65845203399658,
-17.3582153320313,15.6936721801758,
-33.2345733642578,13.1938734054565,
0.614695906639099,8.59164524078369,
45.3771171569824,6.98975944519043,
47.6113586425781,7.80239057540894,
9.97841453552246,5.57404851913452,
-17.4325809478760,-0.730998873710632,
-0.765749692916870,-8.73231697082520,
33.2592163085938,-20.4571475982666,
38.1061325073242,-39.2179260253906,
15.3705148696899,-61.0857925415039,
7.65500307083130,-67.8878021240234,
29.2710990905762,-38.6666679382324,
47.7655715942383,15.7323246002197,
24.5600814819336,54.0833740234375,
-23.9973373413086,43.3139991760254,
-45.1038665771484,1.34823751449585,
-19.5862026214600,-26.1322746276855,
15.0973262786865,-20.7372570037842,
26.9895801544189,-8.57825374603272,
23.8377933502197,-14.0006179809570,
25.8578319549561,-23.6309852600098,
23.4772644042969,-8.58438491821289,
-5.58052682876587,18.6434345245361,
-42.0480346679688,16.3177528381348,
-34.8676605224609,-22.7958507537842,
21.6487503051758,-52.5173873901367,
68.4422378540039,-30.8174190521240,
56.2243881225586,22.6193237304688,
4.61603927612305,58.6226081848145,
-26.3137512207031,53.1586494445801,
-17.4692783355713,33.7587585449219,
-7.13202905654907,21.1211280822754,
-27.6337795257568,6.24747514724731,
-56.2275352478027,-15.3028793334961,
-53.5122337341309,-19.5564327239990,
-18.8041381835938,11.1269044876099,
11.4498128890991,48.8267402648926,
5.18692731857300,47.8084983825684,
-28.1758155822754,6.50529479980469,
-50.2812271118164,-23.8944377899170,
-33.2253379821777,-11.2300357818604,
4.32588338851929,8.82726573944092,
20.0647869110107,-11.1651630401611,
-2.32783317565918,-54.5302200317383,
-31.6836299896240,-59.6140518188477,
-27.3403282165527,-8.59584045410156,
10.8295040130615,40.0253906250000,
35.5817604064941,33.2743721008301,
16.1127166748047,0.105336189270020,
-17.7427387237549,1.98569893836975,
-23.5768680572510,39.8468818664551,
-6.74568700790405,52.2002716064453,
-2.65476846694946,10.1992301940918,
-17.3223094940186,-35.1732940673828,
-17.5600261688232,-27.9619483947754,
13.9961509704590,18.0870742797852,
50.8916091918945,39.2136611938477,
55.3393783569336,16.1069374084473,
32.8492431640625,-7.36115503311157,
6.82144546508789,-0.972847223281860,
-15.3239755630493,18.9523677825928,
-37.4905052185059,23.3651657104492,
-43.4988136291504,12.8836879730225,
-12.0353240966797,6.56599235534668,
36.8820838928223,12.1013050079346,
48.3226966857910,19.8057994842529,
5.07025623321533,21.2343120574951,
-38.6699562072754,20.9519443511963,
-33.6168289184570,20.4492607116699,
-0.223677396774292,22.6234817504883,
5.92811441421509,30.4483451843262,
-30.2777576446533,37.6666450500488,
-63.2583122253418,19.4052257537842,
-58.7210197448731,-30.1233139038086,
-31.8525180816650,-69.7645187377930,
-16.2581844329834,-57.9748382568359,
-11.5235128402710,-2.98329353332520,
-3.98970389366150,41.1166915893555,
-0.579333961009979,41.6234283447266,
-11.6147823333740,18.2834701538086,
-28.1742858886719,5.24907493591309,
-31.7352943420410,3.01902031898499,
-29.0646457672119,-10.1238203048706,
-32.9514923095703,-30.0067501068115,
-34.4178695678711,-34.5566902160645,
-11.6764049530029,-24.6893444061279,
32.6016006469727,-17.7957401275635,
62.6160125732422,-10.6268711090088,
59.6690368652344,14.6868591308594,
44.1906929016113,49.2013168334961,
37.0176467895508,59.8553466796875,
20.1768684387207,36.6866531372070,
-20.1755619049072,14.9007205963135,
-56.7635765075684,20.3970050811768,
-52.5928382873535,26.6165657043457,
-19.7260322570801,-4.73699283599854,
0.840992391109467,-49.1645317077637,
-0.619589328765869,-45.5715255737305,
9.33093070983887,6.83957910537720,
42.9949417114258,39.3485336303711,
61.7474746704102,13.9520215988159,
31.0339069366455,-18.0003223419189,
-23.9498176574707,1.43750035762787,
-52.9470634460449,43.2116851806641,
-43.6950263977051,33.0117034912109,
-27.5057220458984,-33.3811035156250,
-20.7118816375732,-70.6733322143555,
-7.23186445236206,-28.7498664855957,
14.8119440078735,38.9205818176270,
18.1391201019287,49.0041160583496,
-10.5495624542236,0.431980490684509,
-45.2505302429199,-40.4292793273926,
-50.2381744384766,-37.6195182800293,
-17.4184246063232,-18.1318683624268,
21.7526531219482,-7.78186035156250,
37.1022415161133,0.0489756166934967,
22.9993667602539,8.92038345336914,
-2.07726573944092,2.96020579338074,
-14.3707294464111,-25.2983608245850,
-3.34396123886108,-44.5950088500977,
19.5814056396484,-20.5965938568115,
22.8253002166748,28.4749374389648,
-1.89921879768372,51.8730468750000,
-24.5573387145996,27.9979591369629,
-14.0332984924316,-11.8119535446167,
17.1531448364258,-34.9085350036621,
29.3185138702393,-33.9566764831543,
9.19038009643555,-13.0223827362061,
-19.3082504272461,17.8403549194336,
-30.4033203125000,42.3124542236328,
-26.0632362365723,35.4837722778320,
-23.7452087402344,-6.69359683990479,
-15.9758396148682,-47.4648857116699,
9.10713195800781,-47.6957054138184,
35.3972434997559,-13.2647132873535,
32.2443389892578,13.3081502914429,
-3.04111790657043,4.60316658020020,
-38.1427536010742,-22.3497638702393,
-45.9573783874512,-33.9401817321777,
-36.4530181884766,-25.4704132080078,
-30.9414520263672,-11.3742904663086,
-25.4728374481201,0.226104736328125,
-3.38314247131348,11.8452930450439,
27.5775508880615,30.6955623626709,
33.1561889648438,46.9234924316406,
-1.74614691734314,46.4758491516113,
-45.5356750488281,24.8815536499023,
-55.1101646423340,1.34648692607880,
-30.2721977233887,-1.96627116203308,
-10.5972127914429,12.7498893737793,
-23.4917354583740,21.5372772216797,
-51.6064872741699,6.43351078033447,
-61.5387802124023,-20.6394939422607,
-42.7576217651367,-21.9996185302734,
-13.2240409851074,11.7940845489502,
7.13163805007935,41.3106384277344,
12.8861713409424,27.2060909271240,
7.21158409118652,-18.2364654541016,
-9.26398468017578,-44.7282028198242,
-28.1137771606445,-32.3379325866699,
-36.5047302246094,-14.6518707275391,
-26.7058658599854,-27.8685760498047,
-5.58296871185303,-55.9723625183106,
16.9119968414307,-50.2955169677734,
28.4341201782227,-8.11671257019043,
20.4962100982666,21.6010932922363,
-2.63360881805420,2.82002544403076,
-22.2021064758301,-40.0770492553711,
-15.3477497100830,-61.5228805541992,
16.4485511779785,-50.7002525329590,
42.5352935791016,-36.8299293518066,
35.6215896606445,-36.9189071655273,
10.1769523620605,-36.2698860168457,
-3.61433863639832,-28.0698223114014,
1.46848726272583,-26.9522819519043,
6.12284517288208,-40.4476318359375,
-2.89274024963379,-48.3910484313965,
-6.26690244674683,-25.4064826965332,
13.1195993423462,15.1014633178711,
40.2771453857422,33.2341156005859,
45.7376670837402,13.0759544372559,
24.7693099975586,-10.4452724456787,
5.27050161361694,0.942154645919800,
8.74847030639648,36.8988265991211,
23.2037620544434,53.4394569396973,
23.2918643951416,26.4529209136963,
7.68435668945313,-16.2085189819336,
-1.83600592613220,-26.4399166107178,
6.91370010375977,2.77756786346436,
17.4379806518555,34.9905281066895,
6.83914661407471,34.4617271423340,
-25.8969154357910,8.79118728637695,
-51.6186065673828,-12.9073534011841,
-44.0910453796387,-18.5370941162109,
-4.66074943542481,-19.8620471954346,
35.8782768249512,-23.9859790802002,
44.8438186645508,-14.4775695800781,
18.9163627624512,18.8053245544434,
-17.5002117156982,51.7647666931152,
-27.5402336120605,50.2065277099609,
-4.08666324615479,18.5284118652344,
22.8796768188477,-1.88900518417358,
26.0275859832764,9.29118251800537,
14.7608404159546,24.3506736755371,
15.2739744186401,9.49761772155762,
33.2623634338379,-23.5786666870117,
42.2566947937012,-33.2359237670898,
19.7697257995605,-8.90574836730957,
-17.7660312652588,11.0419311523438,
-36.7649765014648,-4.30234909057617,
-31.7742843627930,-40.2834739685059,
-17.7998600006104,-61.9459190368652,
6.38029766082764,-59.2669601440430,
36.8002052307129,-47.1504249572754,
50.0900573730469,-32.1689071655273,
19.6656093597412,-8.94394302368164,
-31.7452602386475,12.5684871673584,
-43.2454490661621,6.02764415740967,
2.15525531768799,-26.1004047393799,
43.7537307739258,-47.9842948913574,
25.7502746582031,-33.5892677307129,
-23.9757461547852,-3.27262473106384,
-34.7083778381348,2.93504786491394,
-3.05548167228699,-20.6329345703125,
8.97902393341065,-36.1933403015137,
-25.8904285430908,-19.1764602661133,
-45.8264007568359,9.85942554473877,
-0.934930801391602,22.4619083404541,
66.1248550415039,13.5378541946411,
76.6374893188477,-0.505671977996826,
23.6815414428711,-9.38611793518066,
-25.1832122802734,-9.98165798187256,
-19.7287311553955,0.863186001777649,
16.6198234558105,17.1745967864990,
32.6905822753906,18.8930187225342,
18.1468620300293,-5.05247354507446,
2.98244285583496,-29.1304092407227,
6.94944858551025,-13.9691638946533,
23.5565528869629,34.7164840698242,
38.0199890136719,56.7433547973633,
30.5349979400635,19.5827579498291,
-6.73266220092773,-32.5657272338867,
-46.6068305969238,-33.2405929565430,
-50.4691390991211,20.2068386077881,
-19.6767826080322,62.7107925415039,
-2.67152905464172,46.3908920288086,
-27.7015151977539,-3.70836639404297,
-59.1765136718750,-36.1144790649414,
-46.0399436950684,-38.6018104553223,
3.96261072158813,-30.9527492523193,
25.4994201660156,-21.6867351531982,
-4.11940670013428,-1.13748037815094,
-27.7289352416992,22.1012420654297,
-1.92787146568298,18.1908512115479,
38.3638305664063,-12.9533624649048,
37.5379562377930,-29.1403293609619,
4.04635047912598,-1.49590063095093,
-6.49733972549439,44.1024322509766,
20.7158813476563,59.5070533752441,
38.3687477111816,28.7769184112549,
17.8687973022461,-11.6061897277832,
-7.10907697677612,-17.5305023193359,
-3.70070648193359,6.30632352828980,
9.71210765838623,24.9635086059570,
-1.73846077919006,13.5155820846558,
-21.2905464172363,-19.7710781097412,
-3.43485999107361,-39.9127464294434,
45.7984504699707,-19.5343456268311,
61.0881462097168,21.9891071319580,
15.9803047180176,39.5094146728516,
-41.2782821655273,12.7098999023438,
-50.5273857116699,-20.5723857879639,
-14.1917247772217,-14.2327804565430,
14.6800994873047,23.4286575317383,
3.57337474822998,33.0761985778809,
-25.0495243072510,-14.0295267105103,
-37.6427688598633,-69.8925476074219,
-27.2243499755859,-65.9346542358398,
-9.30999755859375,-5.09542274475098,
2.90866327285767,44.3252716064453,
1.03909218311310,41.8583030700684,
-14.6328954696655,14.3334541320801,
-26.3576450347900,10.9439363479614,
-9.61806488037109,33.6089973449707,
26.9318447113037,47.2717170715332,
45.9651374816895,35.5586662292481,
27.8275756835938,21.6525764465332,
-7.61967039108276,24.1410598754883,
-22.6134586334229,36.0638542175293,
-5.25425863265991,35.7471656799316,
16.1219310760498,21.2963104248047,
22.1377696990967,0.617874026298523,
18.4188861846924,-23.4473762512207,
16.0647106170654,-48.6088180541992,
15.8657398223877,-57.3949165344238,
17.6442871093750,-29.8182601928711,
20.4365024566650,19.7527999877930,
16.0121364593506,54.2164878845215,
-10.0273895263672,54.2099342346191,
-48.0860137939453,33.2106819152832,
-62.8387565612793,21.7867259979248,
-31.7693138122559,26.6778202056885,
12.3069124221802,33.7384948730469,
17.4726200103760,35.7568969726563,
-23.3245067596436,43.3566474914551,
-62.2289886474609,56.5441398620606,
-56.7237777709961,57.3609237670898,
-20.1579208374023,33.9762916564941,
7.98595714569092,-4.79121208190918,
10.7395906448364,-31.2280025482178,
-1.66269171237946,-26.7750396728516,
-21.1835079193115,-4.32117271423340,
-48.8679199218750,8.40508651733398,
-68.8862075805664,-9.69431400299072,
-58.4956665039063,-44.7681770324707,
-12.9110889434814,-61.8576850891113,
33.1882934570313,-40.2872238159180,
46.9756469726563,1.83007025718689,
29.2991733551025,17.7290515899658,
7.86062955856323,-6.80151748657227,
0.746524035930634,-36.5226631164551,
-0.689839243888855,-28.6254158020020,
-4.75628280639648,10.8948936462402,
-12.2300968170166,34.5873031616211,
-22.9192276000977,16.0180702209473,
-29.8895206451416,-25.7865066528320,
-18.3551940917969,-48.3694992065430,
16.2519721984863,-38.2699966430664,
53.2369842529297,-10.1864929199219,
58.7428474426270,20.5206375122070,
20.4510555267334,44.6672477722168,
-25.8085021972656,50.7062988281250,
-47.2357978820801,28.5702934265137,
-46.2279586791992,-9.35912036895752,
-46.2128448486328,-33.5343666076660,
-44.0318794250488,-25.8172836303711,
-18.0009193420410,-5.52065277099609,
23.7179126739502,0.739524245262146,
42.2426414489746,-7.21847772598267,
21.5441150665283,-8.66931343078613,
2.31133651733398,10.3335475921631,
22.1830768585205,35.5117034912109,
54.0841140747070,44.8551902770996,
37.7807693481445,32.3583374023438,
-34.2950782775879,13.1687841415405,
-96.6941757202148,-2.31503415107727,
-89.9935989379883,-7.34151983261108,
-32.6505889892578,-4.73816442489624,
5.01049232482910,-2.18695592880249,
-4.30776739120483,-5.20635890960693,
-25.1146144866943,-10.5972204208374,
-15.2421312332153,-7.18244504928589,
18.1891365051270,8.51951503753662,
32.7421607971191,21.6436424255371,
6.42070055007935,14.7927465438843,
-33.6546096801758,-9.56311702728272,
-40.5768165588379,-29.2397708892822,
-6.54798126220703,-33.6906967163086,
33.0193634033203,-37.1335144042969,
41.9395294189453,-51.7237243652344,
20.4851360321045,-60.7279090881348,
-1.80647504329681,-45.5562171936035,
-1.71529519557953,-13.6171388626099,
15.8512077331543,1.07349956035614,
28.6901397705078,-11.7970619201660,
39.2791633605957,-19.7721786499023,
49.7748374938965,4.00338459014893,
42.0045471191406,40.1036872863770,
-4.14956474304199,45.5325927734375,
-64.0284500122070,13.8254299163818,
-82.5528259277344,-16.0786533355713,
-30.6460094451904,-12.9667940139771,
41.5522880554199,6.40041637420654,
58.0222206115723,8.69848728179932,
12.4698200225830,-4.14929103851318,
-29.1075744628906,-4.34749460220337,
-25.0732765197754,21.3823814392090,
-8.37129688262940,48.6787872314453,
-30.4134254455566,44.2686157226563,
-67.7400665283203,5.56772994995117,
-58.3138885498047,-32.7297248840332,
-1.35449481010437,-38.9474143981934,
30.3178195953369,-16.1564407348633,
-5.79376745223999,3.03573203086853,
-57.0440330505371,-4.89443540573120,
-42.9468116760254,-27.6951427459717,
26.8646831512451,-30.1677379608154,
72.5764312744141,-0.949624061584473,
52.2704162597656,25.4146919250488,
8.33607769012451,13.1541833877563,
-0.806267917156220,-20.5799160003662,
22.0405063629150,-28.3586025238037,
40.4622840881348,5.92797279357910,
45.1467399597168,43.7849311828613,
43.9280700683594,44.4621696472168,
36.7119941711426,18.1663341522217,
13.0435476303101,2.92727923393250,
-15.1658220291138,6.51855707168579,
-18.2969570159912,3.04498410224915,
9.92682838439941,-14.1663436889648,
36.4506072998047,-17.6724777221680,
33.4584693908691,9.21864128112793,
9.16576576232910,41.5739135742188,
-10.0830402374268,48.0985488891602,
-18.3368511199951,32.4262733459473,
-19.7594623565674,26.9036026000977,
-12.5488929748535,38.0530662536621,
-0.651236057281494,41.1937675476074,
2.49636578559876,22.1157169342041,
-14.2041034698486,-2.76237630844116,
-35.1441574096680,-16.3165321350098,
-32.5320243835449,-25.4172286987305,
1.73571503162384,-41.4390830993652,
40.7447624206543,-46.3972129821777,
46.7168693542481,-16.6751041412354,
14.1392288208008,29.6528091430664,
-28.0056438446045,45.7872619628906,
-45.9195480346680,16.2471313476563,
-24.7329673767090,-18.0373535156250,
14.9825725555420,-12.7741508483887,
32.7763137817383,21.7563266754150,
13.6528987884521,40.0659561157227,
-13.1808748245239,22.3307952880859,
-12.2134456634521,-0.121547713875771,
11.1180686950684,-2.14740681648254,
10.3851671218872,6.64719676971436,
-33.0439033508301,6.00805330276489,
-74.8747940063477,-3.92744684219360,
-60.6256408691406,-12.3664789199829,
0.592039585113525,-19.8465976715088,
43.0961227416992,-30.7843761444092,
22.8130798339844,-35.3447761535645,
-29.4937343597412,-19.2942771911621,
-53.4399185180664,6.87067747116089,
-33.0615196228027,19.5021533966064,
-4.39104032516480,12.7426366806030,
-1.60388112068176,7.25214147567749,
-17.6619606018066,10.0425920486450,
-22.6081943511963,-0.556715726852417,
-1.85261416435242,-28.4063014984131,
26.8109073638916,-39.2505264282227,
33.9714660644531,-8.67696952819824,
10.5105113983154,36.2378921508789,
-15.9832944869995,47.8016700744629,
-14.1787767410278,22.1633796691895,
17.0187931060791,4.58705043792725,
38.6288871765137,22.1650733947754,
13.3803215026855,51.3482398986816,
-36.6981620788574,56.9993247985840,
-48.1563987731934,39.7696151733398,
-3.04854559898376,20.5675792694092,
44.1353607177734,1.40628516674042,
37.7669219970703,-24.2775878906250,
-7.82866573333740,-40.1458053588867,
-28.3289470672607,-29.2600784301758,
0.00947606563568115,-3.14603233337402,
29.5053901672363,9.85964298248291,
20.7739791870117,5.80710744857788,
7.65886211395264,4.00320768356323,
35.5618972778320,13.3898677825928,
76.2827301025391,21.0345821380615,
60.0199317932129,19.3372287750244,
-15.0640363693237,24.2210960388184,
-64.2734527587891,39.1895027160645,
-30.8670501708984,40.4007568359375,
33.8053436279297,15.3588390350342,
44.2142562866211,-3.62666082382202,
1.34779644012451,12.6974754333496,
-17.8102626800537,43.0979232788086,
19.7677478790283,39.8822059631348,
55.7808418273926,5.53459930419922,
35.2906951904297,-7.93334865570068,
-14.4198493957520,21.3456115722656,
-29.8365345001221,54.6846885681152,
-6.06685352325439,45.6460304260254,
13.8439226150513,6.43639898300171,
13.9781503677368,-9.32793807983398,
13.2131357192993,17.7741966247559,
18.5370101928711,55.4565315246582,
7.40712261199951,63.8829612731934,
-20.6014556884766,41.1839103698731,
-27.5557575225830,8.92085266113281,
10.3391084671021,-7.96365785598755,
49.1998405456543,-0.369946956634522,
32.7374725341797,19.3317642211914,
-27.7021198272705,24.4326400756836,
-69.6761779785156,4.08304166793823,
-64.3234329223633,-19.2434844970703,
-38.0109291076660,-19.7010421752930,
-24.7555065155029,-2.96219801902771,
-28.0981082916260,-0.679850459098816,
-37.2464637756348,-24.4824428558350,
-48.6153259277344,-46.8500976562500,
-56.1780204772949,-39.0523757934570,
-38.1728477478027,-17.4176731109619,
6.99279689788818,-16.8195419311523,
37.6464080810547,-38.4287719726563,
16.1389045715332,-49.5212135314941,
-36.9008750915527,-37.6044540405273,
-58.3555068969727,-19.1542797088623,
-32.8405456542969,-14.8290452957153,
-8.25741863250732,-16.1661891937256,
-20.6550788879395,-9.97881889343262,
-50.8389930725098,-1.48155355453491,
-55.0533485412598,-2.44973707199097,
-30.1751194000244,-11.8734846115112,
-12.2081241607666,-14.8234405517578,
-17.4630279541016,-9.09302234649658,
-22.6051673889160,-6.79158878326416,
-1.92703652381897,-10.3977651596069,
31.4736766815186,-8.90140724182129,
48.9947738647461,0.131898924708366,
33.3071098327637,-0.166122496128082,
-5.80329847335815,-16.3426761627197,
-47.2772445678711,-34.8323898315430,
-64.6696014404297,-38.4727058410645,
-42.7576980590820,-33.2486152648926,
3.66010355949402,-33.2175140380859,
41.9625320434570,-32.3981590270996,
54.0607452392578,-8.49257946014404,
50.5000648498535,31.8723278045654,
47.8452186584473,53.9942398071289,
45.0650177001953,37.1671981811523,
24.5243186950684,6.37125492095947,
-11.4463605880737,-3.80396437644959,
-40.4416961669922,0.115794613957405,
-48.5667572021484,-15.3488473892212,
-41.8890419006348,-49.9343299865723,
-29.2464828491211,-59.9489555358887,
-10.3993854522705,-20.5352096557617,
12.1759443283081,29.4983711242676,
23.8091964721680,31.1705284118652,
13.3862075805664,-11.8668498992920,
-6.65014505386353,-39.0037803649902,
-13.5407228469849,-6.92568159103394,
-4.91889476776123,51.3192634582520,
1.33507955074310,73.5971679687500,
-7.76352453231812,46.5478820800781,
-19.4830150604248,8.65331268310547,
-13.9273223876953,-2.94369149208069,
12.9578037261963,10.1089620590210,
37.7974166870117,24.2010440826416,
35.5686264038086,25.6230964660645,
3.87661695480347,16.4709377288818,
-32.6362800598145,-1.00082540512085,
-44.0768318176270,-22.3792400360107,
-25.2950897216797,-32.3422584533691,
2.73391342163086,-13.7208051681519,
13.0299615859985,24.4849948883057,
1.82698488235474,53.0938186645508,
-16.7546119689941,48.3999710083008,
-31.6585311889648,16.4253749847412,
-37.7006263732910,-13.9889011383057,
-31.9700584411621,-25.6521263122559,
-15.2295246124268,-26.3685951232910,
2.69627881050110,-29.4534301757813,
4.18840408325195,-38.4147605895996,
-7.14458417892456,-42.2456016540527,
-6.39401626586914,-33.2559089660645,
20.3392276763916,-13.6421012878418,
45.5385475158691,9.90638923645020,
34.3827629089356,35.6625938415527,
-11.7842655181885,56.1714019775391,
-50.4184455871582,63.0282554626465,
-42.1771888732910,56.5426597595215,
-3.94681334495544,44.5401954650879,
18.8947772979736,31.8103618621826,
4.30626344680786,12.4643774032593,
-22.7251567840576,-18.9696903228760,
-21.1250591278076,-41.6960945129395,
15.4918594360352,-33.6108627319336,
50.9042701721191,2.09425401687622,
54.3790168762207,26.9770660400391,
33.9267578125000,18.2745761871338,
22.2896251678467,-0.697627723217011,
32.4560737609863,5.99238300323486,
36.9535865783691,31.6068058013916,
9.57180213928223,38.3453407287598,
-31.5992317199707,7.73866415023804,
-46.9209861755371,-31.3244667053223,
-20.3521881103516,-42.4785041809082,
22.4940834045410,-32.5235404968262,
40.9476051330566,-28.0692272186279,
22.9473247528076,-37.4052696228027,
-10.5230646133423,-42.5631599426270,
-29.4712924957275,-40.1435546875000,
-13.0858230590820,-40.8619499206543,
28.3282661437988,-45.0759086608887,
52.0052680969238,-29.7339553833008,
24.8161811828613,8.71004486083984,
-33.6164016723633,35.0114669799805,
-56.7402000427246,18.4842967987061,
-13.9096212387085,-22.0361671447754,
45.4099121093750,-36.1530227661133,
45.1215591430664,-7.61052322387695,
-17.7527141571045,25.9689865112305,
-67.6215667724609,25.5660171508789,
-47.5879898071289,-1.47723710536957,
8.21674823760986,-18.4341583251953,
23.6545448303223,-12.8357677459717,
-17.9434051513672,-2.21543908119202,
-57.5261383056641,-7.19213867187500,
-47.0713119506836,-24.4455299377441,
-4.14303493499756,-43.6786270141602,
22.7889823913574,-52.8319931030273,
20.4399185180664,-48.7593994140625,
17.0379238128662,-33.1696128845215,
26.1693706512451,-12.1319684982300,
27.7544174194336,5.88716411590576,
5.33760833740234,7.41111850738525,
-23.3308334350586,-9.26156425476074,
-24.9891929626465,-31.6209831237793,
5.59735965728760,-44.3312530517578,
37.3230895996094,-33.6473541259766,
45.7016181945801,-5.64872455596924,
40.3154678344727,12.4677124023438,
34.4571838378906,8.81775379180908,
28.9962882995605,3.18608713150024,
14.8884611129761,23.1367492675781,
-3.51078462600708,55.9017601013184,
-11.6721763610840,56.5217590332031,
1.43562459945679,6.33885526657105,
22.2983970642090,-47.1298522949219,
29.7602043151855,-41.1279029846191,
22.2491989135742,15.8102426528931,
11.5823135375977,51.7188186645508,
9.06641674041748,19.2605705261230,
11.4083328247070,-40.6327819824219,
5.17357492446899,-57.2673187255859,
-14.7827367782593,-18.2600421905518,
-33.4886627197266,31.9592056274414,
-35.7700767517090,50.5926704406738,
-31.7326431274414,46.5680847167969,
-37.1906013488770,38.7633705139160,
-51.4323539733887,21.4764347076416,
-47.4306526184082,-13.0114803314209,
-12.8217782974243,-46.6562995910645,
23.0061111450195,-49.5976562500000,
15.7377767562866,-25.5441589355469,
-29.0117740631104,-5.15880012512207,
-60.4921302795410,-6.75985145568848,
-41.3329582214356,-10.1887006759644,
2.53691816329956,6.70754241943359,
17.3536224365234,24.7562427520752,
-5.12236356735230,9.61837673187256,
-21.1979198455811,-38.7038917541504,
3.89107108116150,-78.9721374511719,
48.0694198608398,-73.2454986572266,
60.0061683654785,-28.6057262420654,
26.4545078277588,14.7240982055664,
-14.3264970779419,36.2943725585938,
-18.9875373840332,42.4109115600586,
5.28033924102783,45.0127639770508,
15.9011573791504,36.8505287170410,
-17.5511913299561,9.82651329040527,
-67.9477615356445,-16.9259796142578,
-83.8234405517578,-17.3300209045410,
-47.4902305603027,5.53941679000855,
9.56994915008545,17.1646099090576,
44.0677413940430,-3.22100257873535,
36.8055000305176,-29.1488704681397,
9.93166351318359,-22.8695621490479,
-9.49359130859375,13.0398540496826,
-13.5974321365356,42.4817771911621,
-4.69549798965454,45.1456336975098,
9.19696140289307,32.0253295898438,
10.7145853042603,20.0387535095215,
-11.6023769378662,1.94486629962921,
-46.4161872863770,-25.7779560089111,
-64.6898803710938,-40.0464439392090,
-51.2316932678223,-23.2082519531250,
-29.9321174621582,5.01657199859619,
-30.0504016876221,8.67919540405273,
-39.7865486145020,-17.3315467834473,
-17.6952381134033,-41.6459617614746,
38.0928688049316,-43.4730606079102,
75.5611877441406,-27.9599781036377,
49.5136146545410,-10.3446426391602,
-12.1965370178223,6.82063627243042,
-39.0456123352051,21.3401546478272,
-12.0434341430664,21.2331600189209,
16.8022918701172,4.19587373733521,
2.36008191108704,-7.94690275192261,
-38.3513336181641,-1.51735079288483,
-54.1829528808594,5.85754299163818,
-30.1645679473877,-12.1298141479492,
1.86195886135101,-44.5947952270508,
18.6485671997070,-57.2666320800781,
24.4573135375977,-34.6234626770020,
31.2267055511475,4.13670301437378,
28.4391155242920,33.7908287048340,
8.44011402130127,47.5109405517578,
-18.8922882080078,50.3791084289551,
-34.0043716430664,40.3521232604981,
-31.9551925659180,19.8074836730957,
-17.3741416931152,4.00054073333740,
11.6626815795898,2.57571744918823,
47.7510604858398,2.44259381294251,
64.8232040405273,-10.3977489471436,
41.7025413513184,-19.5844860076904,
-8.46955108642578,-0.00692558288574219,
-43.3187675476074,39.6235656738281,
-36.4628295898438,62.3983497619629,
-10.6181631088257,50.2483825683594,
-4.19536590576172,27.0721454620361,
-21.2014884948730,24.0083503723145,
-36.1510658264160,37.4228096008301,
-29.5054645538330,36.3069801330566,
-8.69931697845459,9.85497570037842,
3.14921092987061,-21.8383388519287,
-2.62245798110962,-41.6719322204590,
-11.0803718566895,-48.2781791687012,
1.54147005081177,-41.5041465759277,
34.7032127380371,-18.9980716705322,
62.9167823791504,7.84206151962280,
50.2765998840332,14.3233060836792,
2.66668701171875,-5.06771087646484,
-31.2409286499023,-24.4279785156250,
-8.14594459533691,-15.9349737167358,
52.5323944091797,15.2276058197021,
79.2362670898438,36.6131553649902,
35.6676101684570,31.8708305358887,
-31.8758811950684,12.6173629760742,
-51.3386802673340,-10.0956077575684,
-11.3546943664551,-35.0643920898438,
36.3301200866699,-50.6610870361328,
42.3401184082031,-30.4666271209717,
21.3554096221924,21.8047637939453,
18.1501216888428,61.9592056274414,
41.6940841674805,56.5094871520996,
63.8830642700195,23.6894130706787,
55.9954147338867,10.0549736022949,
20.3534317016602,23.9928417205811,
-19.1090888977051,26.9627132415772,
-38.9008140563965,-5.66039562225342,
-23.2945346832275,-48.1100502014160,
17.8648338317871,-63.1717491149902,
46.0870590209961,-52.9027404785156,
27.9391002655029,-38.2589759826660,
-17.2498416900635,-26.4735736846924,
-37.7286949157715,-13.8600378036499,
-7.11739587783814,-6.26161718368530,
37.1714668273926,-13.1285810470581,
35.6170501708984,-19.6065406799316,
-12.2496509552002,-0.713779568672180,
-55.8882751464844,28.2977809906006,
-63.4043731689453,26.6290378570557,
-48.4878044128418,-15.8833293914795,
-34.1823120117188,-57.5927581787109,
-14.1121788024902,-47.4084396362305,
17.0594844818115,-2.04471087455750,
36.2887420654297,17.7921733856201,
19.8516483306885,-12.0567398071289,
-8.56746196746826,-56.8016738891602,
-5.33868408203125,-68.4402313232422,
28.3851089477539,-33.0968055725098,
41.8273735046387,15.6143283843994,
0.928720712661743,37.7182350158691,
-52.5367088317871,19.5418834686279,
-52.6982650756836,-14.0291137695313,
0.620616436004639,-22.9881248474121,
45.5233573913574,5.93802213668823,
36.7555503845215,37.0962753295898,
-9.68840503692627,21.7603454589844,
-38.6707000732422,-37.9187622070313,
-19.9198265075684,-79.9562225341797,
20.3495502471924,-49.5596313476563,
41.0642280578613,22.8199501037598,
22.7685985565186,58.7707099914551,
-10.9751777648926,31.8634681701660,
-18.9045486450195,-10.8319807052612,
12.0965204238892,-18.3172111511230,
47.1350860595703,6.28411912918091,
41.0854568481445,18.5896205902100,
-6.86106681823731,8.37504673004150,
-43.3906440734863,6.64218902587891,
-34.8240699768066,25.0870761871338,
-9.39612483978272,42.4603080749512,
-14.1207380294800,38.4020729064941,
-48.8272209167481,19.3940696716309,
-62.2943649291992,-0.383631944656372,
-22.3895664215088,-25.7153949737549,
35.8022155761719,-53.6867942810059,
53.3216056823731,-56.0706748962402,
19.0819702148438,-19.1307411193848,
-27.1646537780762,19.5607719421387,
-42.0049667358398,10.0988340377808,
-19.8378982543945,-40.4355812072754,
16.4584217071533,-64.0745239257813,
45.0595130920410,-19.4224281311035,
52.3171157836914,48.3585891723633,
38.9475555419922,70.7120285034180,
20.0894966125488,35.7326126098633,
6.31195116043091,-10.3659820556641,
-3.10654997825623,-26.5221061706543,
-11.0057849884033,-9.61773300170898,
-14.7901105880737,26.2312431335449,
-7.99420547485352,59.2400131225586,
5.33000993728638,62.5339851379395,
12.1324462890625,19.6500129699707,
9.33164787292481,-42.2126083374023,
17.0700645446777,-62.9226760864258,
40.9243316650391,-24.1783733367920,
45.5732688903809,26.4491405487061,
6.78991127014160,27.3739776611328,
-46.9079093933106,-19.4847526550293,
-56.1660156250000,-56.5634307861328,
-8.87784194946289,-55.0570297241211,
37.3917503356934,-30.4476642608643,
32.6354866027832,-6.61835527420044,
-0.224757328629494,4.64838409423828,
-3.79315471649170,3.26222443580627,
25.0669574737549,-12.8072204589844,
35.0938186645508,-36.2122879028320,
7.00080633163452,-41.9166145324707,
-13.4822111129761,-19.3263263702393,
5.96012306213379,11.9591703414917,
30.9085884094238,31.1659431457520,
9.41056728363037,36.5296707153320,
-41.9250793457031,37.4467926025391,
-57.2120246887207,19.6302890777588,
-20.7627105712891,-27.5300521850586,
12.4160461425781,-71.0448608398438,
0.386167049407959,-61.6772460937500,
-30.2704067230225,-7.25811910629273,
-33.5175857543945,37.0784835815430,
-15.8865337371826,30.0762157440186,
-11.6028289794922,-8.37515544891357,
-13.3704433441162,-34.7052383422852,
12.6851587295532,-36.3146286010742,
55.7121505737305,-27.7312450408936,
60.9209175109863,-10.5808734893799,
12.5696811676025,17.1886024475098,
-39.3958168029785,28.1018238067627,
-39.6720237731934,-8.73466110229492,
3.44105720520020,-65.0226364135742,
38.0831680297852,-76.3421859741211,
39.4969100952148,-36.3498802185059,
29.7999191284180,-8.62335968017578,
29.3261547088623,-35.3609771728516,
30.5087833404541,-67.0750808715820,
24.4782848358154,-38.0718612670898,
10.7896509170532,26.7595844268799,
-11.1182193756104,41.7660255432129,
-28.9423847198486,-10.1917791366577,
-22.3256263732910,-44.3508682250977,
11.7328681945801,-6.87618398666382,
42.6158332824707,46.0639724731445,
36.5419158935547,37.3219223022461,
5.14878368377686,-16.5290737152100,
-6.42053508758545,-35.0842742919922,
16.8653964996338,-2.52894115447998,
29.1880245208740,16.3697090148926,
-2.15005111694336,-12.1349849700928,
-40.0570068359375,-39.7885208129883,
-29.2561454772949,-13.9748992919922,
12.8465347290039,41.4416427612305,
16.5384922027588,60.2185363769531,
-31.1531982421875,31.1144981384277,
-63.5204200744629,7.36247014999390,
-28.2327175140381,20.2849273681641,
34.4949951171875,45.6233100891113,
46.5275039672852,48.8245773315430,
-0.680201053619385,24.0095310211182,
-39.3809356689453,-8.47274398803711,
-21.9863395690918,-24.4343757629395,
20.4066162109375,-9.09559631347656,
29.2125396728516,27.0107975006104,
-5.59350728988648,50.7161178588867,
-47.9858169555664,32.9710464477539,
-62.2006034851074,-15.8912506103516,
-41.1037979125977,-45.7769699096680,
4.73082542419434,-26.7741260528564,
45.9549598693848,8.51641368865967,
50.3976516723633,9.18955802917481,
14.7912960052490,-18.7852916717529,
-22.1316223144531,-30.3061542510986,
-21.0617542266846,-8.73110389709473,
14.6612224578857,19.1215610504150,
36.1985321044922,29.7018909454346,
12.5151453018188,26.5827903747559,
-25.3679332733154,23.9142189025879,
-34.6796493530273,16.0234985351563,
-15.1014328002930,2.09514808654785,
3.87029480934143,4.11370611190796,
4.83718013763428,33.2684936523438,
-9.73601818084717,54.7408218383789,
-28.9323501586914,30.1567020416260,
-44.8995971679688,-17.9766693115234,
-47.7997016906738,-25.6856651306152,
-29.3516960144043,18.3167896270752,
-9.03329086303711,51.3883132934570,
-11.4659214019775,28.3809375762939,
-28.0047893524170,-12.3484191894531,
-22.2741928100586,-10.6447906494141,
17.5515327453613,26.5997562408447,
47.2630004882813,41.6453819274902,
30.3267211914063,16.0346202850342,
-6.74050235748291,-1.33213257789612,
-9.35645103454590,16.0315799713135,
27.0086364746094,31.2400188446045,
52.0846862792969,2.91361808776855,
31.7657127380371,-40.9712409973145,
-7.16154193878174,-44.8312110900879,
-20.0471210479736,-8.15591907501221,
-1.72022199630737,16.7274112701416,
16.5174770355225,2.52962613105774,
22.6048851013184,-23.1229019165039,
22.6797180175781,-27.6722621917725,
19.4370040893555,-12.1721534729004,
-0.616637945175171,1.95833373069763,
-32.0258293151856,13.3004989624023,
-50.2776870727539,29.7820529937744,
-40.4414901733398,44.7004737854004,
-16.7788810729980,43.7618522644043,
1.88150155544281,33.9873237609863,
12.0068988800049,28.6976413726807,
15.0655622482300,24.6126461029053,
9.14743804931641,7.69768810272217,
-8.48290443420410,-15.2163524627686,
-21.7760219573975,-19.5249156951904,
-5.55139875411987,1.01301229000092,
31.0368022918701,26.2971477508545,
52.2796745300293,34.3374099731445,
44.0849456787109,29.8993682861328,
29.9509601593018,33.5514907836914,
30.8389472961426,49.2038192749023,
39.4052925109863,59.2597732543945,
34.6139030456543,50.0180244445801,
19.4184951782227,28.1030387878418,
7.16567754745483,10.6909294128418,
-8.83624553680420,6.76327800750732,
-44.9980697631836,15.5012836456299,
-80.7992935180664,17.4442958831787,
-69.0497360229492,-1.75987958908081,
-9.31916427612305,-28.9363346099854,
33.3614692687988,-33.1805610656738,
9.18278503417969,-10.0020933151245,
-45.5025329589844,11.0847721099854,
-57.2980613708496,2.41711950302124,
-20.0739917755127,-20.3250522613525,
3.70388269424438,-19.8359737396240,
-20.9401512145996,4.62908601760864,
-51.4587974548340,10.1759204864502,
-34.1556053161621,-20.6287231445313,
12.1529111862183,-42.9233322143555,
32.9202003479004,-11.0033397674561,
16.7701778411865,45.9338722229004,
3.09585809707642,56.1283454895020,
10.7191944122314,4.49496412277222,
15.1598358154297,-42.3786125183106,
-2.23472166061401,-21.9153728485107,
-16.7874774932861,37.4046936035156,
-10.0882387161255,63.5689353942871,
2.16539573669434,37.8731040954590,
-3.69069337844849,11.6831436157227,
-18.5086669921875,24.8413009643555,
-14.0317726135254,52.6220932006836,
13.6617355346680,52.3419914245606,
29.3884620666504,29.8892498016357,
13.1628656387329,20.1581192016602,
-15.2394018173218,32.4335975646973,
-24.5459003448486,38.2651519775391,
-11.8734741210938,25.3926143646240,
8.86659526824951,12.3320350646973,
19.0354671478272,19.1130771636963,
7.77907609939575,38.0290870666504,
-16.1280956268311,47.3849792480469,
-27.1462516784668,43.8408737182617,
-13.6193857192993,39.6143035888672,
5.33230590820313,30.9269580841064,
0.518926799297333,14.3606491088867,
-28.1900005340576,9.01370906829834,
-43.1662330627441,21.5082111358643,
-23.5940170288086,30.8206634521484,
2.81375098228455,9.33357715606690,
0.258671969175339,-32.0060882568359,
-13.3777112960815,-59.8660163879395,
5.04746294021606,-58.6990509033203,
44.8504829406738,-55.8352203369141,
51.7523269653320,-64.0891418457031,
10.2586097717285,-56.9194679260254,
-23.8203773498535,-22.6306018829346,
-4.74092817306519,-4.07201528549194,
36.2787132263184,-34.2601699829102,
35.4523468017578,-67.3526611328125,
-7.93581962585449,-36.6540679931641,
-38.4254875183106,40.1338195800781,
-28.8669013977051,74.6598358154297,
-15.2858381271362,34.7040824890137,
-26.8372230529785,-10.5406684875488,
-38.7351455688477,7.14776229858398,
-21.4439620971680,47.1330146789551,
3.23470258712769,31.4387969970703,
-0.295121252536774,-30.6770133972168,
-23.3678951263428,-51.7328109741211,
-30.2104358673096,-5.39204692840576,
-19.7304801940918,38.1276626586914,
-20.1037788391113,26.7458457946777,
-38.7315444946289,-3.93619966506958,
-45.5718879699707,-3.00554180145264,
-24.4501285552979,7.84104871749878,
-2.97604656219482,-14.9883842468262,
-10.5751190185547,-53.2258949279785,
-26.6658878326416,-45.4505157470703,
-16.2490367889404,14.9680404663086,
13.7003822326660,63.4646606445313,
28.3562030792236,53.9744377136231,
13.7126893997192,20.7923030853272,
-11.5772790908813,6.54585170745850,
-27.7335453033447,-0.956947028636932,
-29.5331153869629,-28.1869907379150,
-13.7195930480957,-56.2680587768555,
21.1310806274414,-53.6409187316895,
58.5874633789063,-33.2856369018555,
68.2220993041992,-26.7410545349121,
42.9764251708984,-31.6793289184570,
14.8309364318848,-14.0420227050781,
13.1821317672730,31.0602512359619,
25.5367012023926,56.0448226928711,
20.7216835021973,35.2673339843750,
-1.09838879108429,5.58005619049072,
-8.89089584350586,8.30856323242188,
8.89439964294434,24.6405372619629,
32.7457237243652,16.1393394470215,
41.1139183044434,-11.1010103225708,
34.3820610046387,-20.5229949951172,
26.3128395080566,-4.07860898971558,
21.8923072814941,5.88311195373535,
13.7947425842285,0.778881072998047,
1.59703922271729,8.86181354522705,
-11.1884765625000,38.9304656982422,
-19.5412082672119,51.7522048950195,
-17.3034877777100,9.03069972991943,
-2.76773071289063,-52.7436141967773,
17.5558719635010,-63.2202339172363,
19.2543449401855,-10.9312362670898,
-6.28362846374512,37.5301170349121,
-31.4144363403320,26.9154949188232,
-27.9414749145508,-26.9510803222656,
-1.56872534751892,-61.6940574645996,
12.8448238372803,-41.6690292358398,
-4.30062675476074,15.3845281600952,
-33.5056991577148,58.7437400817871,
-44.7591629028320,51.3226432800293,
-36.9792747497559,-1.53076457977295,
-25.6883335113525,-58.4391975402832,
-16.2060661315918,-68.4353637695313,
-1.80507409572601,-22.9991683959961,
7.69917011260986,28.1698589324951,
-4.83510208129883,35.0069923400879,
-31.5349674224854,3.78100824356079,
-35.7238655090332,-13.3945083618164,
1.43723154067993,1.32071614265442,
48.0859832763672,16.1554965972900,
55.6248588562012,10.4141311645508,
19.8828582763672,3.91872787475586,
-19.4986057281494,20.9071350097656,
-28.3326320648193,41.3297233581543,
-15.0076026916504,20.8643589019775,
-6.06547546386719,-31.4739761352539,
-5.02584886550903,-60.6346054077148,
4.68245029449463,-40.7124328613281,
21.7389202117920,-2.68717455863953,
28.4647541046143,7.30156135559082,
14.0705471038818,-9.25399875640869,
-7.94595050811768,-23.6400756835938,
-20.1194610595703,-29.8799934387207,
-17.3912754058838,-36.0489311218262,
-12.8044815063477,-36.4762039184570,
-13.7419881820679,-16.2953624725342,
-20.0288028717041,12.2535228729248,
-21.7950916290283,17.3905868530273,
-12.8724536895752,-11.1776142120361,
4.29259634017944,-41.0532989501953,
13.0327825546265,-41.8835411071777,
0.280276775360107,-17.7188854217529,
-19.1654453277588,10.6062564849854,
-21.3079814910889,39.0604286193848,
-2.72964859008789,64.6512832641602,
4.70422840118408,64.2750473022461,
-21.7354221343994,22.9393844604492,
-55.3742370605469,-31.8216228485107,
-47.6874008178711,-48.9440193176270,
13.4861602783203,-12.5916938781738,
74.4499588012695,36.0286712646484,
79.7038116455078,52.3164138793945,
38.8970489501953,38.9119834899902,
4.27292776107788,28.1075706481934,
5.60070896148682,32.6184577941895,
18.0429306030273,32.7609672546387,
8.58919334411621,17.6274452209473,
-22.8592243194580,2.56882762908936,
-47.1626167297363,3.56668376922607,
-49.9065551757813,16.5628299713135,
-37.4794464111328,25.5684757232666,
-16.4483127593994,25.8572101593018,
8.91740894317627,24.3090591430664,
22.3847045898438,26.0054779052734,
3.70545530319214,29.3367481231689,
-37.4408950805664,21.3601455688477,
-57.8524475097656,-2.62117147445679,
-28.6466178894043,-29.2099323272705,
18.7742614746094,-41.7709045410156,
37.2154960632324,-27.8704051971436,
25.7190227508545,0.345603942871094,
19.0680313110352,13.3518781661987,
39.5248107910156,6.12847328186035,
58.6216430664063,1.86057245731354,
46.0135574340820,14.8047409057617,
13.3005151748657,19.7781009674072,
-4.71930265426636,-9.16454029083252,
-2.93277549743652,-46.7791481018066,
6.17905139923096,-44.2026367187500,
13.9746246337891,3.01490736007690,
20.1599693298340,36.1868515014648,
17.3810291290283,12.2102737426758,
2.55011439323425,-29.0903797149658,
-1.43737435340881,-21.4686126708984,
23.9119834899902,28.9589347839355,
52.6227188110352,52.2797164916992,
37.6842880249023,21.2030906677246,
-22.2949237823486,-17.7000885009766,
-66.1238327026367,-15.7945728302002,
-47.0946846008301,4.55279588699341,
-5.37767076492310,0.864048480987549,
-4.38947486877441,-13.0703630447388,
-39.0055351257324,5.31226158142090,
-52.0129547119141,48.1760482788086,
-22.5986099243164,54.2480316162109,
10.1109962463379,-1.35667657852173,
14.5568494796753,-64.2405624389648,
11.4572029113770,-71.4674835205078,
27.3028945922852,-34.4319419860840,
45.6985168457031,-3.01693248748779,
36.1426734924316,8.90638923645020,
10.0475053787231,24.2749595642090,
2.17170429229736,47.5408325195313,
9.64362239837647,54.2120399475098,
-2.04805922508240,37.6954460144043,
-36.3415565490723,13.7212200164795,
-52.8514175415039,-1.49453377723694,
-29.2843284606934,-15.6942386627197,
-0.120999336242676,-32.8582839965820,
0.489089488983154,-30.1040668487549,
-14.2465066909790,1.64071977138519,
-14.1704120635986,28.5383358001709,
-3.16594886779785,11.2539005279541,
-10.1941261291504,-32.7914047241211,
-36.7835464477539,-54.7310180664063,
-47.7261276245117,-35.6179389953613,
-22.9683914184570,1.47752964496613,
9.72280979156494,23.8470191955566,
16.5771427154541,24.4477024078369,
6.56419563293457,6.94987964630127,
7.79815149307251,-29.1203536987305,
27.8337230682373,-68.0197830200195,
43.0710906982422,-72.3741302490234,
34.9649238586426,-25.8027210235596,
9.10072326660156,31.2756519317627,
-12.0417652130127,42.6664505004883,
-9.92157268524170,12.2147178649902,
13.9178180694580,-6.64602088928223,
36.8787612915039,14.5933666229248,
33.3967781066895,42.5774917602539,
-0.513211727142334,35.6630477905273,
-40.2179412841797,2.97061848640442,
-50.4836540222168,-14.4482059478760,
-23.1927394866943,-1.66410350799561,
12.5250110626221,16.3493747711182,
28.0442047119141,18.5539722442627,
19.2306175231934,18.3340492248535,
-2.18890023231506,29.8026714324951,
-23.7683544158936,43.9939575195313,
-34.4202575683594,45.8081283569336,
-29.3577251434326,42.0897369384766,
-19.2171821594238,44.8116531372070,
-18.2499675750732,46.5139579772949,
-29.9106979370117,35.8334999084473,
-30.2345199584961,14.4658060073853,
2.87455058097839,-6.46628904342651,
45.9027862548828,-16.0445022583008,
52.3301467895508,-11.3036489486694,
15.8175945281982,9.12693595886231,
-15.9870367050171,44.0512123107910,
-3.45900511741638,65.1580810546875,
22.7643089294434,46.0623779296875,
12.7013883590698,8.43911361694336,
-30.3926982879639,0.673461019992828,
-50.6380195617676,24.4926109313965,
-24.2285842895508,25.9786376953125,
2.54151368141174,-21.6905269622803,
-16.9567279815674,-64.8137893676758,
-52.8502922058106,-41.2011337280273,
-45.6286735534668,21.2718505859375,
7.78200244903564,33.7884674072266,
41.6825790405273,-20.9547023773193,
18.6771335601807,-62.9214134216309,
-26.4774589538574,-21.8299694061279,
-40.6103515625000,53.9249801635742,
-26.8841781616211,69.9971389770508,
-22.2590446472168,16.6900215148926,
-38.9185447692871,-28.9837303161621,
-50.5332832336426,-18.6779174804688,
-37.5125007629395,7.76431512832642,
-11.0265817642212,-3.17528486251831,
7.79238224029541,-45.6782722473145,
17.8700141906738,-64.8466644287109,
28.7596817016602,-35.8683509826660,
36.0333061218262,15.0584983825684,
38.3749961853027,42.9943847656250,
39.8604354858398,26.1473922729492,
41.3553886413574,-18.4685726165772,
33.8093681335449,-59.0732917785645,
16.0079421997070,-60.2253990173340,
3.41845703125000,-19.0950164794922,
4.15647983551025,17.1733646392822,
10.7691297531128,10.0406370162964,
9.12471008300781,-24.0714244842529,
7.24869775772095,-36.4983444213867,
20.9884510040283,-4.87377262115479,
37.4501609802246,40.9395751953125,
19.4673290252686,61.7716636657715,
-28.7698364257813,52.8938407897949,
-57.0233192443848,34.1252899169922,
-29.1876773834229,16.2530975341797,
24.7519092559814,0.940726935863495,
44.0562782287598,6.43645858764648,
16.8580589294434,43.3397789001465,
-19.9245052337647,79.4157562255859,
-34.4960289001465,67.7205429077148,
-41.6428260803223,3.81833600997925,
-52.9100418090820,-53.5172615051270,
-47.7923202514648,-55.6060523986816,
-7.23898315429688,-18.0689163208008,
34.4818534851074,12.7521448135376,
26.8726215362549,17.2122192382813,
-21.9078464508057,13.1881179809570,
-53.0085105895996,17.3363037109375,
-34.9119415283203,19.1359615325928,
1.75784993171692,7.69828510284424,
16.3265151977539,-6.08742380142212,
8.86559104919434,-15.0097265243530,
0.433913201093674,-22.6183242797852,
-7.90774250030518,-31.5090560913086,
-29.1983814239502,-34.6968612670898,
-50.1602668762207,-33.4193382263184,
-44.3201675415039,-41.5714721679688,
-20.7925510406494,-61.8440971374512,
-14.5557794570923,-64.0238113403320,
-26.3369140625000,-32.6221427917481,
-22.7951221466064,9.38766098022461,
4.50090694427490,18.2555751800537,
18.0480194091797,-8.70233345031738,
-6.51108360290527,-29.9849662780762,
-38.0156631469727,-17.6570625305176,
-28.0405216217041,8.64272403717041,
16.4947853088379,10.6857614517212,
39.7426795959473,-9.54329967498779,
24.4756660461426,-25.4627342224121,
7.82255792617798,-19.7121543884277,
17.0360317230225,-3.00937461853027,
28.9793853759766,5.64321708679199,
19.2631072998047,0.745951831340790,
4.86455345153809,-16.7339248657227,
11.6942787170410,-36.2512550354004,
23.4637355804443,-45.4402046203613,
8.88304710388184,-39.2271308898926,
-19.7831897735596,-28.0673637390137,
-17.8931217193604,-20.1531753540039,
21.8728237152100,-14.1050443649292,
48.3613777160645,5.09394168853760,
22.4995594024658,41.4854888916016,
-27.8698253631592,73.6547317504883,
-50.1504325866699,81.8541183471680,
-39.3250923156738,62.4143524169922,
-28.6694335937500,24.6496582031250,
-26.1545352935791,-11.7950077056885,
-14.0115709304810,-24.2333106994629,
11.1526107788086,-3.48619079589844,
22.1589851379395,26.3276195526123,
1.95958042144775,27.1319007873535,
-27.0054969787598,-8.92257976531982,
-35.2378425598145,-38.3940582275391,
-27.0687942504883,-20.7583141326904,
-26.3531723022461,26.9624233245850,
-35.9325828552246,45.1995201110840,
-34.3537292480469,7.50577831268311,
-16.5980834960938,-43.3916473388672,
1.55065870285034,-53.6533241271973,
13.2290172576904,-21.8932666778564,
27.2064800262451,12.5829858779907,
41.5807456970215,28.0847301483154,
38.6992034912109,31.3492641448975,
7.53379726409912,36.0258598327637,
-29.8814640045166,30.6118736267090,
-43.7722129821777,3.89484024047852,
-25.3874492645264,-26.1390724182129,
5.74184560775757,-37.5128211975098,
24.3206653594971,-35.1241683959961,
24.8211917877197,-42.0270957946777,
9.84432029724121,-55.4736022949219,
-11.6877346038818,-45.8949317932129,
-23.7694950103760,-5.93307924270630,
-21.1827430725098,24.6654720306397,
-16.8120384216309,7.93343305587769,
-21.7480621337891,-31.1505432128906,
-21.8128757476807,-35.6483421325684,
-6.19075870513916,6.43090057373047,
9.42843723297119,37.3210220336914,
-3.53004074096680,16.8087062835693,
-30.5738277435303,-25.0634765625000,
-28.1599559783936,-42.2965126037598,
18.7864017486572,-39.2868652343750,
58.2639274597168,-47.4585647583008,
36.9112167358398,-57.2349662780762,
-17.3058986663818,-32.4230308532715,
-36.0984344482422,17.8231601715088,
-8.57677555084229,31.1114196777344,
9.69363307952881,-13.3420410156250,
-9.95528411865234,-49.9618568420410,
-26.5184116363525,-23.6583652496338,
2.44621515274048,27.9347648620605,
49.0602416992188,25.0571517944336,
57.7763023376465,-32.7936096191406,
33.6224250793457,-66.7219161987305,
29.2293014526367,-38.4600334167481,
59.6786117553711,-1.36419951915741,
74.6529388427734,-5.93761110305786,
36.5742912292481,-29.4419479370117,
-21.9152088165283,-23.5796375274658,
-47.8986129760742,5.99155282974243,
-40.7243881225586,4.13567829132080,
-30.9949169158936,-41.8457183837891,
-19.1439666748047,-80.1003417968750,
9.01583957672119,-62.3424835205078,
43.3365020751953,-6.70557641983032,
48.9950065612793,33.5429725646973,
19.4987926483154,30.4036617279053,
-11.7952308654785,1.26368045806885,
-18.7764568328857,-18.0623741149902,
-17.9988594055176,-1.89700484275818,
-25.2979412078857,41.0482940673828,
-21.3007774353027,62.5602645874023,
6.16781473159790,31.7780055999756,
27.6452369689941,-26.9972305297852,
6.54880285263062,-54.9842643737793,
-27.9390029907227,-24.1940956115723,
-19.4740829467773,28.3948020935059,
33.7061119079590,43.9379615783691,
68.3164749145508,15.6178016662598,
41.2381401062012,-13.3401374816895,
-11.9609031677246,-12.4060764312744,
-30.2759647369385,6.65989685058594,
-16.5977630615234,26.7944946289063,
-17.0518836975098,35.8052253723145,
-45.7786483764648,21.9011230468750,
-61.0207595825195,-16.5812187194824,
-39.1038208007813,-55.6045989990234,
-0.339952588081360,-51.1207466125488,
24.2044830322266,5.41731643676758,
33.4060554504395,56.8578453063965,
34.8582038879395,46.9656181335449,
26.0395374298096,-8.57926177978516,
9.69315147399902,-38.5151557922363,
9.50131702423096,-10.7764015197754,
36.2586326599121,27.2225685119629,
61.1742439270020,28.7047328948975,
43.0503997802734,12.6447057723999,
-12.9784593582153,20.2616024017334,
-53.2412033081055,40.3448143005371,
-49.3408203125000,25.1925907135010,
-31.8783111572266,-29.5896625518799,
-34.0605964660645,-65.2739028930664,
-51.9880447387695,-38.4354705810547,
-54.8005332946777,15.5188264846802,
-37.1506958007813,35.3770370483398,
-18.2933921813965,15.6474313735962,
-14.1779651641846,-0.196696743369102,
-22.6668186187744,9.24214172363281,
-33.5538864135742,13.5586652755737,
-38.5331001281738,-6.78905677795410,
-29.3929500579834,-30.4653224945068,
-7.95274734497070,-33.6601676940918,
5.78636884689331,-23.1752490997314,
-7.61773967742920,-20.3897571563721,
-37.7892723083496,-27.6841297149658,
-44.6709251403809,-27.6712150573730,
-9.09693336486816,-17.4744834899902,
39.6081390380859,-12.7228279113770,
65.4801330566406,-13.5168781280518,
56.0049629211426,-2.38776326179504,
30.2257289886475,25.0501575469971,
4.74825668334961,47.3643531799316,
-15.3181009292603,52.8538398742676,
-31.7860984802246,45.3079414367676,
-41.7047843933106,28.2617454528809,
-42.7735366821289,1.90152132511139,
-35.5154304504395,-24.4065132141113,
-21.9165229797363,-23.6527729034424,
-9.04203128814697,9.22068023681641,
-5.14288377761841,32.4241867065430,
-9.16100788116455,4.68660116195679,
-7.20847368240356,-49.5689735412598,
13.5614433288574,-63.0240936279297,
45.2056121826172,-16.2885208129883,
60.4680976867676,33.4489784240723,
50.3539962768555,33.9130210876465,
28.4464054107666,6.23750543594360,
9.64151573181152,6.43913984298706,
-0.576114773750305,34.7678222656250,
-1.83334445953369,34.5620422363281,
8.20817756652832,-17.3311386108398,
19.4722690582275,-68.6670837402344,
19.3962841033936,-63.5577621459961,
11.3625030517578,-11.4766750335693,
15.2506446838379,29.5450344085693,
33.2737083435059,34.7507934570313,
38.4476852416992,26.4206161499023,
4.18238162994385,21.3239994049072,
-44.3924980163574,5.27337169647217,
-60.2657394409180,-26.5464458465576,
-36.1434440612793,-46.0068817138672,
-8.89211940765381,-29.4705715179443,
-0.811386644840241,5.35445499420166,
5.43528747558594,16.6636810302734,
22.1508159637451,-5.34185123443604,
27.7484130859375,-27.0117321014404,
2.73461818695068,-18.5805931091309,
-21.9229679107666,9.85120296478272,
-6.20427179336548,33.1676139831543,
35.1602249145508,44.0754890441895,
39.4606399536133,42.1465034484863,
-17.7603569030762,32.2615165710449,
-76.4431686401367,17.2295913696289,
-73.0875015258789,5.19095420837402,
-18.0774097442627,5.27974033355713,
16.8843154907227,15.0716762542725,
-3.11429858207703,25.2999248504639,
-41.6921615600586,29.8240966796875,
-46.4480895996094,26.3024959564209,
-10.1729068756104,19.1004676818848,
26.4963455200195,11.9588298797607,
31.4061355590820,18.2057170867920,
6.49412822723389,39.0945167541504,
-28.6196002960205,48.8942413330078,
-51.8436813354492,26.0870018005371,
-48.4264030456543,-16.4497146606445,
-14.2814340591431,-41.9949188232422,
35.8331146240234,-33.8240051269531,
67.5745849609375,-16.2951717376709,
62.2660903930664,-9.04752826690674,
37.9809951782227,-10.9873018264771,
26.3433265686035,-11.2405872344971,
34.1164436340332,-17.3639755249023,
34.2087097167969,-38.0259552001953,
15.5533828735352,-52.5388526916504,
5.51895570755005,-31.0300159454346,
22.7487144470215,14.7152137756348,
37.7427711486816,38.3349876403809,
13.8376598358154,14.0423088073730,
-36.1098670959473,-28.4209499359131,
-51.1569442749023,-50.3260841369629,
-8.70528602600098,-44.6475219726563,
37.9710655212402,-22.7154731750488,
35.4128608703613,12.1004371643066,
6.45018148422241,52.1566123962402,
2.04225063323975,73.5883712768555,
23.5117855072022,53.7361145019531,
21.9221153259277,9.28875446319580,
-6.68059301376343,-19.7899551391602,
-13.7572546005249,-17.9166736602783,
23.8186302185059,-8.50709533691406,
50.9934005737305,-1.46027266979218,
19.2598037719727,15.0612325668335,
-34.4029502868652,42.0690040588379,
-34.4864692687988,49.7082977294922,
21.7721347808838,22.4623966217041,
58.3576202392578,-4.38894891738892,
30.6461162567139,6.35020351409912,
-13.4951124191284,36.1052780151367,
-15.0500926971436,34.3052482604981,
16.0865726470947,-8.22551345825195,
32.1383247375488,-41.5264892578125,
19.8404521942139,-29.0703182220459,
10.2806510925293,-0.143974900245667,
22.6678047180176,-7.77990150451660,
41.1508598327637,-50.8091125488281,
40.2172546386719,-75.9606094360352,
20.2909622192383,-48.0222892761231,
-6.72638893127441,10.9296407699585,
-27.9020347595215,50.6578445434570,
-31.7352447509766,46.8306579589844,
-8.79715156555176,16.0774345397949,
18.6046676635742,-5.75523138046265,
11.3825340270996,0.303249835968018,
-32.9156951904297,16.5958728790283,
-63.9721679687500,16.4334030151367,
-41.3812294006348,-8.34234333038330,
15.4426469802856,-38.0587577819824,
49.3502502441406,-46.6152610778809,
39.0699462890625,-35.4807624816895,
19.4822483062744,-25.1884021759033,
25.9474086761475,-24.0638141632080,
47.6954421997070,-16.2494621276855,
53.0622940063477,4.46917533874512,
39.8850822448731,11.7067108154297,
30.5799922943115,-9.85639953613281,
35.0273895263672,-39.3905754089356,
40.2788238525391,-41.1408195495606,
33.9877014160156,-13.5940246582031,
22.3580055236816,-1.46212542057037,
12.0578155517578,-28.4446964263916,
2.69902372360230,-58.1415481567383,
-7.08674573898315,-37.7283935546875,
-13.7994804382324,22.3159179687500,
-14.0603237152100,64.2521514892578,
-5.59207439422607,56.9585189819336,
5.77813053131104,28.5932807922363,
11.9870290756226,11.0207233428955,
9.22712516784668,-4.84291267395020,
-3.77237844467163,-35.1337280273438,
-20.5812511444092,-50.9247360229492,
-24.1611270904541,-16.5428428649902,
-15.6454448699951,41.0525283813477,
-9.67184352874756,54.8923530578613,
-16.6629276275635,14.3344297409058,
-28.3113040924072,-13.3526802062988,
-37.0023002624512,18.1458873748779,
-42.3861007690430,56.9253768920898,
-43.0827865600586,33.5579299926758,
-27.2432384490967,-33.7011032104492,
6.19285774230957,-62.6845550537109,
27.3395214080811,-29.1127090454102,
7.37834167480469,4.22270441055298,
-34.2655639648438,-14.7068538665771,
-42.0852050781250,-53.3875808715820,
3.76677727699280,-51.9269294738770,
56.7909317016602,-13.8942146301270,
58.8213958740234,12.7816715240479,
14.8544645309448,11.8060789108276,
-16.6562728881836,9.68159580230713,
-8.33996486663818,14.4423074722290,
13.4688806533813,2.37936186790466,
9.12526226043701,-26.9731349945068,
-18.7215347290039,-36.3460006713867,
-34.4657402038574,-8.41742897033691,
-16.9401264190674,24.4579391479492,
16.4188232421875,21.7342910766602,
32.8630790710449,-8.52207183837891,
18.0966358184814,-17.5839195251465,
-9.80890560150147,10.1807565689087,
-20.2980365753174,38.2936668395996,
-0.422160208225250,34.3511886596680,
27.0525245666504,10.4672231674194,
28.1010532379150,-3.62292695045471,
-10.3310050964355,1.05531513690948,
-53.7383346557617,13.5258111953735,
-67.1079940795898,13.6458349227905,
-44.1217880249023,-6.01119804382324,
-6.99789381027222,-41.6463317871094,
22.7348270416260,-69.7769622802734,
40.2952995300293,-63.2423133850098,
43.3205261230469,-18.9131793975830,
28.5907478332520,30.5274658203125,
-1.84875595569611,43.1747398376465,
-24.2352313995361,15.6599617004395,
-19.6597290039063,-16.7781505584717,
6.65713214874268,-29.9088420867920,
31.1981372833252,-31.3118610382080,
40.4613304138184,-33.9555511474609,
41.9444503784180,-29.3829650878906,
45.4935188293457,-4.02519893646240,
48.4097137451172,33.0103683471680,
42.7903213500977,56.3959503173828,
27.6002101898193,53.9061660766602,
4.80350494384766,37.9547386169434,
-18.2885761260986,24.1869640350342,
-38.8224716186523,10.2261314392090,
-53.2536888122559,-2.79868221282959,
-60.9089088439941,-7.84637498855591,
-62.8334388732910,3.79564213752747,
-53.8241310119629,18.3825778961182,
-27.5396976470947,19.0739517211914,
9.91525840759277,6.37465286254883,
33.9060020446777,-6.05270242691040,
24.8865776062012,-8.49098968505859,
-5.27120828628540,-2.46553754806519,
-23.1968727111816,9.57599258422852,
-16.0430221557617,28.2054710388184,
-0.716573059558868,39.6274337768555,
-1.37010467052460,25.4762115478516,
-15.5995607376099,-17.8713512420654,
-20.5548725128174,-57.6600112915039,
-13.1002674102783,-64.2129898071289,
-10.0482807159424,-40.1224441528320,
-19.0371570587158,-20.5855751037598,
-29.1426277160645,-24.5285491943359,
-22.4076042175293,-38.6139945983887,
-7.10388946533203,-40.9925956726074,
-3.62150979042053,-29.4970378875732,
-18.2698574066162,-18.9556293487549,
-30.9932556152344,-19.8127994537354,
-23.2760353088379,-24.9512348175049,
-11.5508737564087,-20.0107917785645,
-17.4031295776367,-0.667646646499634,
-29.3845367431641,23.5957584381104,
-13.3131895065308,39.2990112304688,
35.1716766357422,40.7345771789551,
69.4633636474609,35.6415138244629,
46.3178176879883,37.2226715087891,
-12.8655347824097,44.2769508361816,
-48.2009048461914,40.2661476135254,
-34.7126235961914,19.7975635528564,
-6.54950141906738,-1.84557187557220,
10.8182411193848,-4.97646713256836,
28.8287868499756,5.87965393066406,
52.2130737304688,17.8862724304199,
46.1077880859375,24.8804435729980,
-6.77021408081055,32.5732231140137,
-57.3701896667481,34.0954780578613,
-44.1334915161133,18.4880027770996,
15.6422348022461,-10.0723619461060,
42.9474525451660,-21.1180324554443,
8.01496601104736,-2.28950381278992,
-28.4444160461426,24.8663597106934,
-16.0162887573242,32.4967994689941,
9.02117443084717,25.9319629669189,
-11.9077501296997,26.0021152496338,
-57.9034385681152,25.8439197540283,
-60.1179046630859,3.31631231307983,
-13.4559202194214,-35.3972702026367,
17.9205398559570,-53.5749282836914,
-1.49729108810425,-33.7471656799316,
-25.5469951629639,-11.4288072586060,
-4.75410079956055,-25.6092300415039,
33.6514587402344,-59.2956085205078,
35.9425582885742,-60.3730239868164,
2.95841503143311,-16.8579540252686,
-14.4838581085205,28.4518146514893,
5.61986541748047,41.4209175109863,
24.8735160827637,36.9809455871582,
11.5748577117920,40.4245300292969,
-10.6041727066040,39.5795707702637,
-5.62770557403564,5.68604135513306,
17.5093574523926,-44.9336624145508,
24.3658485412598,-60.4049224853516,
3.09363770484924,-19.5819072723389,
-26.0418930053711,32.4981346130371,
-32.2249488830566,43.0245780944824,
-10.7656822204590,11.1892242431641,
14.9015779495239,-15.6220035552979,
27.0110683441162,-14.0764312744141,
29.5446491241455,5.29955387115479,
33.6529006958008,28.3355770111084,
40.5119323730469,50.1029586791992,
35.7850608825684,58.9099388122559,
9.07342910766602,41.7114601135254,
-19.3072624206543,-0.610207855701447,
-13.5208511352539,-36.2803497314453,
25.3875617980957,-42.1237144470215,
47.0193862915039,-32.9119567871094,
15.8396186828613,-30.6597156524658,
-36.5712738037109,-36.1093673706055,
-43.0629806518555,-36.4091529846191,
8.63919639587402,-38.8514976501465,
58.5602836608887,-54.2534675598145,
46.6652374267578,-61.0046348571777,
-7.36681079864502,-25.0447044372559,
-41.1308250427246,38.1145515441895,
-31.8188629150391,66.0196533203125,
-14.1949119567871,24.9367122650147,
-22.6915302276611,-35.0573730468750,
-39.1724090576172,-36.6663818359375,
-33.0672340393066,24.0601844787598,
-6.61739444732666,75.8569183349609,
8.45667266845703,60.6070785522461,
-1.99915122985840,2.21401786804199,
-19.2378616333008,-34.7338066101074,
-27.8253993988037,-24.2883682250977,
-31.6592006683350,10.5147552490234,
-39.9157524108887,27.5747394561768,
-49.6880722045898,9.51347541809082,
-47.0007019042969,-29.4182224273682,
-30.6174278259277,-58.1961059570313,
-10.0025253295898,-52.0913810729981,
15.1260957717896,-19.8263740539551,
37.9798202514648,5.27859401702881,
38.1199722290039,-0.741367936134338,
11.1362285614014,-29.8767700195313,
-20.2844333648682,-49.5390777587891,
-25.6289119720459,-41.7768783569336,
-4.46398258209229,-20.4828681945801,
17.6298122406006,0.485524654388428,
25.0517559051514,21.6075725555420,
33.3580436706543,38.7504920959473,
48.5469436645508,47.8498497009277,
41.1640090942383,44.4525489807129,
-2.99202156066895,34.6419868469238,
-36.2375259399414,24.0653629302979,
-9.82766723632813,11.0811529159546,
43.4742927551270,2.09678030014038,
46.8561859130859,9.28623008728027,
-12.2462739944458,26.0527172088623,
-55.4900512695313,24.0017204284668,
-24.5506095886230,-15.5238361358643,
30.9605102539063,-60.8311271667481,
29.8743705749512,-55.9742240905762,
-17.6411056518555,2.86786174774170,
-35.4977607727051,51.3656044006348,
-4.94720935821533,41.0935440063477,
9.12062549591065,-11.5504970550537,
-19.1755790710449,-51.4320831298828,
-29.3669319152832,-56.1962585449219,
17.0049438476563,-41.4594383239746,
63.9933319091797,-18.4262657165527,
41.7472763061523,10.9233655929565,
-18.9708805084229,34.6030120849609,
-32.7458457946777,26.9169006347656,
12.6770410537720,-3.51612472534180,
39.4084129333496,-12.9800815582275,
0.120503902435303,16.6789512634277,
-52.8282089233398,42.0195236206055,
-60.0284881591797,19.8923492431641,
-38.3435592651367,-28.8824882507324,
-28.1982822418213,-41.9003601074219,
-18.3399581909180,-5.14690923690796,
10.7146492004395,36.3283233642578,
31.8526897430420,43.9963722229004,
8.33434486389160,27.4972534179688,
-33.7077636718750,15.0745935440063,
-30.8056182861328,5.16207075119019,
17.4146041870117,-19.2974910736084,
38.6455383300781,-45.5042114257813,
0.0496931672096252,-45.6015663146973,
-38.8940582275391,-23.0135803222656,
-14.5965614318848,-12.4329547882080,
41.7672882080078,-32.1737937927246,
52.3399085998535,-57.5515060424805,
17.1573143005371,-57.9009819030762,
3.72043800354004,-32.0895729064941,
40.9171714782715,-2.07638359069824,
78.4105606079102,11.7872076034546,
61.3072547912598,7.75061655044556,
10.2216110229492,-3.51664519309998,
-16.9288063049316,-13.7692670822144,
-3.73708200454712,-14.3918914794922,
11.0389328002930,-3.63148784637451,
-5.14816093444824,1.76657629013062,
-36.8417854309082,-10.3923130035400,
-48.3035850524902,-33.7791061401367,
-28.2875556945801,-47.0165786743164,
8.11651229858398,-41.9407882690430,
42.4892005920410,-31.7979354858398,
56.3549385070801,-26.0468120574951,
47.8284454345703,-17.4105453491211,
32.0244750976563,-0.122198581695557,
19.5023593902588,15.5161800384521,
9.38525199890137,7.84687805175781,
-3.73497700691223,-19.7687892913818,
-14.0112962722778,-43.0283050537109,
-15.2856111526489,-44.3044738769531,
-5.17368698120117,-34.4117736816406,
0.973667383193970,-32.4262619018555,
-2.45997667312622,-38.5752220153809,
-2.19814515113831,-39.2408828735352,
9.20723533630371,-28.0919437408447,
9.05658245086670,-11.9127807617188,
-18.2587223052979,-0.506801545619965,
-46.4268760681152,4.10295343399048,
-37.2972488403320,1.96560418605804,
2.65977001190186,-4.53880453109741,
22.7301731109619,-9.94774246215820,
1.74365901947021,-10.7031946182251,
-19.6298217773438,-12.2723388671875,
7.35777854919434,-25.3911705017090,
56.4770622253418,-39.8495368957520,
62.9440803527832,-29.8880195617676,
12.2513856887817,8.72461128234863,
-38.8865623474121,39.8046569824219,
-44.5359725952148,31.8220767974854,
-29.2319660186768,-3.89216804504395,
-35.5440635681152,-21.4077930450439,
-52.7452011108398,-2.92861700057983,
-44.3042030334473,21.5066013336182,
-11.9326210021973,21.9897766113281,
1.47802817821503,11.3197193145752,
-20.1893653869629,15.1917905807495,
-37.0425910949707,22.8667888641357,
-14.2582693099976,4.15402364730835,
31.9755706787109,-31.7469043731689,
59.3443374633789,-45.2650108337402,
53.1133041381836,-22.0189609527588,
31.4267654418945,1.98044300079346,
9.96708869934082,-8.53185558319092,
-6.75592565536499,-33.7504158020020,
-6.67030429840088,-36.1288337707520,
10.1272411346436,-15.9788970947266,
19.1922149658203,-7.73546886444092,
-3.23900508880615,-23.8401165008545,
-42.7886810302734,-37.4867820739746,
-55.5754585266113,-31.3351612091064,
-21.1342449188232,-22.9797420501709,
27.4702930450439,-25.7877349853516,
41.8611679077148,-15.6670341491699,
19.1926574707031,24.0146541595459,
-12.1513795852661,68.3665008544922,
-29.0025024414063,70.4926605224609,
-29.1801452636719,27.7085971832275,
-15.3157997131348,-17.0492706298828,
5.54670572280884,-29.1389198303223,
21.5497951507568,-20.6500797271729,
20.4549961090088,-16.2470798492432,
9.36252021789551,-12.1149110794067,
5.47661733627319,7.87911462783814,
7.07848453521729,35.0294647216797,
-8.17909812927246,45.1332473754883,
-45.8667831420898,30.2190799713135,
-73.7058334350586,4.37700939178467,
-55.6220626831055,-20.5845890045166,
6.75198364257813,-42.4514503479004,
62.3488006591797,-60.3928718566895,
71.1922683715820,-64.1382904052734,
40.8677978515625,-49.3071060180664,
7.13309192657471,-26.2210140228272,
-5.07131099700928,-9.45938396453857,
-0.978450000286102,3.08982610702515,
0.921221375465393,14.5960731506348,
-6.09249114990234,18.0192298889160,
-8.90009212493897,12.0720310211182,
2.09147882461548,8.93102741241455,
12.4575576782227,15.6441402435303,
2.56650424003601,18.0778350830078,
-23.7544021606445,1.57994377613068,
-35.3953399658203,-20.9308319091797,
-6.58818292617798,-21.3048915863037,
41.2866210937500,2.16923975944519,
60.4944801330566,13.0847396850586,
30.4891357421875,-5.21152114868164,
-7.90288305282593,-21.5935821533203,
-6.36056089401245,-2.08688759803772,
25.3193187713623,33.0848121643066,
37.2375907897949,34.6357192993164,
6.05089378356934,-1.03223633766174,
-30.2741909027100,-23.2365760803223,
-22.9893684387207,1.82795166969299,
15.3663549423218,37.2305297851563,
28.3498840332031,29.8788299560547,
-5.97904729843140,-16.7197227478027,
-48.9959106445313,-50.0074920654297,
-55.0646057128906,-40.9180946350098,
-26.9208850860596,-14.7523498535156,
-2.57180833816528,-10.9141530990601,
-0.108388289809227,-28.6309146881104,
-2.87009978294373,-38.4114074707031,
0.541018187999725,-33.3736038208008,
-0.775013208389282,-30.6468009948730,
-11.0855789184570,-41.3516654968262,
-12.6260633468628,-48.2274360656738,
10.8406276702881,-28.2611923217773,
43.9004058837891,15.9790248870850,
49.0664634704590,47.6685180664063,
17.0941944122314,35.9979705810547,
-19.1512241363525,-3.29811716079712,
-26.0377807617188,-27.0325164794922,
-3.37841916084290,-10.6787528991699,
20.5719242095947,24.0088138580322,
23.3164272308350,36.4213409423828,
8.39768695831299,18.6618499755859,
-2.10334944725037,6.20047426223755,
2.26475095748901,28.0047473907471,
15.2972364425659,61.3567352294922,
22.5824127197266,63.0431327819824,
16.1813774108887,28.6241455078125,
6.85607290267944,0.303634703159332,
11.1718769073486,11.8645935058594,
30.4348011016846,41.1407356262207,
44.5990829467773,41.0925445556641,
31.3631095886230,0.647413492202759,
-0.388015985488892,-37.1440467834473,
-25.2804126739502,-42.5845947265625,
-25.7258701324463,-25.3049793243408,
-8.95392608642578,-8.16701412200928,
4.00882625579834,12.4877643585205,
1.66762804985046,45.8268814086914,
-13.1797304153442,68.4943161010742,
-36.4187812805176,44.0689315795898,
-58.2236862182617,-14.2901248931885,
-66.6897888183594,-52.7625198364258,
-56.4251403808594,-40.3553314208984,
-34.5657577514648,-11.0186576843262,
-15.8041467666626,-8.27411270141602,
-3.88287496566772,-24.3454761505127,
10.9601202011108,-16.3524551391602,
27.8548164367676,19.5076351165772,
34.3478889465332,46.9818496704102,
23.6236228942871,46.8289031982422,
3.23155641555786,35.7398262023926,
-8.14946365356445,28.3618640899658,
0.102022051811218,17.1238059997559,
22.1245727539063,2.78067421913147,
40.4382934570313,8.60088443756104,
38.4283294677734,40.6714210510254,
7.85186767578125,60.6082344055176,
-34.6334381103516,38.1754188537598,
-51.9916915893555,-3.20525312423706,
-27.5885047912598,-9.86311531066895,
10.2222833633423,18.1912117004395,
12.4210233688355,24.7040004730225,
-23.8004016876221,-9.72441291809082,
-49.8948287963867,-42.5791549682617,
-27.7107505798340,-29.8294410705566,
20.6069030761719,10.4975843429565,
40.1875457763672,35.3120002746582,
21.8599433898926,34.9194946289063,
7.54192066192627,28.9620513916016,
24.5656719207764,22.7567577362061,
46.5955047607422,6.81451034545898,
38.1730270385742,-8.37501716613770,
11.1407451629639,4.34602165222168,
2.04483079910278,40.3025856018066,
14.5550432205200,56.2885437011719,
17.8981952667236,29.5002632141113,
-2.57784056663513,-2.56570816040039,
-20.1307735443115,2.29205298423767,
-13.1303119659424,35.6801795959473,
-2.07374405860901,55.0763511657715,
-17.7075443267822,44.2237739562988,
-47.1885337829590,22.5150070190430,
-54.2964820861816,6.24372243881226,
-27.7243289947510,-5.52487993240356,
0.383987367153168,-18.3066024780273,
10.8608617782593,-21.2669982910156,
11.4631710052490,-10.6630802154541,
9.23924541473389,-1.06583678722382,
-8.62568187713623,-8.92175197601318,
-41.7914619445801,-21.7790527343750,
-58.6137924194336,-18.4305515289307,
-33.4354133605957,-0.973302125930786,
8.35743331909180,12.7983388900757,
16.9231586456299,12.9200077056885,
-11.7546529769897,1.07433915138245,
-26.9141998291016,-13.0472488403320,
1.52254080772400,-17.7419109344482,
42.9911651611328,-1.78197145462036,
57.3653221130371,27.9968070983887,
48.6968193054199,46.5881729125977,
41.3936767578125,29.6696777343750,
37.7047080993652,-3.06758451461792,
23.1297473907471,-6.43125391006470,
0.100330591201782,29.4162197113037,
-10.5761423110962,55.1476058959961,
-10.0715093612671,27.5760459899902,
-17.5446357727051,-30.0623626708984,
-29.9059143066406,-60.1142234802246,
-21.1098003387451,-41.2088088989258,
12.6739940643311,-4.46401166915894,
27.9429378509522,18.9323940277100,
-0.312089979648590,33.7177352905273,
-39.3148155212402,48.1419067382813,
-42.9813270568848,45.5572967529297,
-19.7376289367676,9.74800300598145,
-15.2126607894897,-31.5761280059814,
-40.6322479248047,-38.1452178955078,
-57.0103492736816,-10.8691444396973,
-32.3496475219727,6.63805580139160,
9.79175662994385,-9.67385482788086,
26.5622158050537,-26.4774112701416,
14.4780635833740,-8.46576118469238,
1.20898652076721,32.8759422302246,
-2.71594762802124,54.5377807617188,
-11.5750617980957,34.9592208862305,
-30.0174674987793,-5.22186326980591,
-43.2844696044922,-31.6701374053955,
-37.2246475219727,-34.0525741577148,
-18.6580028533936,-20.8288955688477,
-1.74497568607330,2.05103731155396,
5.20879554748535,25.3359699249268,
0.137154683470726,39.6774597167969,
-9.06472873687744,42.4601936340332,
-10.9573659896851,38.7552871704102,
6.89670705795288,26.4977340698242,
37.9310607910156,-2.60423564910889,
51.6639976501465,-37.4137573242188,
29.9416198730469,-51.3371200561523,
-2.02372741699219,-32.4198226928711,
-4.63764286041260,-5.65904712677002,
25.3609485626221,0.104553729295731,
54.3899421691895,-7.33072090148926,
58.6052742004395,9.43785381317139,
40.6949043273926,49.4261817932129,
11.9004344940186,64.3788833618164,
-19.0092716217041,26.6157550811768,
-43.4575386047363,-28.1233520507813,
-40.8732948303223,-44.3987503051758,
-10.3692569732666,-20.3441810607910,
11.8706188201904,3.23035025596619,
-7.45379400253296,7.59479045867920,
-44.4284477233887,7.23643302917481,
-52.6603050231934,17.1919555664063,
-27.4635086059570,21.2954406738281,
-10.6918611526489,9.34025764465332,
-17.2816028594971,2.83702182769775,
-8.63274192810059,18.6621685028076,
32.2273902893066,32.8760833740234,
59.5150451660156,18.8000907897949,
25.4418029785156,-8.28540897369385,
-40.5809020996094,-13.6065959930420,
-57.1874809265137,-2.27082490921021,
-13.4460287094116,-4.91276788711548,
19.5283374786377,-20.4922370910645,
-6.22632503509522,-23.2199497222900,
-43.4841041564941,-10.0587329864502,
-26.8606719970703,-15.4958553314209,
29.1899242401123,-50.5880889892578,
62.2099227905273,-67.0145492553711,
51.9983978271484,-24.9775943756104,
29.4848880767822,30.6509571075439,
13.5907592773438,29.1781482696533,
-5.70180416107178,-20.3961677551270,
-28.9858531951904,-45.4981117248535,
-26.4911365509033,-24.7406501770020,
7.89238739013672,-12.6881599426270,
34.4532127380371,-41.3637924194336,
26.2339076995850,-61.3672294616699,
18.6508464813232,-21.9680118560791,
42.5415763854981,42.6473731994629,
64.8933639526367,59.8569297790527,
41.9961433410645,25.8109321594238,
-3.87511253356934,4.72653388977051,
-16.8286342620850,20.9730625152588,
3.14957618713379,24.9338645935059,
5.83309745788574,-8.95351314544678,
-24.2772674560547,-34.1415672302246,
-34.3713150024414,-8.62177753448486,
7.95164871215820,30.0602073669434,
44.9851150512695,25.0998973846436,
16.2993316650391,-13.4471006393433,
-38.2099571228027,-34.3766937255859,
-33.8237609863281,-23.9832019805908,
29.0068931579590,-13.1777324676514,
67.3622589111328,-13.7458057403564,
43.0701866149902,1.12775588035584,
7.11091899871826,35.5806655883789,
8.80083370208740,41.7459144592285,
19.4217453002930,1.51136255264282,
-5.48009729385376,-32.6803627014160,
-47.9771308898926,-14.1180171966553,
-51.9569702148438,26.0276012420654,
-16.2377662658691,30.1057834625244,
5.32701396942139,0.153148889541626,
-3.84706306457520,-18.7814464569092,
-4.93016147613525,-13.4879703521729,
23.8353404998779,-13.3433647155762,
42.8604087829590,-26.2152156829834,
25.1540985107422,-14.9419240951538,
-1.11109423637390,32.0124549865723,
-3.54439043998718,57.5506706237793,
6.24892377853394,19.5624446868897,
0.119740128517151,-40.7839736938477,
-15.5045471191406,-60.1302185058594,
-9.76934814453125,-43.0095138549805,
13.6602869033813,-38.8604087829590,
14.1771163940430,-51.6547622680664,
-18.0117568969727,-39.6935348510742,
-40.2620735168457,-3.32846665382385,
-24.0909500122070,5.11539363861084,
4.54719781875610,-35.2588539123535,
22.4783611297607,-64.2786178588867,
39.8925781250000,-26.6741485595703,
64.6781692504883,37.1503562927246,
71.7372207641602,42.6410255432129,
40.9043655395508,-10.9772605895996,
1.86634874343872,-39.9446868896484,
-4.47499322891235,-3.83500003814697,
9.09866905212402,41.7292900085449,
-7.92951679229736,35.4077415466309,
-51.7122230529785,-8.18518161773682,
-57.3112297058106,-39.0264816284180,
-3.30961298942566,-39.7078018188477,
42.1320838928223,-38.3043708801270,
17.4773063659668,-45.9303474426270,
-31.8464317321777,-43.8054504394531,
-26.1150188446045,-19.7193164825439,
26.6737632751465,10.7243194580078,
48.0453681945801,30.4127311706543,
5.93167257308960,39.7619781494141,
-35.2113571166992,31.7081451416016,
-17.9470577239990,-2.45001554489136,
20.9510383605957,-41.3134574890137,
19.0135612487793,-47.8135490417481,
-19.1781806945801,-23.8501186370850,
-32.7750282287598,-14.0090322494507,
-7.71388339996338,-39.1847381591797,
18.1114196777344,-63.8308563232422,
25.7476139068604,-44.0853347778320,
39.9202880859375,4.83704996109009,
62.5401687622070,28.4392280578613,
54.4945602416992,18.4743366241455,
1.03723931312561,16.6800785064697,
-54.5274276733398,38.6316223144531,
-59.1235885620117,38.9460906982422,
-18.7519950866699,-9.48617744445801,
13.3695440292358,-63.0318832397461,
10.8711156845093,-64.8379592895508,
-0.334788858890533,-20.2685432434082,
-5.45148372650147,13.8019046783447,
-15.9931716918945,15.9296646118164,
-32.8533363342285,9.75681400299072,
-37.2357406616211,12.9778184890747,
-25.9487133026123,6.55388736724854,
-17.5268001556397,-19.8360443115234,
-12.8401784896851,-32.6678276062012,
7.71549892425537,-6.75414085388184,
43.5056610107422,26.1663303375244,
53.5007553100586,20.7632026672363,
15.5757160186768,-9.49226665496826,
-28.7630233764648,-15.7255315780640,
-17.4272632598877,13.6070127487183,
34.0410537719727,37.0564575195313,
45.7321586608887,29.5666522979736,
-4.65843629837036,6.06128072738648,
-51.0061302185059,-11.1419191360474,
-39.9604301452637,-30.7465801239014,
-1.08769059181213,-63.1969566345215,
9.86709880828857,-78.2891082763672,
-3.60097646713257,-42.2846641540527,
3.98875761032105,23.1693439483643,
28.0275287628174,59.8821754455566,
20.9771366119385,50.7142486572266,
-21.1951522827148,27.5278339385986,
-36.3047866821289,15.7747707366943,
5.95229530334473,9.62180519104004,
53.0011367797852,5.07257175445557,
39.1967086791992,18.6294059753418,
-13.1314535140991,52.2210235595703,
-38.8145828247070,72.1891555786133,
-28.1506786346436,46.4405250549316,
-27.5083675384522,-6.15186786651611,
-47.8281631469727,-33.6448059082031,
-47.5946998596191,-24.4510517120361,
-1.61960470676422,-10.0694608688355,
49.8035812377930,-2.57718300819397,
55.4406433105469,15.1592426300049,
25.2619915008545,46.3204727172852,
9.53926086425781,56.7631645202637,
23.0572929382324,31.5081424713135,
37.7684020996094,-2.17948150634766,
38.2484397888184,-10.5924634933472,
37.8133087158203,-9.55885410308838,
41.8459663391113,-25.7611274719238,
40.9889945983887,-42.9063606262207,
34.0171966552734,-18.2063808441162,
31.7473430633545,34.2200965881348,
31.4214572906494,47.7814941406250,
19.1873035430908,-2.28289389610291,
-9.55801296234131,-48.2573165893555,
-32.6089019775391,-28.9725303649902,
-31.8334407806397,22.5550785064697,
-20.6555519104004,33.7638664245606,
-21.7956142425537,-1.79500079154968,
-24.4911651611328,-19.4045429229736,
-7.79321670532227,15.5497159957886,
13.1985769271851,61.0294837951660,
10.0387544631958,66.5798721313477,
-12.4042329788208,45.8651237487793,
-24.9189167022705,39.9202270507813,
-21.0283737182617,43.2086372375488,
-32.6267280578613,28.4995098114014,
-65.2351074218750,2.24796414375305,
-76.0924682617188,-5.33518457412720,
-29.4257698059082,7.07197618484497,
35.6671562194824,14.7861309051514,
52.8275413513184,13.7059192657471,
15.6083602905273,20.9069442749023,
-13.6118488311768,30.7821769714355,
5.49796962738037,17.2381191253662,
35.2852668762207,-15.1581926345825,
26.9028816223145,-16.7855319976807,
-10.9557847976685,32.2698860168457,
-27.2637634277344,69.9749603271484,
-3.59836244583130,30.5310211181641,
28.8192844390869,-48.1561431884766,
37.6804695129395,-68.0943450927734,
22.3723754882813,-9.05395698547363,
7.91648292541504,47.9450607299805,
7.51257419586182,35.3531417846680,
16.7619209289551,-17.6630496978760,
22.9799098968506,-39.1951637268066,
18.7387142181397,-22.2366886138916,
-2.89516949653626,-13.9326219558716,
-27.1311817169189,-33.8573837280273,
-28.9000949859619,-50.1643142700195,
-7.93173694610596,-40.1407127380371,
12.7967023849487,-21.2180709838867,
17.0858135223389,-10.8079271316528,
10.7516746520996,4.74151706695557,
4.12578201293945,32.9783706665039,
-8.47556591033936,42.3759880065918,
-34.2085762023926,8.81342887878418,
-51.9926986694336,-38.9538536071777,
-26.9867973327637,-52.9319458007813,
22.8336830139160,-14.5242528915405,
32.7107734680176,40.4325561523438,
-19.3351440429688,62.6097488403320,
-69.6668548583984,43.2792053222656,
-56.0876579284668,7.08853340148926,
-5.07900047302246,-16.9601173400879,
5.78000164031982,-13.6023225784302,
-35.8685989379883,7.99800968170166,
-54.4350204467773,19.4585838317871,
-7.12959957122803,4.54874992370606,
46.9859199523926,-8.95373725891113,
35.0643844604492,9.52074909210205,
-13.2076072692871,47.4957046508789,
-15.4157009124756,51.4971046447754,
30.1670589447022,5.11882209777832,
43.0283126831055,-38.4000358581543,
-7.74117851257324,-26.3113136291504,
-45.8266372680664,25.5228042602539,
-10.0008201599121,48.4429855346680,
48.7090682983398,23.7343311309814,
40.3354187011719,-0.260378092527390,
-28.6782932281494,12.9885730743408,
-69.3988037109375,35.5830421447754,
-37.3020629882813,23.2837944030762,
13.9431591033936,-10.3693809509277,
25.9223785400391,-17.8187580108643,
14.4171895980835,13.1972351074219,
21.6746616363525,46.8198852539063,
38.4220504760742,53.9443092346191,
31.8341941833496,41.4862632751465,
8.33950042724609,26.3435516357422,
-4.36513423919678,3.75838565826416,
-1.59711074829102,-29.0542316436768,
-8.04356384277344,-53.3726463317871,
-29.2270755767822,-53.5184135437012,
-42.8885955810547,-45.2374038696289,
-29.0231571197510,-44.9232330322266,
1.07402503490448,-36.5767936706543,
22.1722431182861,-0.812819480895996,
30.9038124084473,42.1679878234863,
29.0903854370117,51.5758514404297,
9.56593894958496,33.8429298400879,
-16.3754673004150,32.8896179199219,
-23.0731945037842,62.7997474670410,
-9.10782527923584,74.0839614868164,
-3.62491273880005,24.4421977996826,
-23.1257076263428,-42.7976341247559,
-46.1266555786133,-48.2869262695313,
-45.7747268676758,8.00847244262695,
-30.0024070739746,47.1746749877930,
-27.5327835083008,20.9744510650635,
-29.0806789398193,-29.0679855346680,
1.22635793685913,-43.8049240112305,
53.9401702880859,-20.8745079040527,
65.2972030639648,4.70737838745117,
14.3640441894531,22.5745716094971,
-36.7854881286621,44.7794876098633,
-22.5826435089111,57.6387062072754,
29.5522747039795,33.7723922729492,
34.2029418945313,-17.1850814819336,
-21.1268711090088,-38.6661643981934,
-58.4932022094727,-10.1593637466431,
-26.9577732086182,26.8441314697266,
26.2997055053711,31.7479515075684,
24.6716251373291,21.6933479309082,
-26.5910434722900,25.4494686126709,
-51.3478965759277,31.7272777557373,
-14.3475904464722,16.8568267822266,
31.1432800292969,-3.79548597335815,
23.7592220306397,5.99296617507935,
-27.0643577575684,41.7904586791992,
-61.0022430419922,53.7126197814941,
-44.3969535827637,31.1770381927490,
4.16348028182983,18.1448707580566,
37.8140792846680,39.9522056579590,
29.0878143310547,55.2425689697266,
-8.98801612854004,21.0000267028809,
-44.6527328491211,-26.7338314056397,
-57.3830680847168,-23.9854412078857,
-51.9739799499512,25.4465408325195,
-43.6816062927246,50.5783920288086,
-41.3793144226074,15.9508380889893,
-34.0276565551758,-29.7707481384277,
-18.7236022949219,-26.9717578887939,
-9.68205356597900,9.15444946289063,
-17.4544830322266,18.3045215606689,
-25.4562568664551,-16.9748401641846,
-12.4195966720581,-53.5863113403320,
13.0817766189575,-54.2261428833008,
25.7506999969482,-36.4362716674805,
10.4095239639282,-27.0741004943848,
-15.1461696624756,-21.4876613616943,
-27.7071781158447,3.04750251770020,
-25.9156684875488,38.2279624938965,
-19.2125396728516,51.1684150695801,
-8.27139472961426,20.3939170837402,
11.1331968307495,-27.4279956817627,
37.9007301330566,-44.8470916748047,
52.3086395263672,-19.1888904571533,
49.9171066284180,15.6382913589478,
37.9284667968750,25.2759952545166,
22.7112236022949,12.1218795776367,
-0.481098890304565,5.35103940963745,
-33.0428428649902,22.7570495605469,
-57.0386810302734,44.9218177795410,
-49.6289024353027,36.7952766418457,
-19.6963157653809,4.80874824523926,
4.20103549957275,-10.7774085998535,
5.15372610092163,11.8528909683228,
-3.57237672805786,45.4221725463867,
-11.8793478012085,48.1958694458008,
-32.4704284667969,20.4394855499268,
-67.6872711181641,-2.96754407882690,
-82.9776229858398,2.35809636116028,
-43.0697479248047,14.2622766494751,
26.0200901031494,8.93234157562256,
51.6753616333008,2.74789810180664,
7.30958986282349,18.4635944366455,
-53.0062141418457,39.0696907043457,
-54.3991088867188,22.5589351654053,
-1.36615943908691,-37.0302314758301,
42.0627250671387,-81.1479873657227,
42.3678054809570,-59.4715614318848,
22.9974765777588,4.09797573089600,
17.2701568603516,44.8557128906250,
20.3709163665772,38.2263908386231,
15.4177360534668,22.1177310943604,
5.26348066329956,33.9974975585938,
3.92014098167419,58.4438819885254,
7.46748065948486,49.6371192932129,
1.58946061134338,-0.134896039962769,
-10.6538448333740,-46.8662872314453,
-19.0165557861328,-51.1477203369141,
-25.8343753814697,-24.9223327636719,
-43.2341613769531,-11.4589824676514,
-60.4136772155762,-31.5222301483154,
-43.2323112487793,-58.8936042785645,
9.38048934936523,-52.3077964782715,
55.7141914367676,-7.87435388565064,
61.6667060852051,32.0125236511231,
40.4244689941406,34.4835929870606,
24.6175136566162,12.4269762039185,
24.5156612396240,-1.98093068599701,
22.2036819458008,0.843639969825745,
12.8717546463013,-0.886992394924164,
13.3644189834595,-20.0325584411621,
26.6649150848389,-33.5493583679199,
32.5441932678223,-17.2390327453613,
21.6129817962647,10.8889961242676,
13.0158748626709,17.7444171905518,
22.6991271972656,3.84071636199951,
28.5956039428711,0.268265902996063,
6.10276460647583,22.1784343719482,
-33.4561805725098,38.8805007934570,
-49.6526374816895,16.1430778503418,
-33.7485122680664,-31.3366432189941,
-16.1520690917969,-52.5300521850586,
-21.2069129943848,-32.6283493041992,
-36.1391410827637,-8.34683418273926,
-30.7653656005859,-18.0638542175293,
-6.08269405364990,-52.3459243774414,
11.9389429092407,-65.6971282958984,
10.0972681045532,-37.0161933898926,
-5.21985101699829,3.87171554565430,
-23.4791755676270,18.5198326110840,
-39.5951766967773,4.99341726303101,
-41.8186340332031,-15.5485448837280,
-20.0067863464355,-27.6489276885986,
16.9088630676270,-38.2555923461914,
41.6920089721680,-52.6356964111328,
36.7978477478027,-54.1984024047852,
11.6231231689453,-28.7375106811523,
-11.4862623214722,10.6593074798584,
-21.4685440063477,31.1349868774414,
-23.8171138763428,15.3650445938110,
-19.4553680419922,-14.8486461639404,
-7.91020011901856,-26.2218685150147,
6.76412630081177,-3.55113840103149,
13.4135503768921,30.5690536499023,
11.1364374160767,38.7843017578125,
7.12075233459473,5.49972867965698,
2.05932021141052,-45.4647216796875,
-7.83241462707520,-69.2714233398438,
-22.9486274719238,-40.7874794006348,
-27.5371665954590,16.2547931671143,
-13.7502117156982,49.2122268676758,
12.7556066513062,37.8323516845703,
31.6834220886230,12.1653013229370,
29.4981746673584,11.2876939773560,
15.6617889404297,34.4376106262207,
3.84661626815796,50.8916091918945,
3.96094679832459,42.5761108398438,
16.1332778930664,24.2330379486084,
28.0500659942627,19.1259212493897,
23.4566707611084,25.8022689819336,
-2.56583333015442,33.4635276794434,
-30.8668594360352,42.5398750305176,
-42.9711418151856,43.1791419982910,
-40.2383766174316,19.9020671844482,
-43.4356536865234,-23.9803524017334,
-57.0043983459473,-50.0844650268555,
-55.3788681030273,-24.4299736022949,
-21.3731231689453,21.0786380767822,
22.2094535827637,26.6961612701416,
32.5333366394043,-15.0840721130371,
5.22773742675781,-48.7448043823242,
-20.0375041961670,-32.5909271240234,
-14.5843830108643,-1.40992629528046,
3.65627264976501,-8.46598148345947,
4.50143098831177,-42.0841293334961,
-7.47242641448975,-38.3849220275879,
-1.31738448143005,14.8786926269531,
28.5909023284912,63.5142631530762,
51.4580764770508,62.2699584960938,
41.2538871765137,27.2760887145996,
7.02625989913940,-1.59580302238464,
-17.0450725555420,-15.7668619155884,
-19.5127182006836,-29.5102157592773,
-10.3626966476440,-35.0391616821289,
-5.10426616668701,-19.3376350402832,
-9.73605632781982,6.85039329528809,
-24.9260711669922,13.3973388671875,
-38.2552795410156,-1.74245333671570,
-31.9585914611816,-11.3614511489868,
-5.50514030456543,-4.50589418411255,
19.8602485656738,-10.2874622344971,
26.0264434814453,-34.9028625488281,
18.7123374938965,-47.1571159362793,
16.3637733459473,-23.8773155212402,
17.0409107208252,6.63710975646973,
-2.32982015609741,3.67675995826721,
-40.2272491455078,-33.6230659484863,
-56.5594291687012,-62.9900665283203,
-25.1430721282959,-59.9418067932129,
20.5131378173828,-41.7292480468750,
26.8217544555664,-28.7583255767822,
-8.31769752502441,-23.2806415557861,
-31.7957191467285,-24.6984539031982,
-6.80708599090576,-42.5169830322266,
44.1603469848633,-62.4659194946289,
73.3891143798828,-46.9817810058594,
66.6644210815430,12.1494035720825,
45.5900268554688,61.4806327819824,
24.3600463867188,52.7021789550781,
2.17713046073914,7.59609413146973,
-19.4048805236816,-9.72910308837891,
-28.2066612243652,19.3111171722412,
-25.6800956726074,45.2952308654785,
-26.6221427917480,25.5702018737793,
-28.8787975311279,-11.9960832595825,
-14.7341613769531,-22.3775424957275,
9.74163055419922,-9.97088050842285,
16.4128799438477,-4.99099254608154,
-4.85301542282105,-17.5055446624756,
-22.7211132049561,-28.3673267364502,
1.12693858146667,-34.8708686828613,
48.8831481933594,-43.9833526611328,
62.8057365417481,-44.8887977600098,
21.2161102294922,-12.9904727935791,
-32.8937911987305,31.5883045196533,
-58.1044921875000,35.9580688476563,
-47.0019416809082,-16.1535110473633,
-19.7519741058350,-65.2070541381836,
15.0425148010254,-44.0214881896973,
45.7832107543945,30.5394821166992,
45.1102333068848,76.9683380126953,
4.38422155380249,49.6820297241211,
-38.4513702392578,-11.1173229217529,
-28.9570980072022,-45.9959907531738,
27.6471519470215,-41.3917465209961,
67.4863204956055,-26.2159843444824,
44.9452056884766,-22.9248867034912,
-0.765351295471191,-27.3604068756104,
-4.02523803710938,-30.0719814300537,
38.9500999450684,-29.7499122619629,
73.1465606689453,-25.5234241485596,
60.4780540466309,-13.4846868515015,
13.1741333007813,12.5436744689941,
-26.6400470733643,37.5150451660156,
-38.0511665344238,40.8720817565918,
-25.4241619110107,17.4312381744385,
2.56844305992126,-15.3682003021240,
29.5237312316895,-33.2808723449707,
40.2449073791504,-20.7640647888184,
36.7099189758301,4.14206123352051,
40.5309715270996,13.2584676742554,
60.9879150390625,7.42495679855347,
69.5649871826172,11.9127521514893,
35.4999160766602,38.8583793640137,
-16.5805969238281,58.4241333007813,
-33.4380226135254,30.9009761810303,
-3.36813354492188,-31.6680660247803,
26.4140396118164,-61.9566879272461,
8.48610973358154,-20.9029579162598,
-42.8564682006836,47.5232009887695,
-68.3146743774414,63.1208648681641,
-42.8819503784180,19.0261554718018,
4.98949909210205,-14.3752183914185,
36.7667922973633,12.0868539810181,
42.7556152343750,60.2186355590820,
31.4437580108643,55.7097091674805,
15.7815084457397,0.642046451568604,
12.4858121871948,-32.8452301025391,
24.9376945495605,-5.93577384948731,
32.0283546447754,40.5423736572266,
6.96441173553467,47.9860305786133,
-39.8109207153320,20.3921909332275,
-66.0217742919922,-1.35131263732910,
-46.2589912414551,-8.09392547607422,
-9.79315567016602,-24.9053516387939,
0.771475732326508,-50.9916534423828,
-9.87240886688232,-44.3533782958984,
-8.81136226654053,6.57145309448242,
0.633710682392120,51.9925994873047,
-20.2352561950684,40.3857879638672,
-62.3256263732910,-20.4312648773193,
-66.4015274047852,-68.0332412719727,
-3.35192489624023,-61.0930099487305,
64.1284332275391,-18.6951732635498,
58.9848556518555,17.8589344024658,
-6.29298019409180,29.5028533935547,
-44.9305496215820,19.9146709442139,
-11.2969093322754,-0.958033561706543,
42.0025825500488,-21.6947593688965,
48.2293891906738,-36.4046783447266,
10.4721889495850,-38.9231491088867,
-18.5329360961914,-28.2408370971680,
-19.4527053833008,-7.20436763763428,
-8.03542518615723,12.7701206207275,
4.46133184432983,13.2547407150269,
20.3090801239014,-7.18688964843750,
34.5190734863281,-29.7274532318115,
39.1784286499023,-26.8057575225830,
41.5664291381836,7.72026443481445,
58.5394287109375,43.6353836059570,
71.7598724365234,51.5252265930176,
45.1274871826172,39.3011398315430,
-21.1660099029541,26.2329044342041,
-68.4636077880859,22.4463138580322,
-52.5909042358398,19.6462554931641,
-8.76616287231445,17.3074569702148,
1.42626941204071,23.0371074676514,
-20.4985980987549,31.3985824584961,
-25.7703914642334,20.9059658050537,
2.93729424476624,-13.5888004302979,
25.3986358642578,-42.3908081054688,
10.8273248672485,-34.7909469604492,
-11.7200431823730,0.218963623046875,
-0.0268921852111816,20.1430873870850,
33.0361671447754,6.67508745193481,
44.6952857971191,-12.8391895294189,
25.9418849945068,-0.873089075088501,
15.5113468170166,36.4409866333008,
29.0221862792969,62.0985107421875,
44.5120201110840,55.4575843811035,
35.9876670837402,27.3620719909668,
20.0021095275879,8.44010734558106,
17.1386489868164,13.5216178894043,
21.1104831695557,31.8177604675293,
14.4849624633789,44.7756614685059,
-0.699385166168213,34.8697242736816,
-4.70795392990112,2.02479934692383,
12.3327102661133,-33.4677276611328,
33.7421569824219,-44.2611618041992,
38.2054405212402,-25.0254383087158,
26.3280277252197,4.47535562515259,
6.58358287811279,24.1915073394775,
-18.3582420349121,33.8551826477051,
-40.1606063842773,36.5113792419434,
-49.8302307128906,22.4886665344238,
-52.3142890930176,-12.4309358596802,
-49.0557022094727,-46.5812759399414,
-31.4282398223877,-41.6329727172852,
11.6988496780396,5.74347639083862,
54.5527114868164,48.0344467163086,
51.2357139587402,44.0005607604981,
-3.41902089118958,5.80499315261841,
-45.8630676269531,-15.5391759872437,
-16.6136665344238,7.36369276046753,
49.0307350158691,45.8027076721191,
57.5305595397949,60.2407417297363,
-13.2044372558594,46.1720733642578,
-71.9011764526367,22.9711475372314,
-43.6144332885742,10.8804798126221,
29.1608371734619,11.3996524810791,
48.2036170959473,17.6864128112793,
-5.23925399780273,31.0545120239258,
-59.9961280822754,49.6539039611816,
-63.4947395324707,60.0946769714356,
-42.6797103881836,41.0771560668945,
-40.2952690124512,-7.70109796524048,
-40.6640548706055,-52.3023414611816,
-18.4544239044189,-55.3369522094727,
6.26082515716553,-11.7247800827026,
4.68076705932617,31.0239658355713,
-4.67993068695068,22.2793235778809,
16.5126628875732,-28.3225727081299,
47.8069152832031,-60.1369476318359,
39.1955871582031,-34.6145591735840,
0.701558828353882,22.3163700103760,
-6.44195795059204,55.7020339965820,
31.5551548004150,49.2577323913574,
47.2636756896973,28.9068851470947,
-6.07818508148193,16.8045253753662,
-71.1487197875977,4.02179765701294,
-58.2706642150879,-14.6350927352905,
16.1831626892090,-18.2245311737061,
48.6468391418457,6.71035051345825,
-1.03654384613037,31.1453914642334,
-65.7315444946289,22.7712993621826,
-73.3117294311523,-13.6057786941528,
-40.2532997131348,-33.3505706787109,
-24.2550182342529,-18.9868106842041,
-32.0261497497559,-3.06460881233215,
-22.6099624633789,-16.6994628906250,
15.8658638000488,-40.5612945556641,
48.3642616271973,-35.6056518554688,
38.4463233947754,-4.61051082611084,
-0.159832119941711,7.31856632232666,
-31.7341041564941,-16.9833488464355,
-42.2471084594727,-34.0480804443359,
-37.6095352172852,-5.05307197570801,
-21.0083179473877,43.4152030944824,
1.83523046970367,48.7984695434570,
16.8997192382813,0.238152027130127,
20.0950412750244,-46.4985275268555,
16.7634487152100,-46.7376823425293,
7.69589471817017,-21.4612255096436,
-4.82531642913818,-14.2785549163818,
-10.1432704925537,-22.4771080017090,
8.05338096618652,-8.92126274108887,
43.8983955383301,23.3691272735596,
58.8958473205566,32.6431617736816,
27.8367252349854,1.74174118041992,
-20.0254440307617,-32.1798362731934,
-26.5963897705078,-32.1533851623535,
14.0042476654053,-5.16002273559570,
47.6171226501465,14.4354286193848,
38.2156677246094,16.3195858001709,
9.03727722167969,11.9281435012817,
-1.03996539115906,5.04644727706909,
2.54357600212097,-7.02365922927856,
-7.98891687393189,-10.7420778274536,
-26.9559421539307,10.2318992614746,
-22.2471561431885,33.4761924743652,
12.2664661407471,17.4305210113525,
39.7758331298828,-28.3094062805176,
40.5229682922363,-47.4476509094238,
37.9324722290039,-16.6365928649902,
43.6972084045410,18.6132583618164,
31.9475688934326,4.73107528686523,
-15.5174350738525,-38.7340698242188,
-51.4047279357910,-45.3232383728027,
-27.4906673431397,3.70015931129456,
27.7190570831299,55.3718032836914,
42.2652091979981,59.1534538269043,
2.35548114776611,27.6906681060791,
-33.5246887207031,-0.00775516033172607,
-20.3409385681152,-8.13729476928711,
1.61527085304260,-2.42904615402222,
-16.8666954040527,12.5161085128784,
-49.5464210510254,30.3965320587158,
-38.5170593261719,30.9892292022705,
12.5293054580688,3.30244612693787,
42.9472503662109,-32.3185729980469,
37.4690971374512,-47.5714035034180,
34.5307617187500,-34.6357841491699,
53.3283271789551,-14.3479413986206,
53.0804939270020,4.73403072357178,
12.0612497329712,32.7987861633301,
-25.6683025360107,61.9380149841309,
-13.7085361480713,56.2839241027832,
22.3321990966797,11.9986600875855,
15.5907430648804,-25.3149471282959,
-37.1526489257813,-20.7114257812500,
-66.0917968750000,8.22850608825684,
-35.2074851989746,19.4240417480469,
12.2862319946289,11.1319656372070,
27.1822204589844,12.4046020507813,
19.6971702575684,24.5128784179688,
22.7089595794678,12.1629962921143,
34.4112319946289,-30.5858192443848,
33.8530464172363,-54.4686012268066,
23.8907470703125,-26.4666671752930,
23.7397766113281,8.65634250640869,
23.7122039794922,-1.47307443618774,
2.91016507148743,-38.6774978637695,
-31.2339382171631,-46.5801010131836,
-31.6602802276611,-15.9460248947144,
16.2774620056152,1.50309455394745,
62.2286872863770,-14.8213434219360,
57.7397346496582,-27.4911594390869,
14.7426328659058,-10.4053936004639,
-18.0979423522949,4.72484207153320,
-23.3275833129883,-18.1886711120605,
-16.6388702392578,-42.5707740783691,
-20.3584747314453,-13.6508970260620,
-32.8890151977539,40.2737388610840,
-41.9985122680664,42.1627693176270,
-34.9934692382813,-17.7590904235840,
-5.63204002380371,-54.6544303894043,
40.0968933105469,-16.2325172424316,
72.7537918090820,48.6141929626465,
59.2936935424805,63.1759452819824,
6.64662122726440,26.4593238830566,
-40.1067237854004,-5.45772218704224,
-49.8062744140625,-13.4376850128174,
-37.4375991821289,-28.0442008972168,
-27.9336566925049,-52.6293678283691,
-16.6552524566650,-45.9383316040039,
7.41634654998779,1.70267212390900,
35.4560470581055,34.4813995361328,
45.2130355834961,10.2732172012329,
36.8347511291504,-36.8103446960449,
36.4790306091309,-50.6905250549316,
49.5182533264160,-31.5281410217285,
44.5983085632324,-20.2909622192383,
4.00684499740601,-27.0807056427002,
-40.5612754821777,-23.4517669677734,
-48.7693634033203,6.46913528442383,
-21.8071746826172,34.1600608825684,
1.67997157573700,31.9743309020996,
9.18002223968506,17.5884075164795,
14.1838731765747,14.3909959793091,
19.4912681579590,19.0385360717773,
9.64013481140137,14.6748609542847,
-17.8241767883301,5.86266326904297,
-27.2472267150879,4.25759649276733,
1.66693687438965,1.55828893184662,
36.7337341308594,-13.6621751785278,
26.6491146087647,-31.2099437713623,
-22.0935935974121,-29.2146549224854,
-48.5451393127441,-7.99754190444946,
-26.4933757781982,6.41488599777222,
11.0879068374634,0.958299219608307,
27.3008460998535,-7.67072153091431,
26.2045516967773,0.958611547946930,
29.9319553375244,18.7673377990723,
33.5251770019531,27.6163997650147,
17.5512981414795,31.8925571441650,
-11.5425958633423,44.2416000366211,
-27.0900630950928,58.9422760009766,
-31.2812500000000,53.5729598999023,
-46.2877044677734,23.6274509429932,
-63.4279327392578,-9.65871238708496,
-45.0321502685547,-21.3438224792480,
3.91182041168213,-9.32758331298828,
25.7346248626709,6.32952737808228,
-12.6736755371094,4.27364969253540,
-55.3185005187988,-17.6585464477539,
-34.7075614929199,-42.8330535888672,
33.7999801635742,-48.7263183593750,
71.0302047729492,-25.5669517517090,
46.4802703857422,6.02158164978027,
14.5411987304688,16.7205085754395,
23.8500099182129,3.85675549507141,
45.6137619018555,-7.58238840103149,
29.0323886871338,-0.387822866439819,
-8.42459011077881,12.5969991683960,
-9.81859207153320,9.16482734680176,
34.3528861999512,1.34647095203400,
66.3005828857422,12.2668485641480,
37.8526420593262,41.3802528381348,
-21.8060512542725,50.7269287109375,
-57.8147964477539,13.6627845764160,
-52.9800262451172,-38.9680061340332,
-34.7625465393066,-51.8125991821289,
-31.0868110656738,-12.2976646423340,
-36.0870933532715,35.7812576293945,
-33.9761390686035,44.5193405151367,
-29.9221000671387,11.3160982131958,
-29.0219745635986,-26.8562984466553,
-20.5358505249023,-38.3010063171387,
11.4776182174683,-18.3053226470947,
52.9051780700684,15.4094982147217,
67.3584442138672,43.3503684997559,
31.5265388488770,49.7832527160645,
-23.9276618957520,32.0572967529297,
-41.3905868530273,9.19019412994385,
-5.94716167449951,7.44800710678101,
32.4470596313477,22.7740631103516,
21.7399406433105,26.9295330047607,
-27.8523960113525,4.60377502441406,
-58.9345436096191,-17.4797401428223,
-38.0783462524414,-13.5410175323486,
0.522776365280151,3.41718626022339,
10.7449960708618,3.72607326507568,
-6.82799196243286,-11.1037902832031,
-11.9528703689575,-6.11175680160523,
13.2739028930664,26.6160507202148,
41.6115913391113,44.2887611389160,
42.8346290588379,19.6055641174316,
20.0574932098389,-13.7391347885132,
-5.21990871429443,-7.34447145462036,
-20.8668003082275,31.0266494750977,
-30.9711093902588,50.8581161499023,
-33.8963012695313,38.4660263061523,
-20.1478977203369,23.3017978668213,
3.44423341751099,23.7125377655029,
18.8267879486084,15.4418716430664,
16.4734687805176,-17.8723144531250,
5.22207069396973,-43.0429153442383,
-1.08775413036346,-22.9117565155029,
-2.43179130554199,21.6413269042969,
-6.65329265594482,39.7903823852539,
-12.8557929992676,20.6646423339844,
-14.3289403915405,2.69335269927979,
-12.1875324249268,3.37995266914368,
-12.0595417022705,-0.126067295670509,
-13.4252233505249,-16.5274333953857,
-9.86498546600342,-17.1124000549316,
-4.86873340606689,15.1393566131592,
-11.7823200225830,49.0598983764648,
-35.6426277160645,38.4003219604492,
-54.2363204956055,-8.46991920471191,
-45.3899040222168,-35.6063156127930,
-18.9627037048340,-17.1021823883057,
-11.0161390304565,15.2090406417847,
-33.5720863342285,19.3899250030518,
-55.8501472473145,-6.26365423202515,
-42.2345504760742,-35.3140983581543,
-3.65178632736206,-51.4059410095215,
15.3510856628418,-49.0591850280762,
-4.43208885192871,-26.7142639160156,
-35.6208343505859,0.299808919429779,
-44.9713058471680,7.69270801544189,
-37.2745246887207,-18.2436580657959,
-31.6800479888916,-55.1445732116699,
-29.3858852386475,-68.2204818725586,
-15.3010253906250,-47.1140708923340,
6.00772857666016,-18.3768634796143,
10.0728988647461,-5.56773376464844,
-3.91351938247681,-3.97566151618958,
-5.17499494552612,0.238996937870979,
21.6807308197022,7.97033977508545,
53.6995697021484,13.7854480743408,
52.1264724731445,18.5429859161377,
21.2706832885742,17.1376743316650,
-4.96760988235474,0.481902599334717,
-8.71115398406982,-28.1423950195313,
-9.52491855621338,-50.5489082336426,
-24.7340259552002,-47.8554344177246,
-44.5955696105957,-29.2027492523193,
-49.0320014953613,-20.1690559387207,
-29.7294635772705,-30.9950695037842,
4.30909538269043,-44.0726661682129,
40.8893966674805,-43.8464050292969,
58.4815711975098,-34.4469795227051,
39.9970436096191,-18.9993553161621,
-5.91409158706665,4.45963191986084,
-37.9930610656738,24.3844871520996,
-20.6715946197510,13.0111579895020,
28.0687522888184,-29.6467533111572,
53.9742012023926,-57.8345794677734,
31.9112968444824,-29.7479705810547,
-2.01546621322632,30.8325443267822,
-8.81557178497315,52.6923675537109,
10.7184476852417,12.4391946792603,
26.9419097900391,-33.1182098388672,
21.3288745880127,-21.5330390930176,
1.55353879928589,30.0332527160645,
-17.9511814117432,56.6651573181152,
-30.9585037231445,39.4995613098145,
-30.6697196960449,16.2876758575439,
-10.7001905441284,11.2664871215820,
12.8110246658325,5.19698810577393,
19.0015220642090,-19.1090469360352,
4.07667350769043,-37.2144126892090,
-9.60979366302490,-20.3590946197510,
-10.9689311981201,15.1387310028076,
-17.5271186828613,29.9267711639404,
-39.1377792358398,18.1987972259522,
-48.8771133422852,4.29942989349365,
-22.1119632720947,-2.58827686309814,
20.9012489318848,-20.3828659057617,
33.0071525573731,-48.9865531921387,
0.982573986053467,-51.7509498596191,
-28.1407527923584,-16.8261928558350,
-12.0822896957397,19.9121665954590,
32.8960494995117,27.4823665618897,
57.1844711303711,15.2202587127686,
44.0004577636719,16.4025382995605,
19.9178142547607,26.9186592102051,
11.4198932647705,18.8690147399902,
14.4890184402466,-9.20413112640381,
14.9357738494873,-17.4995689392090,
6.80689287185669,15.6171607971191,
-7.07758712768555,57.3192901611328,
-17.8341217041016,65.8832702636719,
-16.0881500244141,38.2348213195801,
4.89085721969605,-1.85509371757507,
36.2290077209473,-34.9150810241699,
55.4101295471191,-50.7392349243164,
50.5131607055664,-39.2503433227539,
38.0644645690918,-0.618785858154297,
36.6282463073731,36.2277259826660,
40.3409881591797,45.8609733581543,
34.3360061645508,33.8548927307129,
24.6151943206787,34.2311744689941,
25.5329189300537,52.3885917663574,
29.3682289123535,54.0980606079102,
12.5299730300903,22.2128067016602,
-24.8021430969238,-13.7452869415283,
-45.0546569824219,-20.1648559570313,
-22.8209342956543,-11.5081853866577,
13.3549661636353,-20.1261978149414,
15.1537542343140,-39.2452697753906,
-18.0360889434814,-39.8440628051758,
-36.5631980895996,-11.0703754425049,
-11.1038389205933,13.2223367691040,
30.6305274963379,15.8778104782105,
47.3020820617676,21.2946605682373,
33.4775581359863,44.9548263549805,
9.30932712554932,61.3032188415527,
-11.9933996200562,34.4227447509766,
-32.9418525695801,-19.1104545593262,
-49.3965606689453,-50.3925971984863,
-47.4293785095215,-46.1769218444824,
-29.7435874938965,-33.9405899047852,
-13.9938554763794,-27.2760810852051,
-9.99342155456543,-7.13375139236450,
-10.8463478088379,31.9318523406982,
-14.6343069076538,53.5068092346191,
-32.6672897338867,20.1377296447754,
-56.8832740783691,-45.6384391784668,
-53.5537376403809,-83.4072418212891,
-6.57798576354981,-62.1561203002930,
44.8511199951172,-11.4483146667480,
51.4807853698731,26.9236602783203,
10.3288822174072,36.8299560546875,
-28.9361209869385,22.1021804809570,
-25.6563529968262,-11.5271320343018,
1.22122883796692,-46.2117958068848,
14.9219379425049,-60.1592330932617,
6.96218967437744,-47.3641967773438,
1.50635766983032,-26.0369930267334,
7.97955942153931,-16.6304759979248,
14.3307027816772,-17.2578830718994,
6.21681308746338,-14.8027086257935,
-10.2634010314941,-9.56192493438721,
-21.7261333465576,-17.0086555480957,
-17.2990913391113,-35.2566795349121,
5.45524930953980,-41.0993003845215,
39.1764259338379,-25.0709686279297,
61.5532951354981,-2.76898789405823,
53.6111450195313,14.1139516830444,
13.6155891418457,26.5154209136963,
-30.3082962036133,37.8782157897949,
-48.4494400024414,36.0431327819824,
-39.3996086120606,18.2320327758789,
-22.1968402862549,7.60911893844605,
-13.0624284744263,24.3472957611084,
-12.9817190170288,48.6092720031738,
-21.8738193511963,35.4316368103027,
-33.0624504089356,-19.2604217529297,
-33.9036254882813,-64.6515274047852,
-12.0811347961426,-54.7930450439453,
24.1531505584717,-13.9388303756714,
45.3494644165039,3.33038091659546,
37.9071846008301,-20.7136993408203,
22.8255577087402,-46.9792442321777,
30.5318222045898,-40.1646499633789,
58.3786621093750,-3.08616113662720,
73.1312866210938,32.3353729248047,
49.8550949096680,48.6263313293457,
4.96823930740356,49.2354316711426,
-33.8004608154297,41.7604141235352,
-53.2563095092773,31.2670269012451,
-63.4340286254883,22.1496677398682,
-68.6751556396484,14.8615560531616,
-60.8397979736328,-3.83855962753296,
-33.4980583190918,-37.8380813598633,
6.01172161102295,-65.4190139770508,
40.9652137756348,-64.2893676757813,
55.1844902038574,-40.5036621093750,
48.1439094543457,-12.5607013702393,
32.1673278808594,9.19955158233643,
17.8134803771973,31.8973617553711,
11.6865873336792,52.4254455566406,
10.5680284500122,49.8032608032227,
5.97291803359985,21.8364658355713,
-12.3826351165771,2.82361054420471,
-42.5108337402344,16.0358085632324,
-69.7776107788086,28.3722972869873,
-68.0216827392578,-3.58527994155884,
-28.4828166961670,-61.0778427124023,
20.8737392425537,-75.2016448974609,
35.4060668945313,-24.9808902740479,
8.86078166961670,28.2377223968506,
-19.2112083435059,19.0494041442871,
-10.3525943756104,-31.7885875701904,
22.6782913208008,-50.9839248657227,
30.8846359252930,-10.5178842544556,
-4.00033330917358,39.4975662231445,
-47.7578353881836,48.4331092834473,
-59.6162414550781,23.9602108001709,
-41.0786056518555,-2.72849488258362,
-22.1040611267090,-19.6259250640869,
-11.4305553436279,-28.3987960815430,
2.50951647758484,-19.0150547027588,
19.4888458251953,11.4813251495361,
19.7313308715820,32.9771499633789,
-2.98778676986694,16.1032428741455,
-22.6112365722656,-22.6498508453369,
-7.30424070358276,-37.9061164855957,
29.8382797241211,-13.2643690109253,
42.4809074401856,16.7346878051758,
12.1197776794434,22.9797668457031,
-33.5538635253906,20.4494915008545,
-54.4831085205078,32.6603622436523,
-45.9149169921875,43.6447753906250,
-30.3828563690186,26.9654884338379,
-14.3168249130249,-5.66846275329590,
17.4885749816895,-15.8588056564331,
55.5363998413086,10.5814914703369,
62.8119468688965,42.8436813354492,
20.9243412017822,50.5871849060059,
-29.5448017120361,39.6185760498047,
-33.0567970275879,33.4480857849121,
7.54946327209473,35.0127639770508,
28.7495784759522,28.9807205200195,
-8.10517120361328,8.34713268280029,
-62.7612342834473,-13.1153707504272,
-70.9990463256836,-21.1943416595459,
-30.9467582702637,-15.6153745651245,
3.72849130630493,-3.66224765777588,
-4.21391439437866,2.65825867652893,
-32.4420089721680,1.04380691051483,
-38.0772094726563,-4.54854106903076,
-24.3277397155762,-2.23860001564026,
-21.3331623077393,11.0480613708496,
-40.9817924499512,22.0375499725342,
-56.6744232177734,17.0914268493652,
-40.7557563781738,-6.69395256042481,
-3.29226112365723,-31.5632743835449,
25.1057376861572,-37.0292167663574,
25.1372604370117,-22.9230556488037,
7.45081138610840,-1.37143373489380,
-2.43673443794251,14.4846839904785,
4.48567390441895,23.6839351654053,
16.9093742370605,31.0125389099121,
19.2701568603516,39.0937919616699,
3.80554294586182,45.9465141296387,
-20.6391696929932,41.5879898071289,
-40.8373374938965,15.8329267501831,
-42.8837966918945,-26.9130649566650,
-23.9209365844727,-64.5770721435547,
7.60029697418213,-69.3910980224609,
33.8702163696289,-35.4863853454590,
38.5181312561035,9.32680702209473,
21.4526996612549,32.6314163208008,
1.27688598632813,23.1123962402344,
-8.70218181610107,1.89805424213409,
-3.82899689674377,-11.1651659011841,
8.94975471496582,-10.0227642059326,
23.5330886840820,0.720834195613861,
35.3791580200195,18.0826015472412,
32.6294288635254,37.5791854858398,
6.11154842376709,43.6051826477051,
-31.7853431701660,22.6179523468018,
-53.7256164550781,-15.1991939544678,
-36.9899024963379,-38.1264419555664,
11.6822738647461,-25.8623943328857,
53.3231353759766,10.9127817153931,
55.9574050903320,44.5116767883301,
15.3365659713745,55.1140594482422,
-36.3151817321777,44.3459243774414,
-58.4861869812012,14.8250541687012,
-34.6367683410645,-26.6338443756104,
12.4205760955811,-64.1244201660156,
38.8396034240723,-76.6193237304688,
23.2606487274170,-55.0588722229004,
-10.4339075088501,-17.0865268707275,
-19.9313468933105,8.85205268859863,
8.52572727203369,6.68576192855835,
42.0146179199219,-12.8917522430420,
39.8612556457520,-28.2213764190674,
1.50824213027954,-28.3866729736328,
-38.4201583862305,-14.9791164398193,
-48.4195442199707,-1.51493871212006,
-39.8659400939941,-2.55104613304138,
-37.7831649780273,-14.2539625167847,
-46.6297760009766,-20.9228038787842,
-49.6538658142090,-13.7564668655396,
-32.3587493896484,1.45603072643280,
-8.92788696289063,10.0099973678589,
-2.41553115844727,10.5568294525146,
-6.99551820755005,6.86675214767456,
-1.82577311992645,-2.96091461181641,
16.3755435943604,-26.3330192565918,
27.1427612304688,-53.7551727294922,
15.8306703567505,-53.1720581054688,
-7.25298500061035,-13.4579868316650,
-20.4045639038086,28.0435714721680,
-29.1865501403809,30.4116859436035,
-45.3410758972168,-2.62605023384094,
-58.1975555419922,-26.0533790588379,
-41.8064270019531,-18.0692443847656,
4.31289577484131,-2.65377616882324,
34.0980415344238,-3.76297116279602,
18.6406898498535,-4.38697147369385,
-17.2419128417969,15.1645994186401,
-31.3206214904785,35.8410224914551,
-21.9913444519043,19.0480957031250,
-14.7625217437744,-29.4636936187744,
-15.9415416717529,-58.1009521484375,
-2.20918250083923,-41.7519111633301,
32.3895263671875,-15.0168209075928,
56.2200775146484,-21.3323936462402,
51.6220932006836,-50.0290756225586,
37.6102981567383,-55.1792678833008,
33.4184646606445,-25.9536056518555,
16.9960289001465,8.08498382568359,
-25.5985984802246,12.4949321746826,
-60.8838768005371,-11.2500772476196,
-38.2017745971680,-34.1484909057617,
26.3496589660645,-40.4778823852539,
60.2506790161133,-31.6121177673340,
32.4672012329102,-13.6160850524902,
-5.67497920989990,5.04385757446289,
3.87951064109802,13.6948060989380,
39.3860435485840,11.1255064010620,
35.3471908569336,3.39725756645203,
-18.0124645233154,-9.71249198913574,
-61.2128486633301,-27.8617668151855,
-48.4244155883789,-33.5479621887207,
-12.0878057479858,-7.96136713027954,
-12.8841924667358,37.6528244018555,
-49.9231986999512,54.4582443237305,
-66.9971008300781,10.6198387145996,
-33.2474632263184,-52.4926605224609,
17.6218452453613,-58.1734695434570,
32.1217994689941,-3.37412261962891,
5.06941699981689,34.4212379455566,
-11.7377662658691,5.29458999633789,
12.7314252853394,-42.1935005187988,
45.5902099609375,-27.7625503540039,
41.7737083435059,34.9324302673340,
6.06334209442139,60.1733665466309,
-11.7168989181519,14.3892793655396,
9.88711547851563,-36.8147125244141,
34.6700439453125,-28.1695938110352,
20.1839885711670,12.8127374649048,
-18.9153060913086,15.8554363250732,
-26.5077934265137,-16.2231597900391,
9.13362884521484,-19.5628585815430,
42.0230941772461,25.8743953704834,
30.5324249267578,66.8949279785156,
-9.83330249786377,54.3609886169434,
-33.8917198181152,11.1486387252808,
-25.6749649047852,-20.9237766265869,
-6.38950824737549,-33.6894874572754,
5.62453460693359,-41.8806152343750,
13.1515893936157,-41.9460182189941,
18.1323070526123,-17.0948524475098,
9.27904796600342,21.9118690490723,
-11.7738962173462,43.1551856994629,
-21.5826339721680,40.1033058166504,
-0.707630634307861,38.5382957458496,
32.3067703247070,44.6692543029785,
42.3360595703125,32.8575363159180,
22.2007923126221,-4.69560623168945,
1.97905540466309,-35.3460121154785,
7.85406112670898,-36.0985260009766,
23.7698059082031,-26.2355575561523,
18.6440296173096,-30.8077144622803,
-7.90945243835449,-41.1236610412598,
-23.1754474639893,-24.6705398559570,
-10.1615819931030,16.7761955261230,
6.55911254882813,42.6617240905762,
1.91476130485535,31.2814674377441,
-12.7693834304810,7.34216165542603,
-10.1179924011230,6.65344524383545,
3.07960319519043,25.0351810455322,
-3.87697005271912,36.4683341979981,
-31.8949604034424,27.2779159545898,
-39.4739074707031,2.84351968765259,
-2.30770206451416,-22.6774387359619,
39.2934570312500,-38.9980430603027,
34.0330505371094,-34.1614303588867,
-7.66841316223145,-9.96382999420166,
-25.7120590209961,11.7759847640991,
-2.16518020629883,10.8344860076904,
21.6503410339355,-4.39855337142944,
13.7880687713623,-8.15448665618897,
-9.90114212036133,8.38061809539795,
-22.1684665679932,20.6885070800781,
-29.6872158050537,1.14678287506104,
-44.6351928710938,-34.8206291198731,
-47.4274024963379,-54.2229118347168,
-15.2313671112061,-43.3243522644043,
25.8258934020996,-21.0239181518555,
24.6557159423828,-12.3145275115967,
-11.1076946258545,-21.3563117980957,
-25.4932727813721,-26.7633113861084,
-2.02305030822754,-14.0690927505493,
9.08988666534424,9.35351276397705,
-22.1298408508301,18.2072486877441,
-48.8422927856445,-3.40563249588013,
-17.3880481719971,-36.0584297180176,
43.7856178283691,-39.5373344421387,
62.5534629821777,2.62717437744141,
30.4716053009033,59.5110282897949,
9.14124107360840,82.6975326538086,
24.6157054901123,54.3474121093750,
26.7802276611328,6.19393348693848,
-17.4449615478516,-18.5397090911865,
-58.8779182434082,-12.0612010955811,
-27.6487617492676,2.76687216758728,
52.4167938232422,-2.36667537689209,
84.7567062377930,-25.3982696533203,
32.5966529846191,-42.8385391235352,
-31.4985942840576,-36.1745605468750,
-29.4882068634033,-13.7834911346436,
26.3789691925049,-3.60510206222534,
53.3303718566895,-17.3823204040527,
17.1656074523926,-32.5122909545898,
-29.2373256683350,-18.2102928161621,
-22.8057842254639,20.6746063232422,
16.5087795257568,43.1870803833008,
26.2353305816650,25.7929363250732,
-11.5078792572021,-14.5017280578613,
-46.2233123779297,-38.0902175903320,
-28.3271369934082,-36.3453903198242,
22.9797782897949,-28.0054531097412,
40.4991073608398,-19.3018436431885,
-0.278019428253174,0.356420278549194,
-42.6035919189453,26.4803447723389,
-25.8823528289795,34.1770935058594,
33.6014289855957,10.0757150650024,
71.8802795410156,-22.2786426544189,
54.7077941894531,-29.0034770965576,
19.0490322113037,-12.7853412628174,
21.3025684356689,2.59565901756287,
53.0034599304199,7.52991628646851,
53.2124862670898,15.6668663024902,
1.81912016868591,30.7176132202148,
-46.0644149780273,32.0402946472168,
-33.7802085876465,2.32172298431397,
17.0588150024414,-33.8446540832520,
37.3129577636719,-35.4861602783203,
3.99506306648254,2.49862623214722,
-30.7650432586670,45.0733566284180,
-21.7652301788330,49.0517616271973,
1.31105053424835,11.7369079589844,
-12.0423612594605,-33.5141868591309,
-44.9799652099609,-48.0750045776367,
-39.1941032409668,-20.8961200714111,
14.3018035888672,22.8470382690430,
53.7062072753906,44.4280662536621,
36.9106788635254,26.6348247528076,
0.108453303575516,-11.4409255981445,
-6.52601099014282,-29.8220882415772,
5.40361976623535,-11.5476093292236,
-3.69401359558105,19.3695392608643,
-27.8969268798828,26.1395454406738,
-23.7116889953613,-0.952596902847290,
14.6271476745605,-34.0413398742676,
34.7635536193848,-43.7401618957520,
4.17886209487915,-30.5614528656006,
-38.7158889770508,-19.8622817993164,
-45.6105117797852,-24.7210941314697,
-24.2210121154785,-29.2589721679688,
-6.60696887969971,-18.3926162719727,
6.09124994277954,0.00280094146728516,
30.4790229797363,8.16122341156006,
51.7237815856934,3.58395481109619,
45.7811851501465,3.41067147254944,
21.8111629486084,14.3414106369019,
15.1343688964844,11.4903659820557,
31.7442169189453,-19.2516555786133,
33.1126747131348,-48.2627677917481,
0.638192176818848,-40.4491996765137,
-28.0444049835205,-2.94560861587524,
-15.5225963592529,16.6843585968018,
15.6966266632080,-0.910169601440430,
20.5943050384522,-22.3237762451172,
2.22488832473755,-13.7685518264771,
-5.05546712875366,8.73788166046143,
8.89669418334961,5.72492122650147,
23.5874423980713,-19.3292694091797,
26.4528770446777,-31.9612541198730,
33.8596000671387,-24.8156414031982,
51.2032127380371,-27.7688026428223,
51.6307601928711,-47.3807868957520,
22.2259159088135,-44.1958312988281,
-10.1938447952271,2.93353080749512,
-11.3837795257568,53.1367721557617,
9.34138488769531,53.3154449462891,
13.8769741058350,17.0260372161865,
-0.239334762096405,2.29831361770630,
-2.10655713081360,26.9147548675537,
22.9056320190430,47.7170333862305,
45.2293052673340,25.2200202941895,
31.6088771820068,-13.7575225830078,
-6.96437072753906,-24.3846378326416,
-33.2013702392578,-9.75244808197022,
-29.4477443695068,-4.67697429656982,
-18.5130577087402,-16.9629478454590,
-24.7936096191406,-24.1493282318115,
-41.4035453796387,-16.8379631042480,
-42.2629737854004,-8.18817234039307,
-14.8749694824219,-12.1405010223389,
20.4583435058594,-18.3148803710938,
41.8862342834473,-14.6986522674561,
49.6326866149902,-4.63925743103027,
54.1641845703125,9.41528034210205,
55.7225112915039,34.0291519165039,
39.4351730346680,64.9574432373047,
0.208747982978821,73.9389266967773,
-39.2970046997070,41.9910087585449,
-52.2488365173340,-0.321985244750977,
-46.5131111145020,-8.82825851440430,
-44.0082511901856,15.6905269622803,
-46.4698524475098,22.3231277465820,
-34.9793319702148,-19.3660545349121,
-4.78058862686157,-71.7014923095703,
13.6173973083496,-78.8279113769531,
1.42834222316742,-38.2760467529297,
-19.2229003906250,-5.74672937393189,
-4.49386692047119,-18.6130485534668,
39.1858024597168,-50.0117149353027,
60.1528739929199,-45.0079956054688,
30.8646888732910,1.43061161041260,
-15.4876728057861,40.6485519409180,
-23.1392002105713,36.5979118347168,
12.1587409973145,10.3633155822754,
45.1722259521484,5.50691127777100,
38.8645515441895,31.7351226806641,
7.90715074539185,47.7765159606934,
-14.3876056671143,22.0336685180664,
-19.9145889282227,-23.0944328308105,
-23.7551460266113,-47.2524147033691,
-25.0504245758057,-43.7352066040039,
-2.66113138198853,-38.3184051513672,
43.8083305358887,-39.7436065673828,
77.3930130004883,-28.3548564910889,
60.9377975463867,9.22006797790527,
7.81279850006104,44.5535850524902,
-30.1162757873535,36.3809165954590,
-30.4999046325684,-11.4832401275635,
-22.3590984344482,-44.4844932556152,
-34.7117118835449,-28.8641662597656,
-49.8276100158691,11.7029409408569,
-33.2435951232910,27.7277603149414,
11.5483016967773,4.04808616638184,
38.6365432739258,-29.3003425598145,
34.5588378906250,-39.2633934020996,
31.2900295257568,-29.6396694183350,
53.3495063781738,-17.2661972045898,
69.4125823974609,0.182991504669189,
34.1631660461426,34.1137046813965,
-41.2007713317871,66.9781494140625,
-93.5504455566406,61.4810371398926,
-80.8642578125000,18.1524581909180,
-25.7744674682617,-16.0424365997314,
19.3929843902588,-2.08434319496155,
33.8785133361816,34.4307479858398,
31.7718448638916,37.7838706970215,
30.2425842285156,6.39552307128906,
35.7945327758789,-10.0599927902222,
44.5031127929688,11.7833147048950,
49.6897697448731,33.7860603332520,
46.8082237243652,15.9172601699829,
37.6096038818359,-12.4572811126709,
31.0869007110596,3.60827207565308,
30.4554805755615,54.0165443420410,
23.0837554931641,75.6510620117188,
-2.80050945281982,36.3752365112305,
-37.2725181579590,-22.3258876800537,
-50.0944175720215,-41.2070236206055,
-27.2695350646973,-20.4070587158203,
8.85357093811035,3.79515981674194,
27.6668968200684,7.82671451568604,
19.1558208465576,-1.66445803642273,
5.24269580841064,-16.2083816528320,
7.06509304046631,-29.4795608520508,
19.8486862182617,-27.8060989379883,
19.9895381927490,1.75930142402649,
-3.01266503334045,36.7032012939453,
-30.0804405212402,31.8026256561279,
-36.5769424438477,-12.1663856506348,
-26.7077999114990,-43.1378211975098,
-21.9650707244873,-17.9154796600342,
-29.3120021820068,40.0448455810547,
-28.6770172119141,69.1409759521484,
-5.83202743530273,46.2718353271484,
16.9441928863525,13.6371011734009,
9.29952526092529,16.6236534118652,
-23.5376243591309,41.3035888671875,
-40.1590652465820,45.2526092529297,
-15.5465679168701,10.5611124038696,
26.8118324279785,-34.7262802124023,
45.9162940979004,-49.0713500976563,
31.8865375518799,-21.5543365478516,
9.34900951385498,26.0633621215820,
-0.318086981773376,59.0284080505371,
4.08295631408691,56.6799774169922,
9.55690097808838,27.2134838104248,
3.68599939346313,-4.31790828704834,
-18.2781105041504,-22.2775917053223,
-44.3224449157715,-29.0643119812012,
-48.5036430358887,-39.5964126586914,
-17.2445907592773,-58.5686225891113,
22.9405517578125,-64.4119186401367,
31.5304107666016,-45.5561981201172,
1.86225283145905,-12.1748704910278,
-24.4837703704834,8.91958618164063,
-10.7020854949951,3.67263913154602,
23.7142181396484,-20.8481292724609,
29.6206493377686,-40.4405860900879,
-2.54583239555359,-42.0718879699707,
-30.2456970214844,-31.0966300964355,
-21.6810607910156,-21.0689735412598,
9.42662620544434,-26.2556514739990,
28.6807823181152,-40.4864311218262,
26.0875911712647,-41.5345802307129,
18.3535900115967,-11.9862356185913,
10.9384508132935,35.3207092285156,
-4.74247932434082,65.0313110351563,
-25.6909294128418,53.6445312500000,
-32.2359886169434,20.6084384918213,
-8.66169357299805,3.08552503585815,
29.4804267883301,6.09743356704712,
53.2814521789551,7.49903488159180,
50.9341812133789,-13.5200929641724,
30.1111965179443,-41.8414611816406,
5.57544422149658,-44.1332168579102,
-15.5733232498169,-14.3030090332031,
-24.2808742523193,18.9054985046387,
-16.0251770019531,24.3909149169922,
7.35703706741333,1.75053691864014,
30.8709125518799,-23.3496913909912,
40.5085105895996,-20.0972232818604,
35.6336517333984,19.5106830596924,
22.3017578125000,70.6930160522461,
6.13772249221802,88.0300369262695,
-16.1132812500000,46.1372299194336,
-38.3100242614746,-20.7944908142090,
-37.2948799133301,-55.0600700378418,
-1.58811378479004,-30.7181701660156,
45.2200698852539,17.8925933837891,
56.7007904052734,40.6643486022949,
16.1724300384522,26.4726638793945,
-37.1551055908203,1.48960864543915,
-55.8250122070313,-18.9104919433594,
-40.3455581665039,-43.2597351074219,
-29.9023208618164,-63.3237495422363,
-42.4504394531250,-59.7366600036621,
-46.2706642150879,-30.5753898620605,
-12.9276628494263,-1.79489970207214,
35.1338043212891,7.90030908584595,
49.9289321899414,13.3878307342529,
21.8606681823730,30.0003395080566,
-13.2166576385498,36.0801162719727,
-23.9984283447266,12.3703107833862,
-15.9425487518311,-15.6901817321777,
-13.3681774139404,-5.85700416564941,
-24.1753635406494,34.5132713317871,
-38.7273559570313,42.1692504882813,
-48.4643516540527,-7.60519886016846,
-43.8934707641602,-54.5530052185059,
-20.2902202606201,-36.1960716247559,
12.5513544082642,29.0718765258789,
32.2578125000000,65.7048110961914,
18.2425346374512,41.7312469482422,
-12.6738367080688,0.775760769844055,
-29.1766796112061,-8.49549388885498,
-18.3016319274902,8.54274463653565,
-3.32089996337891,13.3638038635254,
-4.65783977508545,-5.00555515289307,
-14.7288846969605,-29.7289867401123,
-8.85480117797852,-43.0369873046875,
18.8865623474121,-41.7111816406250,
43.9189643859863,-23.1143760681152,
40.8518371582031,7.65606212615967,
12.6320552825928,29.0669021606445,
-10.8559951782227,17.5955371856689,
-8.08252239227295,-14.2054920196533,
16.2300624847412,-33.3515434265137,
38.3984184265137,-26.1190853118897,
46.5971374511719,-11.9405517578125,
44.9088134765625,-16.5987224578857,
40.7852363586426,-33.1268196105957,
30.6696739196777,-29.0315570831299,
8.08567237854004,-0.380472660064697,
-18.1942729949951,26.3654899597168,
-27.2787113189697,29.3335647583008,
-10.7800025939941,14.5812406539917,
10.0406570434570,3.55203914642334,
13.3130588531494,13.1603240966797,
-2.29500889778137,36.3464851379395,
-12.9960222244263,56.0269813537598,
-0.731922924518585,54.5790252685547,
23.6795463562012,32.5893173217773,
37.2738342285156,10.0960006713867,
30.8234443664551,9.00677680969238,
16.6310138702393,23.6779098510742,
9.10432624816895,24.1344051361084,
11.4913520812988,-6.09118366241455,
16.5019245147705,-41.1704940795898,
18.8138828277588,-42.2724113464356,
11.1848726272583,-7.83913707733154,
-8.10596942901611,15.3419256210327,
-38.4582824707031,-1.78193807601929,
-61.5020294189453,-37.6908378601074,
-61.8804435729981,-50.6510047912598,
-42.0732231140137,-28.8938827514648,
-23.4933471679688,-4.90121936798096,
-17.0669689178467,-10.8048000335693,
-11.4485168457031,-37.0755653381348,
6.58616542816162,-49.8010940551758,
28.8938751220703,-31.0329570770264,
33.3034629821777,2.68816614151001,
20.1177310943604,19.9559955596924,
10.8055524826050,4.66173458099365,
15.9859437942505,-22.0959262847900,
16.8532238006592,-19.6046447753906,
-8.34494876861572,25.6014041900635,
-47.8580513000488,71.6056747436523,
-66.2423095703125,58.9830017089844,
-50.4103393554688,-11.5976076126099,
-27.4047470092773,-69.8936004638672,
-24.6287479400635,-57.1268272399902,
-33.9764671325684,0.498518407344818,
-28.8326454162598,19.9379444122314,
1.78791403770447,-21.3196258544922,
35.2362022399902,-62.6727714538574,
40.8342361450195,-49.4007949829102,
16.7467117309570,-9.72032165527344,
-9.67056941986084,-5.97590065002441,
-11.4452638626099,-41.4709739685059,
11.6679801940918,-55.9226112365723,
33.1606445312500,-19.5511875152588,
28.0222301483154,25.2039070129395,
3.41412973403931,25.5123939514160,
-4.84831857681274,-4.71516704559326,
24.8308467864990,-19.6595153808594,
61.4853744506836,-8.37414264678955,
58.5939216613770,-2.60355472564697,
16.8523788452148,-24.8196620941162,
-16.1849060058594,-48.7483024597168,
-0.0735917091369629,-40.3847885131836,
42.4834556579590,-5.40275096893311,
53.4607696533203,23.3125000000000,
15.2973499298096,26.1410694122314,
-31.7983894348145,7.15031623840332,
-48.5495452880859,-13.4748430252075,
-31.2337169647217,-23.3172931671143,
0.792310655117035,-19.0661926269531,
34.2436485290527,1.22432589530945,
53.4336204528809,36.8032836914063,
35.4427108764648,67.1736373901367,
-21.5202064514160,68.2660064697266,
-70.1342239379883,36.8720207214356,
-56.7447700500488,-6.01451063156128,
9.18192291259766,-23.2262344360352,
59.5034141540527,0.474596977233887,
46.9701919555664,33.7622184753418,
1.14414310455322,31.4177665710449,
-20.4485588073730,-11.1803655624390,
-3.32927846908569,-45.2450218200684,
20.7382259368897,-27.5245704650879,
31.2021141052246,23.5498409271240,
31.9137630462647,45.1469917297363,
25.6781864166260,9.77794933319092,
5.43542480468750,-36.5720939636231,
-22.1615009307861,-39.2620010375977,
-32.9962768554688,-7.77354717254639,
-16.1574726104736,-0.591161251068115,
6.89737987518311,-36.4854774475098,
14.3705015182495,-65.4228439331055,
14.8350639343262,-44.8167419433594,
30.2582530975342,9.56271743774414,
54.7288589477539,44.4302482604981,
57.9017601013184,45.0938339233398,
37.8849143981934,38.9408378601074,
13.6050767898560,38.6827354431152,
-1.26992094516754,26.5582141876221,
-4.14395427703857,-5.81055879592896,
7.84692287445068,-33.2507896423340,
37.0087699890137,-30.7960109710693,
61.3018875122070,-13.0362796783447,
48.1512489318848,-12.1820154190063,
3.75267934799194,-27.5877418518066,
-20.7702827453613,-32.6475028991699,
5.71533536911011,-24.1688117980957,
39.3898925781250,-20.3557987213135,
19.8712139129639,-32.9338836669922,
-33.3250846862793,-43.9456748962402,
-45.2805976867676,-37.1872558593750,
6.44092655181885,-16.5658264160156,
55.4660110473633,-2.05650043487549,
39.2528877258301,2.98845505714417,
-14.3725500106812,6.24891042709351,
-40.2105407714844,8.78863906860352,
-31.2297840118408,8.37841701507568,
-29.6201725006104,7.53638792037964,
-47.4317436218262,7.22827625274658,
-41.4625167846680,-5.69554376602173,
11.1011524200439,-32.1534423828125,
65.9822082519531,-49.2547302246094,
67.9127502441406,-28.0968513488770,
32.2083892822266,20.0842075347900,
13.0449285507202,55.1569709777832,
29.4567451477051,51.0049209594727,
49.3994178771973,27.8244228363037,
41.1270294189453,21.4205741882324,
8.52541160583496,31.6907558441162,
-21.2539443969727,30.4246520996094,
-24.8735561370850,10.4213390350342,
2.88685274124146,-12.5208721160889,
43.6829605102539,-26.7106742858887,
61.7736473083496,-36.0742835998535,
29.7026329040527,-40.0900115966797,
-25.8948211669922,-34.5966987609863,
-42.7627029418945,-26.2488536834717,
2.46578121185303,-36.7849731445313,
56.9779510498047,-61.0046539306641,
57.2038955688477,-55.2959861755371,
12.4065685272217,1.86527276039124,
-22.0289916992188,66.7906570434570,
-16.3380374908447,71.2376785278320,
3.42315149307251,12.8565540313721,
2.64459180831909,-33.4537467956543,
-12.7011060714722,-18.4483261108398,
-18.4293956756592,21.2348518371582,
-17.5597763061523,27.2973270416260,
-21.6042022705078,0.534321784973145,
-21.6903400421143,-9.47184944152832,
-6.41069030761719,21.7670421600342,
15.1605644226074,56.5539283752441,
22.3381233215332,55.8809700012207,
20.6267242431641,23.3614616394043,
31.6746520996094,-6.10985660552979,
46.8374137878418,-16.8198204040527,
30.4497489929199,-11.1471242904663,
-17.5912647247314,2.01213407516480,
-46.3973693847656,11.7139377593994,
-15.5429506301880,7.14809226989746,
43.5994758605957,-2.91274118423462,
57.8451881408691,10.2563314437866,
11.8068733215332,51.7775421142578,
-32.5947914123535,80.3213043212891,
-24.1502761840820,55.4305839538574,
18.5391712188721,-6.76791763305664,
35.2870254516602,-47.1211700439453,
5.47813224792481,-39.0931396484375,
-30.8780918121338,-19.8956966400147,
-28.5597057342529,-31.0394477844238,
11.5767202377319,-48.5027122497559,
43.4434890747070,-29.4143104553223,
30.6290035247803,20.0484161376953,
-19.4207534790039,50.3853187561035,
-58.3276977539063,39.6900482177734,
-48.4993438720703,19.5139789581299,
1.03171718120575,25.8846759796143,
42.6286582946777,52.0587463378906,
31.9003906250000,64.8461990356445,
-23.9526653289795,52.7211875915527,
-73.0192947387695,26.6009769439697,
-79.2253265380859,0.0916827917098999,
-45.8443107604981,-14.8388462066650,
-4.67243576049805,-2.87743258476257,
19.2859878540039,35.7928619384766,
22.1708946228027,64.7802200317383,
18.1871433258057,46.1809196472168,
16.7229690551758,-4.69156217575073,
22.6983261108398,-27.2745971679688,
29.5912857055664,2.43654274940491,
17.7859287261963,39.5026550292969,
-13.5190219879150,28.7336025238037,
-37.5849876403809,-26.2075538635254,
-25.3527259826660,-66.3473815917969,
21.7884826660156,-55.8033905029297,
58.5191040039063,-17.3537483215332,
41.7657814025879,10.9451551437378,
-12.2495403289795,24.6183414459229,
-52.1201171875000,37.5559310913086,
-48.5203018188477,50.6007995605469,
-25.0482730865479,46.1419715881348,
-23.6331405639648,14.8721437454224,
-45.2147674560547,-24.0786457061768,
-47.9526023864746,-43.9782905578613,
-5.75013303756714,-29.2233581542969,
48.8747596740723,5.30752611160278,
60.9898109436035,31.3786678314209,
16.9261455535889,28.2454109191895,
-31.4395236968994,-0.493956923484802,
-29.3126602172852,-33.4421463012695,
21.3559360504150,-49.1002960205078,
63.4098472595215,-43.6354370117188,
52.1067619323731,-30.5434551239014,
5.75639343261719,-16.1228446960449,
-27.1356163024902,-0.481801509857178,
-30.1821918487549,16.4412631988525,
-26.3588504791260,29.4650306701660,
-38.3726119995117,33.9504547119141,
-53.3342628479004,32.5799446105957,
-41.6037826538086,28.5520896911621,
-5.14343547821045,27.3983039855957,
25.8508567810059,29.3256111145020,
30.5252075195313,32.1408615112305,
23.5696411132813,30.2652606964111,
28.1369113922119,16.9506034851074,
41.9700202941895,-8.13903713226318,
38.3893661499023,-27.4101600646973,
5.46244525909424,-25.0618801116943,
-34.4811019897461,-3.25573062896729,
-49.2428665161133,14.1900281906128,
-38.5974349975586,12.8145351409912,
-26.7263050079346,4.34091520309448,
-31.3753623962402,9.06868076324463,
-41.1731376647949,22.1253223419189,
-34.3838386535645,19.9473857879639,
-9.29208087921143,-5.59577465057373,
12.5951051712036,-26.1190071105957,
13.3877658843994,-15.0916767120361,
-2.15543031692505,9.90857315063477,
-21.5628318786621,6.82360887527466,
-31.6519756317139,-36.1774749755859,
-24.6291770935059,-79.7159347534180,
1.64976441860199,-81.7867813110352,
32.4809989929199,-39.8827400207520,
46.2671051025391,11.2191467285156,
26.3097000122070,39.1963729858398,
-8.82439327239990,34.3123321533203,
-25.2323913574219,8.41827106475830,
-13.6451568603516,-15.6609029769897,
0.278916060924530,-14.6772041320801,
-11.3206787109375,17.5696430206299,
-41.2677650451660,53.4627723693848,
-54.1838607788086,61.3875923156738,
-30.9992237091064,39.5377693176270,
4.32254600524902,14.1715431213379,
14.5286369323730,-4.13607597351074,
-4.44247961044312,-27.0329303741455,
-19.6868991851807,-57.8445739746094,
0.977948427200317,-68.6116943359375,
46.4885711669922,-40.1497154235840,
74.3538665771484,4.32928991317749,
60.1635513305664,17.4916381835938,
27.5091915130615,-3.46236968040466,
20.7255802154541,-14.4800624847412,
41.8950386047363,11.1735095977783,
46.9661026000977,49.1067466735840,
7.13618230819702,56.8754081726074,
-51.4072952270508,33.7447013854981,
-76.0099868774414,12.0078573226929,
-49.2889213562012,5.31715202331543,
-11.7575407028198,-6.25130224227905,
-6.28315305709839,-31.7044830322266,
-18.2434539794922,-55.9550628662109,
-16.6140136718750,-50.9341239929199,
-3.30616259574890,-20.1990375518799,
-2.04398345947266,6.29554748535156,
-9.32323265075684,8.16344070434570,
-1.48412537574768,-0.363056659698486,
19.1636962890625,-1.10586583614349,
11.5059738159180,11.3114166259766,
-29.7941894531250,24.2068138122559,
-51.9601669311523,25.7756042480469,
-13.4975051879883,17.7272796630859,
37.0606803894043,14.9910564422607,
26.6284751892090,27.1582012176514,
-31.2069797515869,33.0465736389160,
-45.6464347839356,7.42655563354492,
15.3757972717285,-44.5152053833008,
69.3045730590820,-78.7230377197266,
47.6990890502930,-57.7701721191406,
-6.05860805511475,-1.23608338832855,
-8.36536216735840,27.6322231292725,
38.3223876953125,-0.562159836292267,
58.6372184753418,-45.7523460388184,
24.6132297515869,-58.0600051879883,
-6.53636932373047,-41.6151847839356,
8.10785770416260,-28.1477870941162,
33.4335327148438,-21.6293334960938,
28.1404285430908,2.45527124404907,
12.2063760757446,38.7542114257813,
16.7258510589600,47.6048927307129,
18.8979892730713,15.9840774536133,
-12.6241779327393,-13.1090717315674,
-48.2819671630859,0.151182889938355,
-38.2845382690430,26.5893402099609,
1.25188565254211,13.0931453704834,
8.92078495025635,-32.8711967468262,
-24.2076816558838,-53.7951126098633,
-36.8076972961426,-27.0536899566650,
5.31066322326660,-0.307599544525147,
44.8084259033203,-14.9430780410767,
19.9889602661133,-45.5934410095215,
-34.9458580017090,-50.6608963012695,
-40.0100097656250,-34.6883316040039,
8.57778453826904,-34.1531257629395,
43.0444145202637,-49.5081253051758,
25.8327560424805,-44.2188568115234,
-10.2675800323486,-5.47803401947022,
-21.2357139587402,27.2981281280518,
-16.9531364440918,22.1990623474121,
-22.7789916992188,2.76033449172974,
-31.1460819244385,4.11484861373901,
-18.2854557037354,20.2521209716797,
10.5998401641846,18.1002101898193,
21.7473468780518,-6.48296642303467,
7.93658685684204,-29.4853610992432,
-7.14409112930298,-31.2474727630615,
-13.4045209884644,-14.3079881668091,
-28.2132797241211,7.36705827713013,
-49.7237510681152,25.6832599639893,
-54.2510566711426,30.6101875305176,
-26.8977088928223,5.93121480941773,
16.8688812255859,-36.3279266357422,
48.5719337463379,-58.5862846374512,
52.3963050842285,-36.9746093750000,
31.7525863647461,6.38734006881714,
-4.20280551910400,34.7266197204590,
-37.5757217407227,39.1112899780273,
-40.1400833129883,28.3915691375732,
-5.17937231063843,5.48594236373901,
30.7213802337647,-30.8432483673096,
24.1370983123779,-58.8198242187500,
-8.66975116729736,-46.9828567504883,
-14.7727794647217,0.413511276245117,
20.3189735412598,36.4741439819336,
50.1367874145508,22.2564754486084,
36.5040512084961,-17.5590820312500,
4.89685678482056,-33.5349349975586,
-2.32344841957092,-14.4350013732910,
15.0863933563232,9.77336597442627,
17.2790889739990,18.2721939086914,
-3.92265748977661,20.5627155303955,
-8.93792629241943,24.3000984191895,
15.2232761383057,26.0492858886719,
33.2707939147949,19.3174896240234,
19.3232212066650,10.3107099533081,
1.15643763542175,6.69165515899658,
15.8701744079590,0.343733489513397,
48.9181709289551,-9.19101333618164,
55.4417304992676,-1.05325353145599,
31.1881504058838,33.5900650024414,
9.33267021179199,62.2972068786621,
0.763789713382721,45.2780456542969,
-17.3605823516846,-5.16305685043335,
-49.5229148864746,-31.9333610534668,
-55.2159461975098,-13.1778964996338,
-12.2723674774170,8.46366786956787,
36.9406089782715,-8.16145515441895,
36.4426574707031,-43.7526245117188,
-4.61294078826904,-45.5346794128418,
-26.0907039642334,-8.31912994384766,
-10.2005176544189,22.1673717498779,
0.420317351818085,15.0726871490479,
-25.2530841827393,-2.71675229072571,
-63.4009895324707,1.46266186237335,
-68.1709289550781,17.7293815612793,
-33.6461410522461,9.46185588836670,
3.68796014785767,-27.3202629089355,
17.4193897247314,-56.7609481811523,
18.2244777679443,-48.2785644531250,
19.8967819213867,-9.13525581359863,
24.9391193389893,31.7769489288330,
28.4207363128662,49.4586181640625,
19.2088260650635,43.8421058654785,
-12.5568246841431,27.5787677764893,
-53.0070114135742,11.4964370727539,
-62.9690246582031,4.91183376312256,
-20.8932266235352,13.4425334930420,
36.7811393737793,28.7523078918457,
46.4139251708984,40.1036529541016,
-3.60670924186707,33.3401145935059,
-52.0387840270996,3.02526569366455,
-40.2711334228516,-34.8691787719727,
7.38230085372925,-50.9542465209961,
18.8407764434814,-28.5514602661133,
-17.1494503021240,8.19022369384766,
-41.0448646545410,19.2483291625977,
-11.9329395294189,-5.42075109481812,
35.5969810485840,-34.8060340881348,
42.0836143493652,-25.6613388061523,
7.03710079193115,14.8557329177856,
-25.1154594421387,39.9317703247070,
-25.5998935699463,15.8016633987427,
-11.1408653259277,-33.9311676025391,
0.0979384481906891,-61.5276031494141,
14.0525159835815,-50.6991348266602,
37.8205986022949,-20.5087833404541,
56.7290115356445,6.13285541534424,
54.5703430175781,17.2465038299561,
39.0784988403320,10.5584974288940,
26.0094909667969,-16.1697311401367,
11.6283426284790,-45.8737640380859,
-5.87208843231201,-44.2102355957031,
-16.1417007446289,-2.86600351333618,
-12.1389131546021,43.8553352355957,
-12.5944604873657,55.0979843139648,
-39.2073554992676,36.2128372192383,
-72.6385192871094,21.9439601898193,
-66.8448333740234,22.3246650695801,
-11.8320178985596,8.02111434936523,
41.3881187438965,-29.1599369049072,
42.8237571716309,-51.1876029968262,
2.89699029922485,-26.2419128417969,
-26.1951675415039,26.4762897491455,
-23.8653945922852,51.5893020629883,
-18.7579002380371,33.9974327087402,
-33.4363136291504,9.24502182006836,
-50.7338523864746,6.39323711395264,
-36.0996398925781,14.3398694992065,
1.68236768245697,13.2954969406128,
21.5775814056397,8.29052829742432,
-1.44440114498138,16.4844455718994,
-39.3832511901856,32.2989959716797,
-43.3912429809570,37.4945144653320,
-6.21597576141357,29.5369663238525,
29.9483184814453,14.0946884155273,
28.5581684112549,-3.95255756378174,
-3.49633264541626,-27.9178752899170,
-29.8008117675781,-45.3108177185059,
-28.4006824493408,-39.4328804016113,
-16.0890941619873,-10.8504199981689,
-7.19897842407227,8.80270481109619,
5.26047229766846,1.29801678657532,
26.6845397949219,-12.5965566635132,
38.0069046020508,-10.0843467712402,
14.1747102737427,5.56195020675659,
-27.3735485076904,11.5292415618896,
-44.0443115234375,2.86210680007935,
-15.1379299163818,-4.99914550781250,
22.1970520019531,-6.48606109619141,
18.2468872070313,-16.3050880432129,
-26.3742618560791,-39.0009994506836,
-57.6834106445313,-57.5178184509277,
-37.0973472595215,-55.0565147399902,
17.1204299926758,-42.2798004150391,
54.6164817810059,-41.1227455139160,
52.5709457397461,-47.7368240356445,
32.2223701477051,-35.9462738037109,
15.5264873504639,1.32788550853729,
1.02131795883179,38.4458427429199,
-26.1208972930908,42.9625663757324,
-54.9776763916016,13.3745698928833,
-58.0410728454590,-23.2528266906738,
-28.5141372680664,-40.6664657592773,
9.62327575683594,-37.1782531738281,
30.2464599609375,-27.6552829742432,
31.2492485046387,-22.7304840087891,
24.3811111450195,-20.3794898986816,
11.5347595214844,-11.9584169387817,
-7.86509037017822,4.40392017364502,
-22.4753932952881,23.0518283843994,
-15.3404560089111,36.0845947265625,
-0.199921309947968,33.2251167297363,
-4.20425128936768,16.5721721649170,
-35.6856651306152,-4.73034095764160,
-61.6924591064453,-22.0581150054932,
-56.0194091796875,-25.4984283447266,
-29.1736106872559,-17.1631927490234,
-12.8386335372925,-6.84255838394165,
-11.3670635223389,4.01365041732788,
-8.35288906097412,15.8456335067749,
-4.53814935684204,30.0677604675293,
-10.4703178405762,36.6761093139648,
-23.7491226196289,19.7554912567139,
-19.0250473022461,-15.8726787567139,
16.7584972381592,-43.4920120239258,
55.3783302307129,-30.5679626464844,
64.0110549926758,18.0353984832764,
45.4593658447266,61.1825256347656,
25.5456027984619,57.9025573730469,
15.5631475448608,9.01064109802246,
15.9618892669678,-43.6325340270996,
30.4021186828613,-52.8663711547852,
59.5277938842773,-12.6775131225586,
72.3801193237305,41.7927780151367,
42.2826461791992,70.7687530517578,
-9.49397563934326,56.0772552490234,
-26.0642318725586,12.5261096954346,
10.6442003250122,-28.3682670593262,
47.2758369445801,-41.1367874145508,
31.2660446166992,-17.8645801544189,
-15.2929935455322,26.2932491302490,
-26.9657821655273,59.6572418212891,
6.31750440597534,54.8774566650391,
29.7278556823730,16.0384101867676,
6.46358394622803,-18.5922546386719,
-33.1082649230957,-15.1381731033325,
-48.6615982055664,21.4709987640381,
-38.9038467407227,47.4053802490234,
-29.3361816406250,25.1992740631104,
-20.4417552947998,-21.5244293212891,
4.44482135772705,-42.8341712951660,
33.8655395507813,-17.2187118530273,
43.7148628234863,18.2689533233643,
29.2099361419678,17.3070945739746,
17.5148792266846,-9.13848781585693,
20.4566249847412,-17.7847156524658,
13.1294021606445,7.33479976654053,
-18.6081638336182,31.4413089752197,
-47.0841674804688,19.2788143157959,
-39.8577308654785,-8.30577564239502,
-7.79814100265503,-8.80547046661377,
7.59666681289673,19.4633922576904,
-11.1065053939819,36.0272865295410,
-38.7913169860840,7.24007272720337,
-43.2038040161133,-45.1454048156738,
-19.6018104553223,-72.9859542846680,
13.8924283981323,-63.1270065307617,
39.1387863159180,-37.7834281921387,
46.3513793945313,-12.9425802230835,
29.2132072448730,14.7393188476563,
-6.30482959747314,43.8376579284668,
-33.6413421630859,49.2881202697754,
-28.0647487640381,13.6883621215820,
9.13753795623779,-30.7599563598633,
42.2452354431152,-28.8621826171875,
38.8037948608398,27.7463035583496,
5.00076007843018,74.2342376708984,
-23.2879257202148,49.5087547302246,
-17.7758598327637,-21.0259361267090,
11.7041683197021,-58.7129554748535,
33.7345924377441,-31.2183227539063,
34.0740280151367,9.56523895263672,
22.8591556549072,10.1059370040894,
10.1457433700562,-12.9601802825928,
-5.30189943313599,-16.7419166564941,
-19.5782642364502,2.73702335357666,
-15.8139438629150,9.08805084228516,
8.37248706817627,0.668533563613892,
29.3038520812988,15.0807905197144,
20.0126819610596,51.3308715820313,
-9.86615180969238,59.8904113769531,
-16.4431610107422,17.2743225097656,
10.8772430419922,-23.9255619049072,
31.9010276794434,-8.86136627197266,
8.73196029663086,40.0093040466309,
-36.7035942077637,57.9315223693848,
-49.5931892395020,37.7567558288574,
-16.5118389129639,22.9811744689941,
14.4465408325195,28.0119838714600,
2.45579433441162,14.2269115447998,
-29.1299839019775,-32.9817657470703,
-31.0911350250244,-61.3228569030762,
2.55411601066589,-27.9816188812256,
28.2315788269043,29.8058795928955,
11.3950347900391,45.4876060485840,
-32.4957809448242,17.3166007995605,
-65.1111831665039,-0.190519988536835,
-66.1867065429688,14.1046705245972,
-49.1736984252930,16.8369331359863,
-27.7425785064697,-18.1829910278320,
-3.68022322654724,-55.7666702270508,
19.6333675384522,-48.2156448364258,
32.7290954589844,-8.21979236602783,
27.8487396240234,8.32208442687988,
7.34533977508545,-20.0294017791748,
-14.6575593948364,-48.0568733215332,
-20.2273349761963,-34.0330047607422,
-8.67303562164307,8.44335746765137,
9.03756141662598,29.5666313171387,
17.6151943206787,13.2942466735840,
18.8106555938721,-11.8751039505005,
27.1122570037842,-11.1357345581055,
47.6125793457031,15.5750732421875,
57.8731803894043,31.2232055664063,
33.9838447570801,19.3500957489014,
-11.9611454010010,-0.475829273462296,
-40.1463088989258,-0.512729287147522,
-24.9380741119385,18.1897850036621,
7.65341758728027,29.4564914703369,
17.5610961914063,17.6917266845703,
-2.66996264457703,-4.64510059356689,
-19.0481300354004,-16.8851737976074,
0.200512170791626,-18.5370101928711,
40.9819068908691,-20.9041919708252,
67.8258743286133,-27.5774173736572,
60.8066558837891,-24.0089054107666,
31.4824771881104,0.529297828674316,
9.16869068145752,39.4101257324219,
7.31258296966553,68.1716918945313,
18.1500892639160,66.1382598876953,
27.1891937255859,32.0067100524902,
23.0287189483643,-8.89446544647217,
2.85313367843628,-22.7199935913086,
-20.9617958068848,-1.28233075141907,
-29.6236114501953,24.3073501586914,
-10.4156513214111,16.4541473388672,
22.5548820495605,-18.0025100708008,
34.1563224792481,-33.4873275756836,
3.25216245651245,-5.75505590438843,
-48.1284866333008,34.8222312927246,
-65.1569213867188,40.1473541259766,
-25.3034591674805,7.34114265441895,
29.7253074645996,-17.2038726806641,
42.0261840820313,-2.02197313308716,
2.11978864669800,30.7606124877930,
-43.5479965209961,38.6103401184082,
-57.0348396301270,13.6848526000977,
-39.9460563659668,-19.3364353179932,
-10.4968919754028,-32.0323371887207,
24.2505588531494,-27.6423053741455,
57.1200141906738,-25.2500114440918,
63.3523216247559,-26.9599761962891,
29.3337173461914,-27.0566768646240,
-8.05532932281494,-26.0592365264893,
0.991683006286621,-30.1789894104004,
44.4518165588379,-34.2280921936035,
60.1112518310547,-25.7056789398193,
22.2120208740234,0.665163278579712,
-23.8638000488281,19.6746406555176,
-34.2923431396484,6.29684305191040,
-27.1013679504395,-21.2033615112305,
-38.3507270812988,-20.8827037811279,
-54.0447807312012,18.4279708862305,
-37.4075851440430,50.1759643554688,
1.56790387630463,26.8158493041992,
6.33441352844238,-34.6404190063477,
-28.8592948913574,-68.7702255249023,
-41.5525054931641,-51.8789596557617,
3.01152133941650,-19.0703144073486,
60.3814773559570,-9.14443874359131,
67.7206878662109,-10.6723546981812,
37.6746788024902,10.2044515609741,
24.4850044250488,52.1257247924805,
34.1952629089356,73.8685302734375,
19.3438472747803,55.4616394042969,
-29.5108623504639,16.1222648620605,
-62.6899032592773,-19.2134323120117,
-41.5531082153320,-41.6922569274902,
0.758648276329041,-47.4481773376465,
4.32897615432739,-37.4601287841797,
-28.1649684906006,-28.7856464385986,
-37.0757865905762,-43.9597206115723,
3.78514862060547,-69.2104492187500,
50.8525352478027,-58.7513122558594,
52.9024772644043,-0.874463796615601,
14.7656917572021,49.2854881286621,
-14.3381357192993,31.8216514587402,
-2.06360816955566,-28.0955200195313,
30.8391971588135,-46.4704399108887,
39.1764450073242,0.0422739982604981,
12.0513200759888,41.8253822326660,
-19.8811378479004,19.1997795104980,
-21.5999889373779,-29.9900207519531,
6.65507745742798,-31.6920356750488,
32.7275772094727,19.1082916259766,
31.6164073944092,55.7607574462891,
9.29738616943359,35.6235847473145,
-6.40158033370972,-9.24575424194336,
2.16197276115418,-26.9140834808350,
21.8435153961182,-12.8189516067505,
29.7344951629639,6.36257648468018,
19.8663883209229,20.8412837982178,
-0.873778343200684,39.5144538879395,
-19.5656471252441,54.1674003601074,
-29.0247497558594,40.8131675720215,
-30.5745830535889,0.247854709625244,
-27.7663116455078,-38.6336174011231,
-19.1861743927002,-51.8577995300293,
-5.25826740264893,-32.7412719726563,
12.8687705993652,4.59166049957275,
27.6431102752686,37.3492927551270,
21.5900726318359,41.0492553710938,
-10.4187278747559,7.65413808822632,
-46.9444313049316,-36.7333030700684,
-49.6829071044922,-48.8453216552734,
-4.55210113525391,-12.9868755340576,
47.9268913269043,30.8529491424561,
52.5131721496582,41.4481735229492,
2.05248785018921,25.3569087982178,
-47.0730094909668,11.6746749877930,
-38.7517585754395,6.23730230331421,
16.3656997680664,-11.8642187118530,
59.1887664794922,-40.8246116638184,
58.5276947021484,-49.5283203125000,
42.1481399536133,-19.7505683898926,
43.3819198608398,23.4114780426025,
53.7673873901367,38.7715568542481,
48.0800247192383,22.8722667694092,
28.4463729858398,0.910127639770508,
15.7811412811279,-17.0848560333252,
14.3723764419556,-34.2556877136231,
4.22005891799927,-42.7776107788086,
-20.4451866149902,-21.1921176910400,
-34.9003601074219,24.2934265136719,
-29.8058185577393,51.6166687011719,
-18.9590988159180,39.8635978698731,
-16.3586006164551,7.88015985488892,
-3.51578927040100,-9.70927238464356,
33.3767738342285,-12.5606031417847,
64.1651687622070,-18.5494880676270,
52.8864593505859,-27.7153148651123,
16.9575786590576,-21.9097824096680,
-0.907938003540039,-3.02835536003113,
8.18922996520996,-0.545821905136108,
8.25546741485596,-22.7135848999023,
-18.8833255767822,-40.4622802734375,
-38.3171424865723,-33.8511581420898,
-13.8899345397949,-19.1680736541748,
30.2134685516357,-14.0388221740723,
48.1929016113281,-10.1052570343018,
38.4943962097168,12.6662950515747,
33.7970046997070,40.6227531433106,
36.5511360168457,49.2584342956543,
26.5880832672119,36.5659179687500,
5.43881559371948,31.3091373443604,
6.31349945068359,42.2663307189941,
29.0968551635742,41.2066574096680,
28.8773651123047,16.0406055450439,
-14.0126199722290,-7.96627092361450,
-54.4383125305176,-7.36023998260498,
-35.5681838989258,-0.408830255270004,
20.6168766021729,-4.93266725540161,
44.2284507751465,-4.62250232696533,
15.6674089431763,23.3650817871094,
-12.2589817047119,58.7408485412598,
-1.63274407386780,63.1756095886231,
15.3671007156372,36.1456069946289,
-2.60220098495483,24.8826389312744,
-39.1658744812012,43.4221611022949,
-57.4829521179199,46.2550621032715,
-51.3083419799805,2.19937515258789,
-42.2629089355469,-46.5415000915527,
-37.6410751342773,-44.6940460205078,
-17.8936843872070,-11.9289436340332,
16.8548831939697,-11.4059820175171,
39.7269439697266,-45.5453224182129,
37.9277534484863,-59.7550926208496,
36.7571563720703,-29.1916084289551,
52.8006744384766,4.94642496109009,
63.9991340637207,5.72574806213379,
52.8404235839844,-1.46231901645660,
32.1789283752441,24.5107593536377,
13.9265451431274,61.0256767272949,
-12.5226697921753,56.8052978515625,
-50.8934173583984,17.3091735839844,
-67.1931915283203,-8.58894443511963,
-26.4762992858887,-12.5652990341187,
41.8716430664063,-28.5566234588623,
64.1673889160156,-50.6242828369141,
28.0094928741455,-33.9346389770508,
-5.45973300933838,23.0655498504639,
13.6019620895386,54.8755836486816,
46.3890228271484,19.9972419738770,
32.8076553344727,-23.5677986145020,
-13.6604108810425,-3.48485517501831,
-29.5698776245117,58.0301513671875,
4.04143142700195,69.2016372680664,
30.0671997070313,16.5617103576660,
10.0894203186035,-17.0155487060547,
-23.0524597167969,15.4042644500732,
-14.2635622024536,60.6094322204590,
28.8143901824951,54.2416992187500,
47.1787414550781,23.2173137664795,
11.6135997772217,26.9736309051514,
-41.8313522338867,59.9651832580566,
-64.8898239135742,62.5587882995606,
-53.7229919433594,20.0587310791016,
-35.9651451110840,-19.9577903747559,
-28.2117633819580,-24.3362731933594,
-21.3890571594238,-23.0600509643555,
0.567836403846741,-44.5255317687988,
30.5366783142090,-59.8948783874512,
40.2133789062500,-29.6688022613525,
13.8051061630249,24.3697109222412,
-28.6358413696289,42.2599830627441,
-49.2949447631836,10.4035739898682,
-30.5835685729980,-27.5975151062012,
4.83387947082520,-33.0236358642578,
17.8432197570801,-14.0147771835327,
-4.71824645996094,-0.938151717185974,
-37.5735855102539,-4.59226322174072,
-49.9336128234863,-7.10700178146362,
-41.6269073486328,-1.51108276844025,
-32.7744331359863,-5.17671155929565,
-35.8058967590332,-27.8801746368408,
-41.4168968200684,-51.7504348754883,
-39.1599311828613,-50.4776573181152,
-26.1519775390625,-20.5182800292969,
-11.5788297653198,10.4661664962769,
-5.31566858291626,10.9949913024902,
-7.47182703018189,-18.9233360290527,
-14.6727647781372,-36.4453468322754,
-16.2991161346436,-12.3502569198608,
-7.48029851913452,28.1047058105469,
4.84894275665283,35.0887641906738,
6.29711389541626,-0.222852230072021,
-5.36785602569580,-33.8147315979004,
-12.8019895553589,-17.4120597839355,
2.88251781463623,29.6184806823730,
26.4357471466064,42.8389587402344,
26.1270160675049,5.15913772583008,
-6.21633625030518,-26.5026702880859,
-36.8905982971191,-2.36633825302124,
-28.1669692993164,43.3061485290527,
13.1895847320557,43.4488945007324,
42.9445915222168,-9.77575111389160,
39.6365280151367,-49.4129333496094,
29.1246986389160,-34.5329666137695,
40.1076965332031,-3.69170188903809,
63.8068771362305,-7.87942457199097,
71.6367492675781,-24.4239120483398,
52.9948577880859,-0.193556174635887,
23.9091873168945,54.5057945251465,
-6.06918525695801,67.4254608154297,
-41.5900306701660,15.6867609024048,
-69.3149948120117,-37.6368789672852,
-60.6597824096680,-32.2751884460449,
-11.6957550048828,1.97127008438110,
34.4732742309570,4.14850950241089,
35.0822181701660,-26.8882751464844,
5.92056274414063,-42.0927505493164,
0.701875865459442,-24.7290592193604,
31.9422645568848,-10.6444005966187,
50.8662719726563,-23.4794540405273,
20.5317420959473,-36.0977325439453,
-32.2783508300781,-24.6474590301514,
-48.6256904602051,-12.1926097869873,
-11.4165544509888,-16.9107780456543,
36.1410331726074,-16.5886802673340,
39.5705299377441,14.3176536560059,
0.289295911788940,53.2374382019043,
-42.7307128906250,57.5848312377930,
-53.1109199523926,35.3582611083984,
-25.8219165802002,29.3549251556397,
8.05065155029297,48.6278648376465,
21.8091640472412,54.2183570861816,
13.8819808959961,19.2779064178467,
10.8612298965454,-18.7433204650879,
25.3697509765625,-13.1517372131348,
32.7094459533691,20.1305236816406,
3.21233797073364,24.9761600494385,
-47.5581398010254,-15.9144268035889,
-66.0946731567383,-52.6960220336914,
-24.1908969879150,-39.5586585998535,
33.6234321594238,9.88431549072266,
41.3004837036133,41.6817970275879,
-2.21559762954712,24.6278152465820,
-32.9788894653320,-14.7902269363403,
-4.73174762725830,-29.8283309936523,
53.8624000549316,-3.99548673629761,
77.2956924438477,32.1776275634766,
43.2810554504395,46.8966331481934,
-6.40781974792481,36.4969100952148,
-26.4901275634766,22.5774726867676,
-18.4704971313477,19.0084724426270,
-10.4258861541748,17.0983448028564,
-13.4450025558472,-3.98293805122376,
-11.7324943542480,-33.2348022460938,
8.46687126159668,-36.2188606262207,
31.4214611053467,-0.544181108474731,
28.2126712799072,46.8234367370606,
0.540236949920654,67.0028686523438,
-29.1200981140137,48.1536598205566,
-41.2289199829102,12.0273666381836,
-37.1054687500000,-17.0339279174805,
-27.6296119689941,-36.4487075805664,
-16.8659152984619,-45.5860176086426,
-4.89188814163208,-30.3429050445557,
-1.51230251789093,8.88796806335449,
-17.3518199920654,38.9505348205566,
-36.4470596313477,24.0940132141113,
-30.4752979278564,-27.9928684234619,
1.80653238296509,-60.8551712036133,
25.2538185119629,-35.7190742492676,
10.7265090942383,18.6720886230469,
-29.0130729675293,45.8027648925781,
-52.1585121154785,32.4244079589844,
-42.8713684082031,9.70089054107666,
-25.0258922576904,10.3585920333862,
-20.9874935150147,26.4178485870361,
-20.1593341827393,31.5302371978760,
-4.58939552307129,29.7056999206543,
15.6252212524414,36.1606407165527,
12.9036417007446,46.9295043945313,
-10.1415195465088,40.7733078002930,
-20.1106376647949,9.31698703765869,
7.41457176208496,-25.9879608154297,
44.6837768554688,-34.1117973327637,
44.8781166076660,-6.98642635345459,
2.38138628005981,30.3659095764160,
-37.8173866271973,41.4902420043945,
-37.8588562011719,7.29068708419800,
-14.5090942382813,-52.0776672363281,
-11.1161823272705,-83.6189422607422,
-31.6371040344238,-52.3402481079102,
-35.6903572082520,13.7162322998047,
-2.75545382499695,48.2966499328613,
31.7466964721680,24.0828819274902,
17.9822502136230,-15.4745693206787,
-33.4750442504883,-21.0797538757324,
-62.2364234924316,-3.74097728729248,
-35.5374565124512,-10.1750354766846,
14.7652473449707,-46.3608970642090,
39.3143730163574,-59.4438629150391,
26.2817268371582,-15.6943206787109,
-2.10688853263855,45.2084503173828,
-26.1238727569580,55.5558700561523,
-39.5102005004883,12.3423833847046,
-28.3580341339111,-34.0069122314453,
9.45225906372070,-45.4101448059082,
46.5404396057129,-32.2928771972656,
44.1324005126953,-20.5299587249756,
2.99188423156738,-10.0233564376831,
-30.7910728454590,-3.95547366142273,
-20.6861457824707,-12.6447734832764,
12.7774200439453,-33.9053840637207,
30.1556568145752,-38.4741668701172,
27.0864562988281,-4.20316028594971,
25.7881164550781,47.1881179809570,
30.2390060424805,70.3855438232422,
23.5541381835938,57.2213516235352,
-3.49689388275147,42.4794349670410,
-29.2195510864258,48.6362991333008,
-32.0111732482910,55.6949424743652,
-16.3785572052002,42.1536788940430,
1.46197390556335,13.6169176101685,
13.1998062133789,-12.0575971603394,
19.3669166564941,-29.3597126007080,
13.0260210037231,-47.3681297302246,
-10.4489336013794,-57.3982276916504,
-33.0155868530273,-47.8295745849609,
-31.8593215942383,-28.4414386749268,
-9.48431396484375,-20.7410144805908,
12.9447441101074,-24.3039875030518,
21.8180656433105,-17.8506145477295,
23.9209861755371,5.42628335952759,
33.3216018676758,18.4815025329590,
48.7498474121094,-2.45587587356567,
58.5502548217773,-31.5938529968262,
51.3498497009277,-23.8098297119141,
25.2960872650147,24.5449428558350,
-16.7102718353272,58.6466178894043,
-56.7659835815430,32.4273262023926,
-65.7877502441406,-35.0960235595703,
-37.1426544189453,-70.2031250000000,
-2.77112483978272,-38.2242240905762,
2.34609436988831,17.7679748535156,
-14.4572544097900,30.8309936523438,
-20.1499729156494,0.959227442741394,
-3.80291914939880,-17.9095687866211,
11.1859941482544,8.77081203460693,
4.95794868469238,42.1512413024902,
-4.65069198608398,30.9759979248047,
5.31424283981323,-14.8217363357544,
17.2460651397705,-32.3106002807617,
0.753523468971252,6.60871505737305,
-34.1359634399414,50.4482154846191,
-42.4115524291992,39.2777519226074,
-15.9145889282227,-16.2541446685791,
5.55286788940430,-53.6985092163086,
-8.76165103912354,-37.1868400573731,
-26.4570980072022,3.19877600669861,
-6.20284175872803,10.5233411788940,
38.2450675964356,-17.8559532165527,
49.2343826293945,-45.6409606933594,
10.2998304367065,-46.5079689025879,
-28.8399734497070,-34.9846992492676,
-23.5606632232666,-28.4331512451172,
7.82521581649780,-19.8072834014893,
14.8077087402344,5.88023853302002,
-9.49267101287842,35.1791267395020,
-31.2482013702393,31.9300441741943,
-27.4462985992432,-3.95503211021423,
-12.1139583587646,-27.8874683380127,
-8.01362228393555,-6.99382400512695,
-15.6180830001831,30.8964443206787,
-26.3661823272705,32.9976043701172,
-35.7922554016113,-8.16008090972900,
-44.2248725891113,-48.3892745971680,
-43.4565048217773,-56.3717460632324,
-24.2932090759277,-52.9343261718750,
6.26289129257202,-60.9963531494141,
29.0760250091553,-67.7111587524414,
40.0450210571289,-49.6584625244141,
48.1065483093262,-10.0247964859009,
53.9152259826660,19.2264690399170,
44.8438072204590,28.5234165191650,
13.7819728851318,32.9371604919434,
-26.0197181701660,35.9536705017090,
-45.5543441772461,23.9550113677979,
-29.2983493804932,2.75356173515320,
6.08330821990967,0.568630218505859,
30.2774410247803,19.2002696990967,
24.9711227416992,24.6952781677246,
1.84193825721741,4.54135513305664,
-14.7500467300415,-5.58505582809448,
-8.43317890167236,21.0053501129150,
8.52343559265137,48.6576652526856,
8.74698638916016,23.9106273651123,
-8.63482856750488,-36.2464828491211,
-14.8639268875122,-59.7891235351563,
5.71934318542481,-18.4674720764160,
31.7840900421143,23.5243568420410,
34.2583732604981,8.90408325195313,
22.1085033416748,-32.2489242553711,
27.5561790466309,-40.7186965942383,
55.2243957519531,-13.6222782135010,
65.5267410278320,-0.622171759605408,
34.9292411804199,-14.2818889617920,
3.53426122665405,-19.5917110443115,
17.8398456573486,2.51421165466309,
50.7819671630859,23.5281867980957,
39.1874046325684,18.6283054351807,
-20.2847480773926,7.95471334457398,
-55.0243530273438,15.5817136764526,
-24.8375854492188,20.7037372589111,
17.6579704284668,-4.94101238250732,
6.39869832992554,-40.3107490539551,
-40.8721389770508,-33.4627799987793,
-51.2813339233398,14.7762832641602,
-10.2064008712769,52.9186744689941,
22.3599910736084,51.2327041625977,
9.18211174011231,30.7071266174316,
-11.4187374114990,23.5495510101318,
-3.98282575607300,28.1525363922119,
8.17277431488037,22.6273536682129,
-13.8762836456299,11.0723667144775,
-46.9275436401367,13.5457763671875,
-47.0499458312988,25.8716201782227,
-18.9309425354004,24.5348320007324,
-10.7377853393555,4.62073516845703,
-27.8027229309082,-15.0510320663452,
-26.3509902954102,-25.5227546691895,
12.8369903564453,-33.4729423522949,
46.3866004943848,-35.7858276367188,
27.9234771728516,-14.6732215881348,
-15.4794063568115,26.9406166076660,
-24.1883087158203,54.1941528320313,
10.1941585540771,37.8653831481934,
39.2401504516602,-6.87413835525513,
32.2423286437988,-35.4670715332031,
4.38291454315186,-34.4720191955566,
-17.1245117187500,-25.8105125427246,
-25.9109249114990,-32.7574501037598,
-33.0148315429688,-42.1792335510254,
-40.9778099060059,-31.6382484436035,
-42.3245658874512,-6.58277845382690,
-32.3733596801758,8.99011707305908,
-13.9021053314209,1.97192680835724,
11.4532966613770,-13.7214670181274,
37.3859024047852,-16.6000938415527,
46.7811851501465,-3.04692101478577,
38.3238029479981,11.6270322799683,
36.1684494018555,8.92625141143799,
51.5987701416016,-4.37617015838623,
60.1128768920898,-5.70011568069458,
32.0653190612793,17.5586185455322,
-20.6288528442383,52.2164916992188,
-51.0922279357910,60.7939414978027,
-37.3421440124512,22.8274459838867,
-13.9312496185303,-29.3285484313965,
-16.5472660064697,-45.3252639770508,
-32.8994293212891,-8.79817867279053,
-26.9412593841553,38.1770362854004,
-3.27288794517517,54.4988288879395,
-6.49694681167603,37.9944725036621,
-45.9637451171875,13.6277475357056,
-77.1716308593750,-7.76750469207764,
-53.9825477600098,-36.2048301696777,
2.76748085021973,-66.6212005615234,
32.9169731140137,-65.3465423583984,
11.9211063385010,-20.4157466888428,
-24.0081615447998,26.3823528289795,
-31.5820693969727,29.5157737731934,
-3.45873641967773,-8.59932327270508,
32.3379478454590,-43.4853439331055,
53.8749885559082,-43.9381027221680,
55.5960540771484,-16.3721733093262,
36.9615669250488,25.0335216522217,
4.73544788360596,64.9380569458008,
-20.6502952575684,78.4809646606445,
-14.3794345855713,42.7851867675781,
20.1111183166504,-21.5631542205811,
52.9732208251953,-49.5029182434082,
53.4229507446289,-8.41319561004639,
20.9412307739258,47.0405158996582,
-15.3894710540771,40.6715621948242,
-24.6162757873535,-24.3245754241943,
-10.1623935699463,-70.6303405761719,
9.07402038574219,-55.3769912719727,
19.4693832397461,-21.0100479125977,
23.8206729888916,-17.0540657043457,
32.7493858337402,-25.9543094635010,
41.7975578308106,-0.675774633884430,
29.5121021270752,51.6178054809570,
-5.64287042617798,66.7848739624023,
-38.1079025268555,20.3807868957520,
-36.7868804931641,-31.4942531585693,
-6.25467920303345,-29.2076244354248,
15.1952705383301,16.2112350463867,
3.87541913986206,44.5054283142090,
-17.6549816131592,28.2020931243897,
-11.3122110366821,-2.91955447196960,
25.2154178619385,-13.5264472961426,
45.3294067382813,4.85230255126953,
19.3801040649414,29.5900611877441,
-24.7290725708008,31.3904972076416,
-30.7189655303955,6.02209377288818,
13.8415479660034,-26.9271888732910,
56.5661773681641,-35.0168228149414,
46.9505691528320,-8.31381034851074,
-2.52925634384155,24.9321079254150,
-31.3253765106201,23.7177505493164,
-9.67802619934082,-7.63164329528809,
32.2266502380371,-23.8098201751709,
44.9463424682617,-4.31545305252075,
17.7831783294678,24.3493251800537,
-13.3578252792358,34.6727027893066,
-22.0304088592529,34.5695686340332,
-16.5793590545654,44.4775009155273,
-18.6150779724121,56.3473243713379,
-25.1580944061279,39.3801498413086,
-19.6992530822754,0.323315978050232,
3.77632331848145,-17.5810298919678,
22.0713996887207,-0.640633821487427,
13.7915334701538,11.7336864471436,
-6.43687152862549,-16.4276638031006,
-7.77875518798828,-58.0244331359863,
11.4546976089478,-61.5143394470215,
25.5192203521729,-25.6598110198975,
14.1950941085815,-1.33913505077362,
-9.54146575927734,-12.3206710815430,
-7.18475008010864,-30.1656455993652,
26.8576602935791,-24.6683998107910,
54.8764915466309,-6.81110906600952,
47.1084518432617,-8.86002445220947,
24.1116046905518,-30.7550716400147,
26.2224254608154,-40.3031768798828,
52.5441398620606,-26.2302379608154,
56.5599098205566,-6.47538280487061,
15.9168100357056,4.31082010269165,
-27.5825195312500,13.6097087860107,
-17.6445426940918,25.8003959655762,
28.2368717193604,36.0031929016113,
37.7637252807617,42.2537460327148,
-17.8869934082031,47.5779609680176,
-82.6526947021484,42.6665229797363,
-90.6459121704102,15.4072456359863,
-50.0587425231934,-27.0898590087891,
-16.6084442138672,-49.5495452880859,
-7.83985185623169,-31.4224510192871,
2.53514957427979,-1.51320266723633,
24.8430728912354,-1.16737627983093,
29.9140167236328,-20.3217411041260,
2.82465839385986,-14.4428739547730,
-22.1298770904541,19.4418888092041,
-9.14632987976074,34.7457618713379,
25.5827922821045,9.39639091491699,
40.6386108398438,-20.8684654235840,
25.7188396453857,-16.1646156311035,
5.13294982910156,6.83619499206543,
-8.05138778686523,8.97283458709717,
-20.2869224548340,-9.37124633789063,
-25.6609058380127,-9.63732624053955,
-4.71474599838257,13.9349803924561,
33.0699844360352,24.7370491027832,
50.4544715881348,9.05554866790772,
26.8660907745361,-1.48320114612579,
-3.82230854034424,14.9900093078613,
3.48842000961304,26.0159835815430,
42.2371101379395,2.54476356506348,
64.0964431762695,-29.8474922180176,
42.6830062866211,-27.3342056274414,
10.1569719314575,1.14216756820679,
3.09511470794678,12.7981863021851,
16.7936096191406,-1.69321072101593,
21.6124286651611,-3.88324117660522,
2.32316112518311,20.2528476715088,
-23.4842796325684,31.0211830139160,
-29.9271907806397,-4.96276760101318,
-11.0163393020630,-52.5028190612793,
18.4047775268555,-60.2234992980957,
36.2185630798340,-33.1114692687988,
32.4996643066406,-12.2722978591919,
16.1110286712647,-6.78498077392578,
-0.680780529975891,7.21824121475220,
-9.51461696624756,33.4631652832031,
-19.9069290161133,43.3181457519531,
-39.6243972778320,26.5488071441650,
-54.4945793151856,12.4978561401367,
-41.8013381958008,26.9092674255371,
-3.44736576080322,49.8756027221680,
33.4329910278320,49.3104934692383,
40.4254302978516,36.7820663452148,
20.9023113250732,40.7633323669434,
-0.493675291538239,51.6702995300293,
-8.79212856292725,37.5449409484863,
-6.04893875122070,2.61026525497437,
2.86830615997314,-15.7201375961304,
19.0596656799316,-5.56139469146729,
40.3298797607422,7.92286348342896,
53.3109321594238,4.00555133819580,
47.3616523742676,1.57837772369385,
32.7799606323242,18.4414958953857,
29.6726551055908,28.1031780242920,
39.1119346618652,2.39268445968628,
45.4759864807129,-33.1000251770020,
29.2694492340088,-27.8698596954346,
-3.58052730560303,17.6649627685547,
-31.6829681396484,42.7421760559082,
-32.1786155700684,16.2026271820068,
-3.60106539726257,-20.3756008148193,
30.0480976104736,-17.5131187438965,
40.4538040161133,11.6404676437378,
16.3552989959717,16.7763404846191,
-18.7379302978516,-13.0043897628784,
-31.3012580871582,-30.6264076232910,
-18.1658515930176,0.269558429718018,
-14.0475730895996,46.0497550964356,
-40.5023612976074,49.8551979064941,
-68.1014328002930,2.33332681655884,
-58.1238517761231,-47.0296859741211,
-10.3438529968262,-47.5815010070801,
33.4348793029785,-1.78966283798218,
40.2117576599121,50.7997207641602,
23.1509399414063,74.1361541748047,
8.36081600189209,60.8066787719727,
-5.70318698883057,33.1522102355957,
-25.4278736114502,13.0462102890015,
-31.2583179473877,7.03096103668213,
-9.95587825775147,9.60493755340576,
9.29521751403809,6.65396547317505,
-11.1610469818115,-13.5906152725220,
-50.5365028381348,-43.1058044433594,
-47.2247581481934,-59.5815582275391,
7.17397975921631,-45.4212074279785,
44.3803215026856,-6.97963857650757,
12.6185274124146,25.6092205047607,
-36.7999916076660,21.3348197937012,
-25.5837116241455,-16.9580669403076,
39.9822502136231,-45.8996200561523,
71.0869979858398,-30.4917449951172,
33.0167694091797,19.3621253967285,
-9.84865570068359,54.2737846374512,
-3.36840915679932,39.8536949157715,
17.9922447204590,-0.946288347244263,
1.59985470771790,-17.5154151916504,
-35.1290397644043,6.03046798706055,
-36.3889236450195,32.7887992858887,
-0.130295991897583,30.7143440246582,
20.3929157257080,12.9411706924438,
0.516123771667481,6.78461790084839,
-25.1671066284180,3.44883823394775,
-30.1443214416504,-18.7390727996826,
-35.0984878540039,-52.1444587707520,
-49.4265441894531,-60.8573379516602,
-35.0820541381836,-37.8918685913086,
22.0199394226074,-23.6168861389160,
68.7966690063477,-39.4844207763672,
60.3557968139648,-46.3943824768066,
29.3089656829834,-3.84530973434448,
31.9712123870850,55.6647529602051,
54.1748390197754,64.5329513549805,
33.8887977600098,14.3040571212769,
-30.2689323425293,-27.0550231933594,
-57.1320800781250,-16.3744087219238,
-4.53900814056397,8.94308185577393,
54.6545867919922,1.99396276473999,
41.9449005126953,-24.5719871520996,
-12.6387968063355,-21.8930969238281,
-20.0828704833984,13.1775245666504,
27.9628658294678,34.4521331787109,
52.1277809143066,20.4860382080078,
6.47948551177979,-3.35598897933960,
-54.0297775268555,-10.3205614089966,
-60.3302993774414,-15.1097469329834,
-19.1554260253906,-34.7354164123535,
17.3409729003906,-51.4905586242676,
25.8786334991455,-43.0379142761231,
31.8340320587158,-21.3984203338623,
42.5598831176758,-8.58943748474121,
33.4175758361816,-2.39760184288025,
-6.95173645019531,13.1157112121582,
-46.1043395996094,33.8633155822754,
-55.0995597839356,34.3590087890625,
-35.1282386779785,10.2137870788574,
-9.07620620727539,-15.7035980224609,
4.16115283966064,-24.5862655639648,
5.31872367858887,-21.8483047485352,
5.00244998931885,-13.5459899902344,
13.2780838012695,13.0482254028320,
27.4231052398682,52.5495643615723,
29.9743652343750,71.4897842407227,
5.80162286758423,45.3613548278809,
-35.5427436828613,1.07701563835144,
-55.4771270751953,-9.48369693756104,
-29.8189449310303,22.9542884826660,
13.2500677108765,55.8700637817383,
21.7392654418945,45.2439117431641,
-15.2076988220215,0.649135768413544,
-54.9287910461426,-36.6791915893555,
-56.7412071228027,-41.9523506164551,
-19.3767166137695,-22.6964206695557,
21.4068641662598,2.58839225769043,
35.7384719848633,27.0682945251465,
18.9218044281006,42.6851615905762,
-14.7869272232056,44.7218170166016,
-38.9884223937988,34.5404357910156,
-29.4842491149902,20.5942420959473,
14.1055908203125,8.48127174377441,
52.6277084350586,-3.18598818778992,
47.8808593750000,-13.7313776016235,
12.9924278259277,-18.3101768493652,
1.63795399665833,-10.8894214630127,
31.3401870727539,4.58415603637695,
54.8250160217285,16.7424602508545,
26.6667537689209,19.3074626922607,
-29.0868721008301,11.6526069641113,
-50.2725486755371,-12.8547410964966,
-21.0471115112305,-49.1416244506836,
12.1634225845337,-71.5190353393555,
13.5217018127441,-54.4993324279785,
6.22287368774414,-9.88680076599121,
17.7716693878174,18.3213691711426,
30.0907955169678,5.16369819641113,
16.1776504516602,-30.2941551208496,
-6.67344379425049,-45.4105606079102,
5.20734500885010,-32.5438919067383,
44.4598426818848,-13.0280923843384,
59.8128929138184,1.34209918975830,
29.8648033142090,16.3105621337891,
-8.73240566253662,29.7497329711914,
-15.1543827056885,24.1612586975098,
-1.73352193832397,-2.17965984344482,
1.62241661548615,-18.5609092712402,
-1.84710216522217,-6.76510000228882,
10.3432283401489,9.48938369750977,
30.4725494384766,-0.883347511291504,
26.0831737518311,-26.8680019378662,
-4.85044240951538,-23.6974220275879,
-28.3654460906982,20.9001350402832,
-27.5682678222656,63.0459671020508,
-28.2926082611084,56.9315986633301,
-49.5343246459961,12.8019638061523,
-70.9526138305664,-23.8281040191650,
-59.3883018493652,-29.7532672882080,
-23.4950141906738,-20.6061553955078,
-4.82707166671753,-21.9758415222168,
-22.2814617156982,-35.6024093627930,
-41.0056457519531,-47.0314331054688,
-23.8717269897461,-45.9845504760742,
18.9809894561768,-27.3246459960938,
41.2874565124512,3.12571740150452,
18.8320655822754,37.6999549865723,
-25.7282238006592,60.1937484741211,
-46.8308410644531,57.1558609008789,
-25.2401657104492,31.1034049987793,
15.4204578399658,6.57858133316040,
37.2850112915039,4.61299467086792,
32.3610877990723,21.1612396240234,
16.0538349151611,34.3405609130859,
9.47646999359131,20.7856693267822,
11.0898046493530,-10.1276245117188,
12.6181917190552,-27.8412837982178,
9.27480316162109,-19.6017208099365,
7.12117576599121,-3.12948441505432,
6.63921213150024,-8.36835765838623,
0.276487290859222,-37.7751922607422,
-18.7354850769043,-63.4666786193848,
-37.5046844482422,-61.6448173522949,
-42.7498130798340,-39.4228096008301,
-31.9457435607910,-23.0385951995850,
-19.5010509490967,-24.0253849029541,
-21.2198963165283,-27.0922012329102,
-38.7144355773926,-10.3903341293335,
-55.4089279174805,22.4699840545654,
-58.6966934204102,44.6981086730957,
-42.8695793151856,36.1426048278809,
-15.2381753921509,3.63770127296448,
9.52516365051270,-25.4840736389160,
16.2962322235107,-30.7706375122070,
-0.888705849647522,-19.8792552947998,
-30.1260051727295,-13.0535049438477,
-42.6563148498535,-24.7773303985596,
-18.8651733398438,-49.5795516967773,
28.5624980926514,-66.1355438232422,
61.2243843078613,-60.0536537170410,
55.4909744262695,-34.4710235595703,
27.5670623779297,-8.14865112304688,
15.4226331710815,2.18015170097351,
34.7193679809570,0.330230742692947,
59.2056427001953,2.48159861564636,
53.3144836425781,10.8014736175537,
16.2407608032227,10.6333494186401,
-20.6609649658203,-12.6081075668335,
-28.4061393737793,-49.0830993652344,
-9.29845428466797,-64.6148529052734,
9.41069793701172,-41.0463485717773,
9.05144786834717,4.39346694946289,
-1.64644908905029,38.6295089721680,
-5.08336734771729,39.9460220336914,
-0.604942142963409,11.2816390991211,
-3.22973155975342,-28.3583602905273,
-19.4636859893799,-55.6832923889160,
-36.3619918823242,-58.6604270935059,
-33.3940658569336,-38.2888641357422,
-13.5151500701904,-21.4501285552979,
-4.17503404617310,-27.0584754943848,
-12.9199094772339,-46.9917793273926,
-11.2352542877197,-49.6725463867188,
24.3807029724121,-19.0507087707520,
65.4080123901367,18.3715991973877,
59.9702529907227,26.2124824523926,
3.36908602714539,4.29881906509399,
-40.1404457092285,-10.5013790130615,
-18.9856109619141,2.50294494628906,
36.0100479125977,26.2686443328857,
53.8210411071777,26.4190826416016,
20.8358192443848,-0.941789448261261,
-4.09912872314453,-24.0272979736328,
15.3229799270630,-15.7687625885010,
46.5181465148926,17.5993556976318,
43.0128173828125,51.0253067016602,
14.1248731613159,57.5798339843750,
2.95909547805786,33.7326583862305,
10.8375482559204,-5.55068683624268,
1.54822874069214,-34.8796844482422,
-30.4901103973389,-35.3818550109863,
-46.5032730102539,-12.6464214324951,
-25.3484897613525,5.87999010086060,
5.31867456436157,4.35566234588623,
6.79882240295410,-13.2535381317139,
-4.19702243804932,-28.0147800445557,
14.8346261978149,-27.4476127624512,
57.2928314208984,-15.8445520401001,
75.1608886718750,-0.474827170372009,
47.0276069641113,18.1594276428223,
2.29823517799377,38.9245491027832,
-15.4117507934570,52.5135383605957,
-0.843368768692017,48.1631546020508,
16.0787792205811,22.6135520935059,
8.08308410644531,-15.4433212280273,
-17.4263916015625,-38.6607246398926,
-35.4132423400879,-24.7132453918457,
-22.9649353027344,23.6328353881836,
20.0609607696533,69.3873519897461,
59.2208023071289,70.9755706787109,
50.0051612854004,26.7031936645508,
-4.02247381210327,-20.2507667541504,
-48.2305870056152,-33.6593513488770,
-37.3945846557617,-18.6372680664063,
9.21277046203613,-11.2142448425293,
32.3416633605957,-19.2089061737061,
15.5645446777344,-18.6147918701172,
-7.84909296035767,3.42219567298889,
-4.57291984558106,21.7711162567139,
5.81601524353027,6.75831270217896,
-10.1187152862549,-27.6640586853027,
-37.6730728149414,-42.4572448730469,
-32.3093566894531,-21.1476879119873,
6.17187118530273,10.2890243530273,
32.0951499938965,18.2294425964355,
14.3540744781494,1.98254001140594,
-24.5700321197510,-23.8267860412598,
-37.7729454040527,-45.6752967834473,
-16.4749355316162,-62.9165000915527,
16.2773094177246,-63.3952560424805,
42.5632057189941,-40.4680213928223,
54.0365562438965,-9.07289505004883,
48.6541213989258,8.88733673095703,
25.6900024414063,6.87408924102783,
5.21131038665772,1.68168103694916,
12.7919759750366,0.430239260196686,
36.4152526855469,-0.0658308863639832,
32.4159126281738,-0.475179910659790,
-15.9276371002197,7.52769708633423,
-66.1859054565430,26.7382431030273,
-63.2986755371094,39.3714675903320,
-12.6596174240112,31.7303009033203,
34.3768424987793,21.8582248687744,
36.0309181213379,32.1788406372070,
0.909386873245239,56.4338912963867,
-32.4769287109375,63.9584388732910,
-48.8429679870606,36.2729721069336,
-52.5482254028320,-4.85535526275635,
-46.9222640991211,-39.6692237854004,
-30.8788299560547,-62.3790245056152,
-4.82746887207031,-72.2316131591797,
15.5473670959473,-57.2498359680176,
17.8648681640625,-12.3739280700684,
0.861386895179749,37.2466888427734,
-19.9334926605225,49.6803970336914,
-21.1708412170410,15.1996841430664,
10.3807449340820,-23.8144207000732,
54.9247703552246,-24.6741905212402,
72.1645736694336,14.8738861083984,
42.2414970397949,53.1857147216797,
-17.3121891021729,48.4570732116699,
-57.1676406860352,-0.256657421588898,
-50.9548645019531,-55.9125900268555,
-17.6682376861572,-73.8273620605469,
12.0307369232178,-43.2815971374512,
24.1484127044678,2.06127905845642,
26.4741020202637,14.7996053695679,
19.8939323425293,-15.9958734512329,
5.62392807006836,-44.3785018920898,
-9.43700695037842,-27.6313190460205,
-13.7232084274292,26.3103866577148,
-11.4514331817627,54.0022697448731,
-16.4650287628174,13.7236728668213,
-27.3356475830078,-53.3395957946777,
-19.8737277984619,-74.1442413330078,
18.1598701477051,-22.4921588897705,
57.3339385986328,49.5936508178711,
59.9752235412598,70.8070373535156,
26.6322002410889,29.0784339904785,
-5.90073060989380,-19.6248493194580,
-16.6954040527344,-28.1598739624023,
-19.0893630981445,-2.44710135459900,
-26.6789188385010,9.07274055480957,
-35.9389457702637,-17.7169952392578,
-36.9156875610352,-57.6978263854981,
-36.5861663818359,-61.0091323852539,
-41.8874282836914,-15.3049459457397,
-40.8892745971680,34.6938400268555,
-21.0290527343750,31.6609382629395,
-1.21839153766632,-21.7063045501709,
-10.2684478759766,-60.1061477661133,
-35.4987106323242,-40.8492202758789,
-34.8970489501953,6.69456958770752,
4.09833288192749,19.0429039001465,
41.2292976379395,-18.2475376129150,
44.7308464050293,-50.8321800231934,
36.4684181213379,-34.9998092651367,
48.5115890502930,-2.70942020416260,
66.9631271362305,-3.52472257614136,
50.2243270874023,-33.5727081298828,
1.54733443260193,-48.0315093994141,
-25.8666744232178,-30.2502746582031,
-3.05327963829041,-8.48742866516113,
29.6204357147217,-4.28509950637817,
25.6196403503418,5.41790199279785,
-5.75383186340332,33.2265205383301,
-17.3528060913086,51.6255760192871,
3.32622814178467,31.0417919158936,
22.2242145538330,-7.88760185241699,
17.9810352325439,-20.2696285247803,
6.87375020980835,-3.82825684547424,
9.26559352874756,-0.366371780633926,
22.2790756225586,-25.4056701660156,
24.0415725708008,-39.5234718322754,
12.2588071823120,-13.7750444412231,
5.91982650756836,24.4943962097168,
11.8861722946167,32.8193054199219,
14.3942852020264,7.58208131790161,
6.28415107727051,-21.3043918609619,
-6.53493928909302,-33.8599777221680,
-11.7358474731445,-40.9505805969238,
4.15283775329590,-47.7512130737305,
41.5647850036621,-43.0130653381348,
70.2665710449219,-26.2494869232178,
57.1450500488281,-16.7203273773193,
5.66422128677368,-25.4762611389160,
-30.3242721557617,-32.5135192871094,
-3.92668294906616,-27.7648372650147,
58.8161582946777,-26.5301780700684,
76.5532989501953,-35.9393730163574,
23.3098983764648,-37.2441101074219,
-32.0247879028320,-12.1831607818604,
-14.8839778900146,16.5630588531494,
44.4813995361328,14.2521152496338,
55.4738769531250,-16.0494232177734,
1.70603096485138,-31.5006904602051,
-37.8781661987305,-14.9149532318115,
-4.46703815460205,0.633270978927612,
58.4619865417481,-4.08795881271362,
72.5192337036133,-3.41258001327515,
33.8333663940430,27.3157958984375,
9.71051502227783,60.6643943786621,
27.5839614868164,55.1799163818359,
49.6548728942871,21.9528827667236,
34.9543838500977,11.4880104064941,
-1.08629071712494,35.8302192687988,
-26.8181571960449,52.7898216247559,
-37.5636100769043,32.3243026733398,
-36.9884071350098,6.56455183029175,
-15.2372016906738,11.8285617828369,
19.6105060577393,30.0342369079590,
33.1637382507324,13.7396106719971,
10.7269096374512,-30.9479751586914,
-16.7085094451904,-49.8169937133789,
-7.06601333618164,-15.1984481811523,
32.8545036315918,36.5730056762695,
51.8724594116211,56.4884757995606,
33.9642028808594,40.2271118164063,
16.2403640747070,13.0092535018921,
10.1558599472046,-9.61831188201904,
-9.98262023925781,-25.9273757934570,
-46.4420394897461,-35.2698860168457,
-50.6725158691406,-24.9144401550293,
-0.346371173858643,1.02379536628723,
49.8794174194336,19.8541564941406,
35.6054077148438,21.1642341613770,
-20.3148040771484,18.8349380493164,
-33.5695152282715,24.4881858825684,
9.75975799560547,34.2997817993164,
30.7825012207031,41.1088600158691,
-18.4638366699219,38.9937515258789,
-77.1483993530273,16.9178142547607,
-57.5120353698731,-19.3791294097900,
23.7022476196289,-41.3979377746582,
67.1626586914063,-21.9958572387695,
34.0332756042481,30.1937007904053,
-18.3141746520996,61.6640853881836,
-25.6940116882324,39.6145095825195,
3.11030244827271,2.19985961914063,
18.6802711486816,4.19947052001953,
11.0300712585449,37.4804573059082,
7.98805332183838,43.4206924438477,
23.2485923767090,13.2492446899414,
31.8169116973877,-0.629247188568115,
11.6535120010376,26.4811420440674,
-24.4992218017578,45.7782630920410,
-48.7067070007324,7.53490304946899,
-46.2948112487793,-45.2099418640137,
-15.7059535980225,-32.3967132568359,
28.4297027587891,34.8385772705078,
48.7769470214844,62.7049140930176,
25.2500152587891,7.79559707641602,
-22.1737785339355,-59.8186264038086,
-51.0920295715332,-59.0255661010742,
-35.0900421142578,-11.5627336502075,
2.44538521766663,4.76974344253540,
23.8255138397217,-15.1785640716553,
23.3756027221680,-13.5584964752197,
21.7209262847900,27.5200576782227,
22.9056415557861,52.5451545715332,
18.0508823394775,16.7125091552734,
9.95330429077148,-44.9658622741699,
12.3813934326172,-63.4563407897949,
18.5383968353272,-27.2198734283447,
1.26601159572601,20.1208209991455,
-40.0509262084961,40.6075019836426,
-62.1196327209473,32.4465065002441,
-29.2402935028076,9.43617057800293,
29.8902740478516,-13.0093460083008,
56.2314224243164,-10.1162424087524,
34.1979217529297,19.9566097259522,
9.37992477416992,42.6995353698731,
22.4943809509277,26.3548393249512,
50.8136825561523,-9.28494262695313,
48.7774314880371,-11.7603158950806,
11.9263534545898,31.2097225189209,
-18.2809638977051,66.7538833618164,
-12.3358602523804,42.8979797363281,
15.2738790512085,-17.7087020874023,
35.3619766235352,-46.2269096374512,
37.6895599365234,-22.3867397308350,
35.8723602294922,15.5966358184814,
33.5488510131836,33.4095802307129,
24.7033157348633,34.6270713806152,
5.92962741851807,35.8641395568848,
-8.47526454925537,35.4397315979004,
-6.54582643508911,30.8758258819580,
2.46521639823914,32.2299766540527,
0.610558152198792,41.3502464294434,
-20.3337192535400,39.6744117736816,
-42.3579444885254,17.3522720336914,
-43.0016441345215,-5.22690534591675,
-17.5002708435059,2.88842248916626,
11.2999057769775,29.9519691467285,
18.3245449066162,31.3347606658936,
-0.379681587219238,-5.93991947174072,
-31.0376815795898,-43.7944908142090,
-53.7845115661621,-48.4778251647949,
-53.7378196716309,-29.8822555541992,
-33.1242141723633,-12.7412261962891,
-3.52708935737610,-2.90820980072022,
17.2510166168213,6.37460041046143,
20.1014385223389,8.51853752136231,
10.7977190017700,-3.74532079696655,
7.96742868423462,-15.5967597961426,
16.2452754974365,0.736734688282013,
24.2256717681885,37.1044883728027,
18.1961650848389,50.6536941528320,
5.65448856353760,26.5314083099365,
6.38122415542603,2.17768812179565,
29.2607822418213,10.2482528686523,
50.6316795349121,33.0987319946289,
42.0327758789063,37.4067382812500,
0.195681095123291,24.3639965057373,
-39.8286094665527,16.2875442504883,
-45.4174766540527,12.3302106857300,
-24.3240890502930,-6.22498369216919,
-12.4519882202148,-30.8418483734131,
-25.3493957519531,-22.9400558471680,
-47.9740905761719,17.8587722778320,
-54.3996963500977,35.5430259704590,
-45.0670356750488,-9.19063663482666,
-32.6082763671875,-67.9219512939453,
-21.6172733306885,-68.6641616821289,
-9.18139457702637,-17.3773841857910,
-8.59766960144043,12.5200576782227,
-28.6573104858398,-14.7009124755859,
-46.1320953369141,-57.1384582519531,
-23.4352703094482,-61.2416648864746,
32.9321327209473,-32.6712722778320,
64.4665756225586,-12.2230262756348,
30.4725399017334,-10.8517036437988,
-28.9395675659180,-8.98542976379395,
-42.8576469421387,-2.42959642410278,
0.578058362007141,-3.53822755813599,
46.0059700012207,-1.82303309440613,
46.6839332580566,22.5191268920898,
22.2847099304199,53.9131202697754,
17.8936462402344,52.4629135131836,
35.8495101928711,11.8188505172730,
42.1578216552734,-23.6736526489258,
21.3621063232422,-20.9381008148193,
-5.72083663940430,-1.00750839710236,
-13.4313049316406,-1.06299185752869,
1.02596807479858,-17.0693626403809,
22.7981605529785,-13.9367561340332,
34.7297019958496,11.8786668777466,
24.0947875976563,25.0789527893066,
-4.60419416427612,17.0176925659180,
-25.6097908020020,16.9158020019531,
-21.7479610443115,42.1615104675293,
2.40007495880127,59.1257133483887,
19.4864253997803,31.3782978057861,
16.4361667633057,-24.1845912933350,
13.4630746841431,-54.3025398254395,
29.0367927551270,-32.6462287902832,
45.5274810791016,12.5667076110840,
39.0290260314941,42.0146369934082,
22.3116950988770,48.9038734436035,
16.9644374847412,46.9105644226074,
21.3405818939209,40.3555145263672,
16.3275852203369,21.2685642242432,
2.15449857711792,-7.96472549438477,
-3.17089748382568,-29.6403255462647,
-0.774357795715332,-32.9009513854981,
-19.3732414245605,-20.7392311096191,
-60.5486946105957,0.381910443305969,
-77.0968704223633,18.5627193450928,
-38.9162902832031,24.9331283569336,
9.39001560211182,10.2384014129639,
5.76117706298828,-23.2306575775147,
-29.4630489349365,-56.1823616027832,
-22.3913040161133,-61.7905654907227,
35.8482475280762,-32.6102561950684,
69.2823257446289,13.2899599075317,
31.1653404235840,45.3151741027832,
-22.2858810424805,38.7579193115234,
-11.8725366592407,-0.139070987701416,
39.7217445373535,-33.9354896545410,
44.1758041381836,-25.8328075408936,
-16.2593650817871,14.0882968902588,
-64.1483078002930,34.5270614624023,
-45.7350730895996,2.36907243728638,
-3.88279104232788,-52.1200065612793,
3.41590309143066,-66.6245193481445,
-11.1073226928711,-25.0204467773438,
1.24296092987061,24.4896621704102,
26.8915901184082,32.6601181030273,
17.4266700744629,14.3101511001587,
-26.7320098876953,10.5929279327393,
-47.7693138122559,24.3888568878174,
-15.1117420196533,21.3288269042969,
27.8966159820557,-10.1858768463135,
26.3406085968018,-36.8950195312500,
-7.71643400192261,-33.6697731018066,
-27.6685523986816,-13.4392337799072,
-19.3736495971680,1.37684810161591,
-9.30788516998291,10.6168298721313,
-9.57120132446289,20.4295158386230,
-3.86448860168457,19.0125160217285,
14.3411350250244,-2.57637023925781,
33.5874443054199,-18.5992336273193,
37.8871307373047,6.07824468612671,
31.5965538024902,59.0847396850586,
23.2120857238770,84.9075698852539,
10.1906156539917,58.8997230529785,
-16.1484470367432,11.4774074554443,
-42.8391990661621,-25.2235050201416,
-43.6645317077637,-51.1984252929688,
-9.53890419006348,-72.0089721679688,
35.3608627319336,-68.9234390258789,
58.5127563476563,-26.2678680419922,
41.9371948242188,27.1161518096924,
-4.90037965774536,37.7855758666992,
-47.8276977539063,1.69210445880890,
-60.7994575500488,-34.9572944641113,
-45.6521759033203,-40.5689239501953,
-22.9620475769043,-35.1572990417481,
-8.48773288726807,-41.3206138610840,
1.86949610710144,-44.5461997985840,
19.9807376861572,-24.8172702789307,
41.3730430603027,-0.614629507064819,
49.0617599487305,-2.01906132698059,
42.6512451171875,-21.7820014953613,
39.9440383911133,-23.6727485656738,
52.9882392883301,1.97888755798340,
58.0878334045410,19.4561538696289,
28.1988735198975,6.19123458862305,
-27.3863525390625,-20.8988018035889,
-60.0157890319824,-28.0006484985352,
-31.9089679718018,-22.5908851623535,
26.4698257446289,-31.4099369049072,
52.9558105468750,-51.0273590087891,
21.4886569976807,-50.1866912841797,
-30.6799869537354,-18.0954265594482,
-46.0447998046875,20.6170120239258,
-15.4712009429932,37.2376480102539,
19.7098808288574,35.5782318115234,
21.5190677642822,37.6998405456543,
-1.85890102386475,52.0901947021484,
-20.2007560729980,60.2043113708496,
-24.9581565856934,45.0171585083008,
-30.0401916503906,7.32331943511963,
-37.8802032470703,-31.9345684051514,
-27.3747539520264,-53.8742103576660,
13.2959976196289,-50.1734580993652,
54.5291481018066,-32.5142364501953,
58.4884796142578,-17.9681110382080,
32.9952507019043,-14.4470891952515,
16.5372028350830,-11.6503181457520,
24.1129322052002,2.69666647911072,
24.0536689758301,24.1591739654541,
-9.53016567230225,39.1647949218750,
-50.9903030395508,33.4856376647949,
-50.2946777343750,15.0039873123169,
-6.23591947555542,3.77315282821655,
34.7290992736816,10.8999118804932,
39.4177284240723,31.1949939727783,
24.3910465240479,42.5436248779297,
20.7338237762451,37.4035224914551,
31.4265861511230,23.6710796356201,
33.4468955993652,22.0159511566162,
18.7021064758301,36.3156623840332,
-0.237421408295631,55.9396171569824,
-14.6730165481567,58.7220687866211,
-30.5089874267578,40.9307174682617,
-46.9670562744141,8.97593784332275,
-55.4003181457520,-26.6848983764648,
-46.1905593872070,-54.9512901306152,
-30.6809501647949,-61.2297859191895,
-24.0248241424561,-39.9267349243164,
-25.1074295043945,-6.06602382659912,
-21.2068214416504,11.8429784774780,
-5.93314886093140,-5.96838331222534,
11.3799276351929,-42.1353263854981,
21.0499877929688,-58.0670585632324,
25.7647151947022,-36.9565238952637,
31.0849113464355,-10.0466871261597,
29.9837875366211,-16.0041828155518,
8.58351516723633,-54.2015914916992,
-20.4377441406250,-79.4254989624023,
-19.9976463317871,-53.4785957336426,
22.3212833404541,-4.30459499359131,
63.6043472290039,12.4969263076782,
53.5352859497070,-16.6684570312500,
-0.846760749816895,-44.7653312683106,
-32.1834220886231,-28.7502841949463,
-3.13931512832642,9.53846645355225,
41.9720230102539,28.1435089111328,
41.0644798278809,20.1562232971191,
5.80662775039673,13.0579195022583,
-3.59072327613831,14.1809015274048,
26.5212249755859,-0.292868375778198,
40.6014633178711,-35.0291938781738,
7.67737483978272,-44.0926094055176,
-26.3316173553467,-2.58606457710266,
-9.28048419952393,54.4870376586914,
32.6882896423340,70.1291809082031,
30.5014915466309,36.9128036499023,
-19.0771694183350,-1.26614570617676,
-47.4836273193359,-20.9048557281494,
-12.1274719238281,-34.2757263183594,
45.1318893432617,-45.1002502441406,
57.0316276550293,-32.9395866394043,
23.6791782379150,-0.530146837234497,
-4.97970771789551,15.7712574005127,
-6.43742942810059,-9.12139320373535,
3.35548424720764,-40.2242736816406,
10.5263986587524,-22.1514472961426,
18.7015419006348,41.4398422241211,
29.9752159118652,87.3283615112305,
31.6034049987793,75.9750442504883,
20.8967533111572,32.8672142028809,
6.58818149566650,-0.295692145824432,
-3.54405927658081,-10.2849655151367,
-15.7486810684204,-6.57366418838501,
-30.2170162200928,3.59944272041321,
-24.6893234252930,7.55206871032715,
5.85273838043213,-6.41647005081177,
26.1447448730469,-36.0998229980469,
6.28284168243408,-50.3691978454590,
-32.9657897949219,-33.0682373046875,
-51.3792228698731,-6.78046131134033,
-37.7570991516113,-4.71532487869263,
-23.1517353057861,-17.5737876892090,
-28.8186225891113,-4.72693443298340,
-38.6314811706543,31.3844757080078,
-37.4695777893066,37.8388099670410,
-34.3832740783691,-7.61256742477417,
-42.0252037048340,-56.0563468933106,
-41.3775939941406,-59.8136749267578,
-7.67418956756592,-30.2144088745117,
37.5381088256836,-20.8395137786865,
47.7004737854004,-42.4246864318848,
13.7995738983154,-58.5519714355469,
-17.5376262664795,-47.5770912170410,
-6.24090623855591,-30.9320240020752,
31.4793014526367,-21.0944309234619,
52.1479034423828,-0.712858915328980,
33.7859687805176,38.1893959045410,
-3.32338523864746,55.7820281982422,
-23.3079032897949,23.6570396423340,
-12.0923204421997,-25.1720123291016,
25.1700763702393,-36.5680656433106,
65.0776977539063,-11.0917959213257,
76.6501846313477,1.06464481353760,
46.5811576843262,-22.6278495788574,
1.32053494453430,-46.2750740051270,
-22.3376007080078,-36.6170310974121,
-16.5478992462158,-13.4370851516724,
-6.58953332901001,-14.3112211227417,
-5.14672565460205,-34.6367950439453,
5.70150184631348,-41.1741638183594,
36.3315467834473,-28.6211795806885,
58.0679893493652,-21.7744216918945,
37.4836158752441,-30.1779022216797,
-13.1923961639404,-29.1225128173828,
-38.8348045349121,-2.21229624748230,
-13.9283885955811,27.5350532531738,
26.7331924438477,34.2578010559082,
36.7164878845215,26.5004253387451,
14.7069282531738,33.7642478942871,
-4.00139904022217,58.8502578735352,
1.84613335132599,64.4163742065430,
10.8405942916870,24.9353713989258,
2.63898444175720,-31.5320072174072,
-15.4607505798340,-54.1603431701660,
-19.5392513275147,-30.6992912292480,
0.0301110744476318,8.48824596405029,
26.2327899932861,22.8017673492432,
38.0104141235352,7.94385766983032,
30.0357685089111,-2.91729736328125,
13.0204401016235,7.82607984542847,
-4.28674030303955,22.6671028137207,
-11.9237899780273,9.27323818206787,
-7.56458139419556,-23.1692237854004,
3.80824446678162,-30.8384876251221,
9.70078754425049,10.2019367218018,
-1.12799596786499,66.2519226074219,
-23.0483913421631,71.0612182617188,
-32.6882896423340,12.4337272644043,
-15.8304615020752,-45.8574142456055,
15.9263944625855,-32.9055099487305,
34.0777359008789,33.6440277099609,
25.0540084838867,74.3546524047852,
4.36374855041504,47.8158721923828,
-7.24942111968994,-11.7956132888794,
-2.54607343673706,-44.3182373046875,
13.5543479919434,-45.4090042114258,
31.8960571289063,-47.2745018005371,
44.9289283752441,-54.8113250732422,
42.9997215270996,-37.2510108947754,
20.3075466156006,9.56765937805176,
-10.6472177505493,43.6596298217773,
-22.3492145538330,34.1230583190918,
-7.35317325592041,3.72846150398254,
11.9668083190918,-13.4271373748779,
8.00633144378662,-20.3416023254395,
-14.6444072723389,-36.7482261657715,
-24.1550292968750,-46.2894477844238,
3.30838537216187,-15.2953300476074,
43.4025955200195,42.9308967590332,
44.1138114929199,73.2724533081055,
-8.01223945617676,54.4487953186035,
-65.2030410766602,22.0810203552246,
-68.5405578613281,19.7086601257324,
-20.3517971038818,26.2919998168945,
18.5278911590576,9.50078582763672,
6.23155927658081,-13.8888015747070,
-35.4402351379395,-0.961330890655518,
-51.0716438293457,35.6085014343262,
-31.4349060058594,40.6616706848145,
-11.2649841308594,0.626431703567505,
-4.35668992996216,-37.4682083129883,
10.7189245223999,-28.5397262573242,
38.1357688903809,8.75995063781738,
43.9426994323731,25.0720310211182,
10.1976394653320,10.3210258483887,
-27.6302795410156,-13.8786840438843,
-23.2776832580566,-39.0218467712402,
6.27703619003296,-68.0185317993164,
10.0450220108032,-79.6887435913086,
-12.0007438659668,-49.2768936157227,
-13.3391199111938,-2.17536449432373,
27.6298618316650,7.82274818420410,
58.1693267822266,-18.5275669097900,
31.0649948120117,-24.4603042602539,
-18.6746368408203,15.5591163635254,
-25.1543178558350,51.7511520385742,
9.98105430603027,30.0609626770020,
27.4833259582520,-25.6997776031494,
-3.69632291793823,-42.0842742919922,
-47.1496887207031,-7.41233921051025,
-55.3840789794922,18.2803592681885,
-23.2631416320801,0.806377768516541,
20.7608127593994,-20.2769660949707,
47.4617767333984,-9.18592262268066,
42.4254264831543,17.6796512603760,
2.10785698890686,28.5103168487549,
-51.3636932373047,27.1838893890381,
-68.0192489624023,35.3340034484863,
-28.9124851226807,36.5995674133301,
21.8554439544678,6.55361366271973,
29.4974689483643,-32.6662254333496,
5.06933784484863,-30.3770961761475,
-5.93544340133667,19.9253711700439,
4.66001033782959,59.6116943359375,
0.993821859359741,49.3297576904297,
-34.5199279785156,18.6355056762695,
-65.9735412597656,8.51397323608398,
-59.0542793273926,3.78035783767700,
-35.6800537109375,-27.0788879394531,
-36.1743354797363,-67.7238616943359,
-45.9819145202637,-67.5884246826172,
-22.6497879028320,-18.2124671936035,
27.6988449096680,28.9150009155273,
53.7384414672852,29.3104953765869,
34.3101501464844,-2.71640706062317,
13.2099285125732,-23.3540515899658,
23.1462783813477,-23.3500518798828,
40.1693000793457,-27.7736129760742,
22.2111225128174,-43.7039451599121,
-21.1883487701416,-52.1776695251465,
-42.2666587829590,-42.8791351318359,
-20.5130004882813,-29.9578571319580,
11.8082008361816,-25.2848682403564,
25.1977863311768,-30.2657566070557,
25.0371398925781,-34.0219688415527,
24.6930828094482,-27.7744846343994,
16.1549682617188,-9.67691612243652,
-0.827318012714386,10.6026163101196,
-11.1896944046021,15.8578720092773,
-2.81325888633728,-4.10089254379273,
2.28274393081665,-34.0000534057617,
-17.5737380981445,-37.3452758789063,
-44.7334022521973,-4.11168098449707,
-47.7165069580078,30.6852226257324,
-28.6087493896484,32.0130996704102,
-23.1558284759522,14.5376462936401,
-45.9966506958008,15.9906253814697,
-61.7700347900391,35.9463157653809,
-35.7399177551270,36.7545089721680,
10.1056270599365,6.11883831024170,
28.5624294281006,-15.8443470001221,
13.1085681915283,6.12329673767090,
2.14553022384644,48.1320877075195,
23.5052909851074,51.4748954772949,
57.3771743774414,9.89269161224365,
63.3376197814941,-28.1983299255371,
30.2014141082764,-25.7819843292236,
-13.1643781661987,3.00477790832520,
-30.6923408508301,22.0654621124268,
-15.0523862838745,23.1778411865234,
11.0338287353516,24.1646499633789,
18.7302894592285,27.6207790374756,
0.876680135726929,28.5657215118408,
-18.9514732360840,28.5268535614014,
-11.5616941452026,37.2449340820313,
17.6998081207275,43.2059288024902,
28.9396228790283,25.4939498901367,
2.73004531860352,-22.4028224945068,
-32.9289550781250,-67.7930221557617,
-36.8590965270996,-73.6204452514648,
-7.38417243957520,-45.3728370666504,
17.0712318420410,-23.0219211578369,
12.2390775680542,-27.6125087738037,
-2.74309039115906,-42.4066925048828,
1.17950212955475,-33.6989440917969,
14.4358911514282,7.24029922485352,
12.4028863906860,45.5695877075195,
0.404797077178955,46.5410766601563,
4.01434278488159,18.5119457244873,
28.2297725677490,3.57286047935486,
43.6419372558594,30.9307117462158,
27.1097297668457,75.9280776977539,
-1.69425594806671,81.4579010009766,
-10.4741153717041,31.9830646514893,
-1.06591701507568,-26.4989261627197,
-0.688565969467163,-31.7859268188477,
-17.8349304199219,8.98491477966309,
-31.9761695861816,23.9797401428223,
-24.4528369903564,-20.4068050384522,
-9.14948368072510,-75.7126235961914,
-6.88427257537842,-69.3181991577148,
-8.80643367767334,-3.00959920883179,
6.47152566909790,49.7706375122070,
34.2016220092773,35.8201217651367,
41.5958671569824,-11.1245441436768,
12.4983549118042,-30.5673122406006,
-25.0293483734131,-15.8929882049561,
-31.4810333251953,6.17925453186035,
-1.37327909469605,26.8977012634277,
22.8210296630859,52.4652748107910,
9.81324005126953,67.1787033081055,
-24.3635635375977,39.9067497253418,
-40.2171897888184,-12.1599054336548,
-20.9235992431641,-34.6890983581543,
11.3091831207275,-14.1623792648315,
21.9790077209473,-0.115367025136948,
3.35248756408691,-27.4640541076660,
-17.2070350646973,-54.3184547424316,
-15.5986785888672,-23.9823417663574,
-0.616665840148926,35.9756431579590,
3.53029727935791,44.9662971496582,
-4.91303634643555,-9.36100769042969,
0.505510389804840,-48.3168411254883,
34.1652984619141,-24.6312599182129,
68.2217712402344,14.9444942474365,
55.8371276855469,14.1496849060059,
2.36828565597534,-9.09889793395996,
-32.3691062927246,-2.94318771362305,
-14.2088699340820,22.4869422912598,
22.1599636077881,18.4505996704102,
26.5802574157715,-17.6724338531494,
2.42857789993286,-24.4478797912598,
-5.73449754714966,26.1453247070313,
12.1323127746582,73.4740982055664,
13.2558908462524,55.7100105285645,
-20.0711174011230,-7.25777673721314,
-43.6002960205078,-51.2853393554688,
-18.0939483642578,-53.5056457519531,
23.5688533782959,-33.2418746948242,
18.4626407623291,-9.56670284271240,
-29.7707901000977,11.9961366653442,
-53.7306632995606,22.3488712310791,
-19.0686473846436,11.5678806304932,
25.5516834259033,-3.23191404342651,
21.9645290374756,10.0573253631592,
-15.8886260986328,39.8671798706055,
-26.0025596618652,38.3756027221680,
11.6196050643921,-7.65261077880859,
51.3952445983887,-43.7855911254883,
47.4039649963379,-23.8128356933594,
8.02310943603516,22.0524711608887,
-25.6981277465820,31.1642436981201,
-33.9964294433594,3.49633622169495,
-27.9052906036377,-5.84796762466431,
-18.9086456298828,27.3276386260986,
-2.45256233215332,55.3728637695313,
16.7125549316406,26.8818416595459,
25.4237709045410,-32.4589767456055,
17.7566242218018,-52.2191658020020,
4.03318977355957,-10.0739669799805,
3.89237523078918,43.8553466796875,
22.2861347198486,54.4927978515625,
32.7407150268555,24.0259075164795,
13.6755437850952,-0.639036536216736,
-20.9095191955566,6.06836462020874,
-37.0515136718750,26.9709930419922,
-20.1654472351074,30.3860301971436,
6.03255844116211,4.18515443801880,
-1.70301866531372,-24.0979156494141,
-43.6395950317383,-23.8885574340820,
-67.8054733276367,2.83017301559448,
-39.2945632934570,27.0969810485840,
11.9597148895264,23.5760688781738,
21.9058513641357,-6.36127853393555,
-19.9562950134277,-34.4826812744141,
-48.0141716003418,-36.7195434570313,
-13.9640140533447,-16.1464195251465,
46.0433235168457,13.2493753433228,
54.2912864685059,37.5879478454590,
-1.07746958732605,42.0129814147949,
-41.9495429992676,16.2060585021973,
-11.8846521377563,-34.1071510314941,
46.5936698913574,-74.4852066040039,
53.5176658630371,-65.7200622558594,
-1.19845390319824,-13.4004144668579,
-53.6839637756348,26.7042236328125,
-57.9197387695313,10.5985202789307,
-30.2469749450684,-39.6002616882324,
-11.4198894500732,-56.7711830139160,
-14.1301345825195,-12.6562585830688,
-32.1979331970215,45.3726158142090,
-56.6545295715332,46.3484840393066,
-70.4482803344727,-11.9248943328857,
-44.2591209411621,-63.2459526062012,
17.3418865203857,-55.3732528686523,
59.8471832275391,-5.61435461044312,
40.6901893615723,24.2154808044434,
-3.28233599662781,6.62599754333496,
-9.04082775115967,-27.5330734252930,
21.4026203155518,-36.9884910583496,
26.7822780609131,-14.6660776138306,
-13.6464099884033,13.9061861038208,
-45.6731033325195,30.6094074249268,
-27.7700653076172,33.8379554748535,
4.62859487533569,29.6659393310547,
-8.20129108428955,17.0450782775879,
-43.3266487121582,-6.23275995254517,
-30.7658023834229,-35.0070800781250,
33.0233116149902,-47.2682533264160,
68.1546020507813,-27.8366336822510,
32.3804130554199,8.97572326660156,
-21.0840034484863,30.8890419006348,
-18.1256732940674,13.9170894622803,
30.5075321197510,-26.0636730194092,
57.1081352233887,-45.1660156250000,
33.5796356201172,-23.0301132202148,
-8.67001628875732,10.3215122222900,
-36.0202789306641,18.4270229339600,
-49.8170776367188,-1.97686028480530,
-59.5611381530762,-24.5801792144775,
-52.8439788818359,-33.7044944763184,
-19.8338871002197,-33.6956520080566,
16.1805400848389,-27.9122123718262,
32.2959442138672,-10.0788230895996,
37.6129035949707,14.7258739471436,
47.3275604248047,18.8595790863037,
53.4199829101563,-9.69760513305664,
35.9757270812988,-39.4790115356445,
4.36080455780029,-38.4867935180664,
-13.9511852264404,-18.4488391876221,
-8.52818298339844,-18.7251224517822,
5.56433105468750,-45.2275238037109,
11.2636613845825,-55.3806419372559,
14.1877365112305,-26.8659954071045,
18.5370349884033,7.69192981719971,
11.5005512237549,0.798813104629517,
-9.90715312957764,-39.4795875549316,
-20.7849559783936,-61.3618278503418,
1.87471902370453,-32.0290756225586,
35.4258956909180,20.3468132019043,
37.5697937011719,53.3538551330566,
-5.42124414443970,55.1338233947754,
-59.4619140625000,44.5924758911133,
-79.3276672363281,34.0855979919434,
-54.8190193176270,22.3011093139648,
-5.64591598510742,6.48051166534424,
38.6022300720215,-5.93330717086792,
55.7019882202148,-13.2857923507690,
35.9485588073731,-17.8610916137695,
-4.42833518981934,-23.2849540710449,
-25.3433628082275,-30.6337642669678,
-4.07076549530029,-41.3110008239746,
34.2969589233398,-52.0548820495606,
39.7128868103027,-57.4315910339356,
2.32644915580750,-47.3625488281250,
-37.9387130737305,-23.6299533843994,
-41.3810043334961,-7.85448074340820,
-14.4684982299805,-13.1364850997925,
9.43972873687744,-29.4151477813721,
9.47487068176270,-33.6498069763184,
1.51045334339142,-11.7232456207275,
3.43419528007507,24.0003032684326,
11.1802730560303,49.6754226684570,
15.0688915252686,44.4585456848145,
12.0542182922363,13.5999584197998,
7.38838958740234,-19.6518840789795,
6.43730163574219,-23.7779388427734,
13.2483777999878,8.39482975006104,
25.8015975952148,47.9725151062012,
34.1598739624023,54.3475341796875,
27.2039546966553,24.1420345306397,
14.4926633834839,-9.86680698394775,
18.6559753417969,-18.0827713012695,
46.2461891174316,-9.87652015686035,
72.6624603271484,-8.89038562774658,
61.7413749694824,-12.4271125793457,
15.4985933303833,4.76714324951172,
-27.0745639801025,37.7837677001953,
-40.8169937133789,47.4215621948242,
-36.7647590637207,5.74885606765747,
-29.1722640991211,-57.0170135498047,
-13.5705966949463,-81.1268005371094,
19.4911594390869,-53.9024925231934,
54.4573898315430,-16.5718288421631,
66.9154968261719,-9.75423431396484,
53.3085670471191,-24.8298835754395,
32.9239540100098,-24.8908329010010,
11.0169601440430,1.53421568870544,
-18.6053543090820,30.8396663665772,
-44.5775260925293,34.9889259338379,
-33.5757217407227,6.88378715515137,
12.5417470932007,-31.9923725128174,
43.7411727905273,-53.5395011901856,
16.7257118225098,-41.6455497741699,
-34.1664085388184,-3.87589597702026,
-43.2021293640137,30.0656013488770,
0.953303813934326,33.2373161315918,
44.8714675903320,9.89398956298828,
46.5063400268555,-10.1480741500855,
28.6332740783691,-10.1804361343384,
32.9431686401367,-1.94098067283630,
53.7779312133789,2.66250991821289,
54.3565597534180,1.98929214477539,
30.1833419799805,-1.58301353454590,
13.3215932846069,-18.0088825225830,
21.2348537445068,-45.0387229919434,
36.1260986328125,-55.2805061340332,
35.9254760742188,-22.7520084381104,
24.2082061767578,25.5376682281494,
10.9413385391235,35.9300384521484,
2.02975988388062,0.552878201007843,
6.87445116043091,-27.6713218688965,
27.7718086242676,2.09280467033386,
48.9114646911621,62.7943649291992,
40.5182380676270,83.3744049072266,
-7.08223342895508,42.9597892761231,
-49.7841262817383,-11.4672422409058,
-38.4720993041992,-24.4804344177246,
14.7217206954956,2.35066151618958,
53.4978446960449,29.0135421752930,
46.9432754516602,33.7235107421875,
20.6297988891602,30.0555725097656,
-0.00749474763870239,34.2373809814453,
-15.4807424545288,39.1790580749512,
-26.9005718231201,28.5776710510254,
-16.0596580505371,0.707162141799927,
26.2243671417236,-30.1388740539551,
60.2886695861816,-41.4778861999512,
36.2473373413086,-17.1800212860107,
-31.9268169403076,25.2755584716797,
-74.7039794921875,45.8132667541504,
-54.2071151733398,24.0771923065186,
-5.39350891113281,-19.8422412872314,
20.8230857849121,-44.1059951782227,
19.3993320465088,-33.5972480773926,
10.9941635131836,-15.2505340576172,
-4.87474822998047,-10.8175992965698,
-33.8062705993652,-5.98263740539551,
-53.5439758300781,19.1233444213867,
-33.8509559631348,42.9856948852539,
10.4768342971802,31.8543739318848,
27.1586494445801,-0.813556194305420,
-2.30773210525513,-6.70965099334717,
-36.8502731323242,29.9559593200684,
-32.1462249755859,55.3078155517578,
-7.84469175338745,14.7717046737671,
-7.50777626037598,-64.7833557128906,
-25.4225845336914,-105.297225952148,
-22.3144664764404,-68.8172302246094,
7.27083301544189,2.10775566101074,
32.3962860107422,40.6089897155762,
23.9805660247803,29.0365123748779,
-1.13756716251373,-4.04423379898071,
-11.1842966079712,-32.7573966979981,
2.04768323898315,-42.8906059265137,
25.9925041198730,-30.9084663391113,
45.3602523803711,-1.00239062309265,
42.4062004089356,29.8377971649170,
1.00920534133911,44.3340835571289,
-59.9866180419922,34.3919143676758,
-83.1472320556641,11.1442003250122,
-43.1330986022949,-13.1494960784912,
10.5394058227539,-29.2238006591797,
13.0383691787720,-32.8521804809570,
-28.5017833709717,-22.2609424591064,
-44.1168441772461,-13.8933086395264,
-1.30430042743683,-25.0223159790039,
51.2556343078613,-38.9637680053711,
56.1040916442871,-24.3445205688477,
25.6245746612549,19.3682403564453,
10.4585418701172,49.5792922973633,
16.0373249053955,30.1866245269775,
3.57397627830505,-11.7054758071899,
-28.3109397888184,-18.1273937225342,
-36.1139526367188,23.3833236694336,
-1.56538200378418,62.8181152343750,
36.6431503295898,54.2246437072754,
34.0568199157715,18.4418201446533,
7.76583480834961,8.97996997833252,
-3.58942532539368,38.2579002380371,
10.0648565292358,67.3874511718750,
18.2235374450684,60.2583122253418,
9.25581169128418,27.0879554748535,
1.69495832920074,2.63417148590088,
11.1840972900391,3.43583512306213,
24.0155735015869,14.8546628952026,
27.6153087615967,16.6115970611572,
36.6934661865234,1.15087866783142,
55.1053619384766,-23.8086452484131,
59.6939353942871,-40.5903549194336,
33.3942909240723,-37.1238899230957,
-7.06519412994385,-16.1573257446289,
-31.4403209686279,0.978415131568909,
-34.8634757995606,-4.38646173477173,
-37.8488121032715,-20.5682430267334,
-54.1252326965332,-23.1778926849365,
-68.8411865234375,-3.18701648712158,
-67.9719543457031,19.3995780944824,
-53.8436889648438,24.0001983642578,
-31.1996955871582,9.20209026336670,
1.82247173786163,-9.07403087615967,
27.4878101348877,-25.3802413940430,
20.7067012786865,-43.3714523315430,
-11.2470169067383,-58.6472244262695,
-21.0605640411377,-55.1340065002441,
15.1901750564575,-31.0390262603760,
56.8690109252930,-3.41290998458862,
44.4073181152344,7.13165616989136,
-10.5397443771362,2.34959602355957,
-39.8516159057617,-1.87877488136292,
-10.3043193817139,2.49638128280640,
30.6902980804443,10.7274942398071,
27.5507926940918,15.1489534378052,
-1.81790852546692,13.3445873260498,
-0.669118642807007,4.51261234283447,
35.0794372558594,-8.33273792266846,
58.3425216674805,-17.7359180450439,
38.9493370056152,-9.88499736785889,
4.71276140213013,12.7988691329956,
-7.70141696929932,32.0440635681152,
-2.88747143745422,28.6739788055420,
-6.52668380737305,3.13772153854370,
-18.1326599121094,-23.3489112854004,
-18.0641059875488,-39.9388008117676,
-3.58396911621094,-42.8868217468262,
8.14021301269531,-36.8460769653320,
6.86433458328247,-26.4300613403320,
7.75476026535034,-10.3026561737061,
21.1292457580566,9.07670211791992,
27.7497863769531,26.5834045410156,
14.5144453048706,36.9985008239746,
-4.91108179092407,38.4625663757324,
-4.11930084228516,35.7361412048340,
14.9777669906616,40.0920410156250,
21.5918712615967,50.7356376647949,
-6.07563161849976,46.7969589233398,
-42.4371795654297,7.66547155380249,
-45.8840141296387,-41.5025825500488,
-13.7041273117065,-49.0493469238281,
12.0938758850098,-4.13066625595093,
-1.26922440528870,40.0757141113281,
-33.6234130859375,25.1866455078125,
-38.5086669921875,-33.7160263061523,
0.374560117721558,-64.5703353881836,
44.6567382812500,-36.9060707092285,
52.0283050537109,2.90084385871887,
24.3112659454346,0.482796907424927,
0.599207401275635,-27.6701030731201,
5.61741304397583,-32.7089920043945,
22.4965877532959,-11.6064252853394,
20.9902572631836,-9.88919639587402,
-1.30313074588776,-43.6202583312988,
-18.3606739044189,-68.6489181518555,
-10.7051496505737,-44.4427375793457,
6.10683631896973,7.30060195922852,
2.05290532112122,33.6095962524414,
-26.7368125915527,20.8790187835693,
-48.8981704711914,-1.64858555793762,
-37.1854438781738,-10.7110223770142,
3.16131877899170,-13.0538282394409,
38.0100975036621,-17.8381671905518,
43.9644203186035,-12.3002586364746,
28.1937904357910,11.7998867034912,
11.2213935852051,33.6629066467285,
2.08577299118042,28.6006183624268,
1.53495347499847,0.852483868598938,
6.19773483276367,-26.4491691589355,
8.82520198822022,-40.1819839477539,
6.43260002136231,-46.4275856018066,
5.84423255920410,-50.4102935791016,
22.6783370971680,-44.4919395446777,
54.3871955871582,-18.0990085601807,
69.7183303833008,14.3563833236694,
37.7031059265137,29.2751140594482,
-26.1671390533447,22.3385276794434,
-68.7508316040039,7.22889804840088,
-61.2220115661621,-0.987199306488037,
-27.8576068878174,-1.19982445240021,
-14.8979206085205,-4.85800123214722,
-25.8984565734863,-18.5893516540527,
-25.5138931274414,-34.1443061828613,
2.80965900421143,-31.2100200653076,
35.1101760864258,-3.55376672744751,
38.9213294982910,27.0350933074951,
17.8970260620117,30.7962627410889,
6.09691381454468,0.305262923240662,
18.5678844451904,-27.2241916656494,
39.2181053161621,-17.1975212097168,
42.1048202514648,19.9368972778320,
23.1542205810547,36.9373130798340,
-1.17294597625732,15.2392215728760,
-13.2507982254028,-11.5446949005127,
-7.90610694885254,-8.46642398834229,
10.3169984817505,13.3184585571289,
32.1815414428711,19.1987304687500,
40.6408462524414,5.90800571441650,
26.3484115600586,3.27704453468323,
-1.78270220756531,18.4224224090576,
-19.0129661560059,21.6686000823975,
-10.4302139282227,-10.7701578140259,
19.8806953430176,-50.7669525146484,
46.4396286010742,-57.3782539367676,
50.4312553405762,-29.7618961334229,
30.1301422119141,-0.623298585414887,
-1.82239055633545,11.9156723022461,
-32.5982780456543,13.9421901702881,
-51.1902465820313,8.62431144714356,
-51.9213905334473,-5.07568693161011,
-37.5676651000977,-12.1841735839844,
-17.4793376922607,6.83351707458496,
-6.36126756668091,42.6742057800293,
-13.9827966690063,58.9500961303711,
-33.4180450439453,39.5207595825195,
-36.8459129333496,20.6231365203857,
-6.44728231430054,35.8269386291504,
41.0346641540527,56.6426086425781,
63.4612960815430,35.3469085693359,
42.9937515258789,-16.8242721557617,
8.03948020935059,-38.2233238220215,
2.78102469444275,-8.35560798645020,
18.5332336425781,23.2112846374512,
10.9772319793701,11.1044950485230,
-31.9636936187744,-20.0117778778076,
-63.4276657104492,-18.6422462463379,
-42.9044036865234,5.32352638244629,
-4.50283479690552,-0.623325943946838,
-0.833542466163635,-47.0793991088867,
-27.4257087707520,-78.6252899169922,
-23.0206680297852,-56.6068725585938,
31.0586738586426,-15.4679212570190,
81.6550216674805,-9.45669937133789,
76.6208877563477,-30.1059455871582,
39.6420440673828,-30.9841041564941,
27.9075145721436,3.24276494979858,
46.6521072387695,32.9425506591797,
52.6428909301758,31.7649040222168,
29.9880981445313,14.4561300277710,
5.02291774749756,12.8194885253906,
-5.55484056472778,27.7575454711914,
-17.6348819732666,37.3590431213379,
-40.5380706787109,35.9825973510742,
-51.5711212158203,32.2230834960938,
-43.1922607421875,26.0662899017334,
-35.1076087951660,11.2820186614990,
-46.9457588195801,-8.70508384704590,
-59.6269454956055,-15.8986425399780,
-46.8203048706055,-7.61498165130615,
-23.5810298919678,-0.190191805362701,
-25.9377365112305,-11.7214775085449,
-43.1059265136719,-34.5072059631348,
-25.4861812591553,-49.4010353088379,
31.6251525878906,-49.8838272094727,
77.6982955932617,-47.3158493041992,
67.5420684814453,-42.7026901245117,
21.4151687622070,-22.8815708160400,
-17.6740837097168,13.0809373855591,
-38.6280746459961,37.8959617614746,
-55.1808128356934,21.1073570251465,
-60.9353446960449,-25.2511177062988,
-38.9015388488770,-50.8515930175781,
3.39485073089600,-30.3478298187256,
28.1029109954834,6.35413312911987,
21.4370899200439,14.9908132553101,
13.5197887420654,-4.78646945953369,
31.1107444763184,-15.5063419342041,
53.9940185546875,-0.685927391052246,
46.1785392761231,16.0805263519287,
3.65383672714233,12.5718832015991,
-37.8462028503418,8.68705844879150,
-48.1980590820313,20.6359672546387,
-29.8992557525635,30.1542758941650,
-5.18709564208984,5.05517196655273,
2.09896540641785,-36.4100341796875,
-8.44227886199951,-46.2319869995117,
-25.6022720336914,-14.9935951232910,
-28.5122108459473,10.0916109085083,
-6.50524616241455,-5.42326831817627,
31.3067150115967,-30.9280147552490,
58.0292549133301,-22.0470943450928,
55.9482498168945,11.4641199111938,
34.0721244812012,20.5691013336182,
15.6573753356934,-4.22862529754639,
15.8266210556030,-16.4585475921631,
24.3386306762695,16.6175327301025,
23.7330799102783,64.6883926391602,
2.59274792671204,77.6044311523438,
-28.0412120819092,52.2106437683106,
-47.4461402893066,25.2975254058838,
-47.8136749267578,16.2179908752441,
-34.3045959472656,5.49080419540405,
-15.7187824249268,-20.0795631408691,
3.87036561965942,-42.9835014343262,
20.5410804748535,-33.0129661560059,
25.5672473907471,2.24955272674561,
13.1260051727295,23.5603675842285,
-6.67301082611084,9.15554523468018,
-8.98582935333252,-16.2987937927246,
15.6418571472168,-14.4707107543945,
42.0106620788574,16.2877807617188,
38.4434432983398,42.2893981933594,
5.78710269927979,37.0669479370117,
-19.0119934082031,11.6430130004883,
-6.23137474060059,-2.95625734329224,
26.2385177612305,0.501882433891296,
32.0791969299316,1.66842567920685,
-1.90941786766052,-10.3141775131226,
-35.0961494445801,-22.9029712677002,
-24.3730716705322,-23.1109123229980,
19.2521877288818,-17.1618785858154,
38.2287368774414,-15.6865673065186,
6.79915237426758,-13.8543529510498,
-41.7748336791992,3.37452912330627,
-55.3429450988770,29.0839252471924,
-35.7689666748047,36.9817008972168,
-23.6624755859375,17.2974472045898,
-32.4304618835449,-15.5262660980225,
-29.5177955627441,-39.1910514831543,
11.5962467193604,-47.0350799560547,
66.2532501220703,-40.5789146423340,
81.9159927368164,-20.2704429626465,
45.4785003662109,12.4724235534668,
-3.14357089996338,42.7462730407715,
-24.7390251159668,51.8193283081055,
-17.8441963195801,41.4299812316895,
-1.93250465393066,24.2197322845459,
14.8104600906372,7.19450187683106,
39.6390151977539,-13.3888530731201,
64.3331680297852,-27.0112915039063,
64.5895004272461,-12.1783838272095,
30.3179206848145,26.3722953796387,
-12.7316665649414,56.9553833007813,
-30.6131629943848,51.9932823181152,
-17.9237537384033,22.8662910461426,
-1.30694651603699,5.16106605529785,
-5.01444149017334,14.3480663299561,
-26.3577404022217,31.1676025390625,
-34.7404975891113,37.0388946533203,
-10.7398891448975,32.6746368408203,
25.2989730834961,29.2061176300049,
42.1844062805176,30.5424461364746,
19.2712574005127,37.4390258789063,
-26.5988731384277,47.3928108215332,
-61.0063476562500,43.3764610290527,
-65.9240493774414,10.6699867248535,
-46.7941246032715,-40.2136993408203,
-17.7404365539551,-70.2880859375000,
17.9809093475342,-55.7025604248047,
46.4517478942871,-24.0718421936035,
42.4579277038574,-14.2956180572510,
0.609200000762940,-26.4553794860840,
-47.0750198364258,-21.4329490661621,
-49.8303718566895,9.09877204895020,
-4.03919601440430,23.4810390472412,
37.5498733520508,-7.24123096466064,
27.9163284301758,-46.7557220458984,
-17.5772037506104,-45.0905303955078,
-47.1141128540039,-3.96728563308716,
-39.3486709594727,22.5344944000244,
-17.2755203247070,7.42549896240234,
-1.66856646537781,-17.2457370758057,
15.7306766510010,-9.30647087097168,
36.6823425292969,24.7942829132080,
36.8514595031738,52.1307601928711,
1.20434188842773,53.2928047180176,
-47.4932250976563,36.8655776977539,
-69.2969589233398,10.5642223358154,
-53.1756668090820,-15.6705837249756,
-22.8837089538574,-23.2769470214844,
1.37326812744141,1.72536349296570,
16.2297916412354,30.1625022888184,
19.0885124206543,21.7774333953857,
4.12889051437378,-21.5642280578613,
-13.9648866653442,-54.0266418457031,
-6.89952850341797,-40.1094017028809,
18.7403869628906,1.87651336193085,
22.3387393951416,21.8932895660400,
-9.56999588012695,8.69444179534912,
-35.6155433654785,-9.25616455078125,
-14.5134334564209,-13.1866607666016,
26.5791339874268,-5.81991815567017,
23.9495735168457,4.38777065277100,
-30.1910152435303,5.90130710601807,
-72.2934341430664,-15.3583707809448,
-49.7070045471191,-59.2285499572754,
5.91158008575439,-87.3723373413086,
32.0858039855957,-56.0431938171387,
18.6319198608398,17.2659549713135,
5.04146003723145,59.9837493896484,
12.3933153152466,33.7229919433594,
23.8110198974609,-12.4776506423950,
21.4409923553467,-6.37014532089233,
7.76137256622314,43.8623580932617,
-3.57046771049500,57.4956359863281,
-10.0329523086548,5.02902507781982,
-11.9299592971802,-54.1507987976074,
-10.4868230819702,-59.2579460144043,
-12.2532777786255,-23.0561504364014,
-27.6331787109375,1.98241209983826,
-43.2551307678223,-1.07726287841797,
-22.9443244934082,-8.26560974121094,
29.4811325073242,-5.74772834777832,
52.7621002197266,-6.88575220108032,
10.6746034622192,-11.8873662948608,
-45.9422645568848,-2.42508411407471,
-41.5777816772461,17.3697433471680,
18.4454269409180,16.4510898590088,
51.8571357727051,-11.7797918319702,
17.8720703125000,-26.6233577728272,
-31.6978607177734,-2.06576037406921,
-31.9215164184570,26.0253448486328,
-7.22134780883789,15.7091979980469,
-16.6574840545654,-15.7124471664429,
-50.6836280822754,-19.1383686065674,
-43.6454772949219,8.12538528442383,
12.5011196136475,16.2859115600586,
53.6805038452148,-18.4678287506104,
41.3078079223633,-44.9733772277832,
11.6022624969482,-7.83600807189941,
6.03475284576416,64.0002517700195,
10.7875728607178,92.3365325927734,
-1.16356956958771,51.5455627441406,
-10.1481771469116,-8.76113128662109,
18.1125907897949,-31.9552707672119,
57.1651077270508,-8.19771766662598,
48.6838302612305,35.9780540466309,
-4.37364673614502,69.4052429199219,
-34.9164695739746,70.5275726318359,
-18.9576606750488,42.1793327331543,
-11.2913866043091,10.3779764175415,
-44.3671760559082,4.01751089096069,
-68.4480514526367,16.4521694183350,
-27.1585903167725,8.11375141143799,
38.1322174072266,-33.1506881713867,
42.3559036254883,-57.7620277404785,
-19.1316833496094,-23.2283668518066,
-59.6067008972168,31.2918167114258,
-20.7199192047119,40.5827331542969,
49.7760429382324,4.35943698883057,
70.2874221801758,-23.0496749877930,
33.6002998352051,-14.0482940673828,
-5.56894588470459,-7.43954133987427,
-17.6643295288086,-37.7312088012695,
-22.6655158996582,-69.3929748535156,
-31.9664478302002,-53.9658737182617,
-32.3177795410156,-14.3554325103760,
-8.97798538208008,-1.59736061096191,
26.9249572753906,-16.8793106079102,
44.9985771179199,-8.99009513854981,
31.9930839538574,31.3915367126465,
-3.28636837005615,43.8125762939453,
-33.7101364135742,-5.95430660247803,
-35.5392608642578,-62.8340072631836,
-6.29950237274170,-55.9050674438477,
25.3061332702637,0.853905797004700,
19.5597705841064,28.8658218383789,
-14.9666528701782,-5.98824691772461,
-23.3239593505859,-47.5556488037109,
15.8391828536987,-31.3538417816162,
54.4076194763184,24.7779140472412,
37.6259155273438,51.9518623352051,
-18.5620632171631,22.7271766662598,
-44.5004158020020,-19.5269336700439,
-10.8350791931152,-26.9748630523682,
36.5005950927734,3.44724392890930,
43.3034553527832,36.9161415100098,
18.5249919891357,43.6135864257813,
0.826327323913574,29.1345062255859,
-8.69184207916260,14.7415103912354,
-28.9626617431641,13.6000642776489,
-44.2439155578613,15.8180875778198,
-25.2772769927979,8.34212875366211,
14.2307786941528,-10.4956645965576,
16.7302246093750,-24.2382678985596,
-29.8985767364502,-15.8656435012817,
-60.6842727661133,5.07478284835815,
-27.1569480895996,12.8827295303345,
33.8323326110840,5.25803232192993,
47.0074386596680,4.38498973846436,
2.47558736801147,22.8366527557373,
-34.9169731140137,39.5205383300781,
-21.8363704681397,21.2853755950928,
5.91938686370850,-27.5901813507080,
7.86810064315796,-62.3593063354492,
-2.87266993522644,-54.6229591369629,
9.79308700561523,-26.2976703643799,
45.0737037658691,-13.8074550628662,
65.7240295410156,-20.3334159851074,
50.5115852355957,-15.8835849761963,
9.60291004180908,10.2152318954468,
-33.8900299072266,29.9682140350342,
-62.7754707336426,15.5160083770752,
-63.9574165344238,-19.3656349182129,
-36.5373573303223,-39.0704383850098,
-8.08843994140625,-25.2372226715088,
-16.1327304840088,3.81513500213623,
-56.5591697692871,19.8897399902344,
-72.9132537841797,15.9501771926880,
-33.3056259155273,7.32171058654785,
29.3479442596436,9.08884906768799,
58.0341224670410,18.6761703491211,
37.1562461853027,22.5012245178223,
3.35006475448608,10.8750343322754,
-12.8525867462158,-9.81105709075928,
-14.9200725555420,-18.1653785705566,
-18.0056934356689,-5.80468988418579,
-18.7978820800781,6.48428392410278,
-6.76319980621338,-4.41818523406982,
10.0595149993896,-30.7575283050537,
20.4627437591553,-43.9458122253418,
28.4394569396973,-31.1527709960938,
46.8432960510254,-10.8683853149414,
63.1562194824219,-9.93192768096924,
57.6413688659668,-24.1352996826172,
33.9295463562012,-29.2969360351563,
18.5515403747559,-23.5583953857422,
24.1177024841309,-21.4961643218994,
40.4975662231445,-25.4478225708008,
46.3481178283691,-19.4642448425293,
41.3499641418457,-8.25965976715088,
34.8691291809082,-15.1811981201172,
25.8805866241455,-43.1224365234375,
10.8226919174194,-54.4298973083496,
4.56006145477295,-23.6019153594971,
15.0562429428101,13.9079647064209,
21.4983654022217,7.88241434097290,
-0.346501350402832,-33.9487609863281,
-32.3266906738281,-45.9983291625977,
-30.4899215698242,1.70141685009003,
10.3730487823486,55.8152961730957,
36.8790740966797,61.0034408569336,
6.89597511291504,30.2710037231445,
-48.7736740112305,11.8465337753296,
-61.8421554565430,8.79793834686279,
-19.1617965698242,-6.60672950744629,
30.2292327880859,-36.4966773986816,
46.4209136962891,-44.3450241088867,
45.7602157592773,-19.8290748596191,
50.6242103576660,4.63537311553955,
52.1583442687988,6.62063312530518,
31.3430252075195,13.6011486053467,
4.67823076248169,44.0439491271973,
-1.36119842529297,65.7365875244141,
6.90817832946777,37.6565246582031,
-0.593199372291565,-17.9825916290283,
-29.9567489624023,-38.9705390930176,
-51.1610527038574,-18.8086795806885,
-43.6410217285156,-8.22369861602783,
-21.4731426239014,-33.7572021484375,
-4.32128047943115,-66.7766799926758,
16.0720748901367,-62.7969741821289,
47.2142410278320,-32.4571685791016,
65.7449722290039,-11.5712928771973,
51.3303222656250,-7.13329124450684,
14.7457923889160,4.73916339874268,
-12.7184782028198,30.5705108642578,
-18.5807247161865,46.5628395080566,
-20.0403213500977,42.1945686340332,
-22.5020713806152,27.9397735595703,
-14.3403844833374,8.45089244842529,
10.4458122253418,-22.6592750549316,
31.4834384918213,-49.1017150878906,
30.2554550170898,-39.4130973815918,
20.6891174316406,13.3293590545654,
25.0948085784912,70.8820419311523,
31.6313056945801,88.8770675659180,
15.2488412857056,69.2265167236328,
-25.0302619934082,44.2707023620606,
-54.8865013122559,31.7873992919922,
-46.9523849487305,14.3464250564575,
-14.0508079528809,-6.54450082778931,
10.0059118270874,-10.5289630889893,
7.70478630065918,8.46539878845215,
-9.37903594970703,22.9023723602295,
-23.4666404724121,13.5863265991211,
-24.3112545013428,0.390707433223724,
-8.15468215942383,7.84908294677734,
15.9885959625244,29.2566547393799,
28.4721450805664,35.5970726013184,
12.4868545532227,21.6945934295654,
-19.6464519500732,5.50229835510254,
-36.2067375183106,-1.42825174331665,
-21.5293197631836,-15.1256904602051,
-0.884401917457581,-49.5578956604004,
-1.12202739715576,-79.3636856079102,
-18.9645442962647,-83.7850418090820,
-24.7282257080078,-61.9806022644043,
0.311096429824829,-31.0730094909668,
29.8727378845215,-0.319414854049683,
31.8285999298096,21.9490833282471,
9.56297683715820,22.7057189941406,
-7.98708820343018,1.42258024215698,
1.56901478767395,-17.5275058746338,
25.6443367004395,-10.2059354782105,
33.9496726989746,7.18342018127441,
12.4969444274902,-3.11092281341553,
-13.2370882034302,-37.8840637207031,
-6.56453752517700,-43.6870155334473,
35.9633216857910,9.13183021545410,
69.1272354125977,75.2709579467773,
42.8329467773438,89.9675369262695,
-30.7965698242188,49.4237785339356,
-79.4217834472656,8.23035812377930,
-47.9229240417481,-5.07005119323731,
29.5434226989746,-10.8151254653931,
63.0775070190430,-32.0213775634766,
21.9172039031982,-45.0044670104981,
-36.1563377380371,-19.4471740722656,
-49.7448768615723,27.2962570190430,
-29.3666095733643,45.4427299499512,
-27.5725021362305,21.7083816528320,
-55.2489776611328,-6.09128904342651,
-70.2216873168945,-10.3357782363892,
-42.5534210205078,-3.57810449600220,
2.82541227340698,-7.77553749084473,
34.3468132019043,-20.5501308441162,
49.6861801147461,-25.3641300201416,
52.6274681091309,-19.3231353759766,
31.9702033996582,-5.20359277725220,
-14.7156867980957,11.4246883392334,
-47.6557655334473,31.1805076599121,
-28.6405830383301,38.7770156860352,
14.2962388992310,26.5651721954346,
28.8889408111572,16.0679683685303,
9.29464626312256,29.7277183532715,
-3.72043681144714,50.5192794799805,
11.5318088531494,30.8314456939697,
20.6220436096191,-27.2068328857422,
-6.48472404479981,-64.0248107910156,
-42.0891532897949,-36.5030479431152,
-43.4353523254395,23.2113075256348,
-17.9230670928955,49.7959594726563,
-5.51683902740479,32.9018058776856,
-3.08597707748413,19.2367610931397,
12.6086940765381,37.6084251403809,
31.0892486572266,59.0489044189453,
10.3180093765259,50.8722877502441,
-46.5479202270508,20.8193454742432,
-76.3504028320313,-5.10059595108032,
-39.9220657348633,-25.3945236206055,
22.7530593872070,-48.7332954406738,
43.3628044128418,-55.2150726318359,
12.3884048461914,-20.2450256347656,
-21.1057968139648,39.1831092834473,
-33.6323089599609,68.4863281250000,
-38.9999618530273,42.5515289306641,
-40.1097412109375,-5.87088251113892,
-14.1266975402832,-28.2346782684326,
35.7318572998047,-15.9854202270508,
60.4700851440430,-0.531993925571442,
33.4320640563965,-2.23943805694580,
-13.6342582702637,-14.1935882568359,
-31.3085765838623,-24.9328880310059,
-15.8821725845337,-29.9640865325928,
-0.342325568199158,-26.0124053955078,
1.18586242198944,-12.6050081253052,
5.33675193786621,4.12509822845459,
18.4823474884033,13.4921665191650,
13.3966045379639,13.6798391342163,
-19.2404937744141,12.2005653381348,
-49.3826560974121,11.7281713485718,
-48.4378242492676,6.99075031280518,
-22.9037704467773,-3.02517890930176,
3.63926887512207,-10.3992900848389,
22.8835487365723,-7.18427181243897,
40.1759567260742,-6.32701539993286,
44.9355621337891,-21.4036636352539,
23.2859916687012,-42.6962394714356,
-10.1313066482544,-48.6301689147949,
-22.2829570770264,-37.2706985473633,
-3.02553248405457,-24.8573513031006,
13.9379291534424,-19.2856197357178,
2.55528736114502,-6.78795385360718,
-23.4475288391113,21.2831134796143,
-31.7195911407471,48.8765335083008,
-24.1258106231689,49.4749412536621,
-25.3073387145996,20.2057018280029,
-40.8570899963379,-14.4305019378662,
-46.6119346618652,-32.3660964965820,
-28.0900344848633,-31.6426258087158,
1.94138932228088,-18.8024291992188,
14.0624990463257,-0.0223972797393799,
3.46649885177612,10.0185432434082,
-12.8629121780396,-0.623682379722595,
-23.0848197937012,-21.9878368377686,
-26.7798061370850,-26.2569236755371,
-26.8511047363281,-6.84655141830444,
-30.1809844970703,14.7574758529663,
-42.8946685791016,11.6863451004028,
-61.5743827819824,-7.06229496002197,
-64.8384780883789,-13.1005229949951,
-46.2050170898438,-5.95901441574097,
-30.2355747222900,-8.13286876678467,
-37.3753128051758,-24.2008762359619,
-52.0600738525391,-24.7433509826660,
-33.8524894714356,-2.73809909820557,
18.5988025665283,10.2231035232544,
53.0487556457520,-9.90106582641602,
29.7469310760498,-38.5596771240234,
-17.7390975952148,-34.8232231140137,
-25.6687602996826,-7.73166608810425,
10.2576217651367,-5.10675764083862,
43.4298133850098,-37.3130493164063,
47.7496833801270,-55.8957099914551,
49.4747200012207,-23.0862407684326,
59.5955314636231,29.6051292419434,
49.4918251037598,49.2688446044922,
-1.28891217708588,32.1879730224609,
-50.9353752136231,18.9561328887939,
-45.5213775634766,27.9598770141602,
4.85654735565186,36.5667800903320,
32.1843338012695,30.4159851074219,
7.18381929397583,26.1168766021729,
-30.8928241729736,36.2750892639160,
-41.4169425964356,39.9954223632813,
-35.0654487609863,15.7417926788330,
-38.7989463806152,-17.8238811492920,
-46.7208175659180,-20.5702285766602,
-41.7978935241699,7.92425394058228,
-36.2796325683594,24.5733757019043,
-48.4159393310547,1.70963501930237,
-58.6446189880371,-37.2955284118652,
-31.5930213928223,-50.7621383666992,
19.5543460845947,-26.5566673278809,
42.8012237548828,9.60439205169678,
14.9194202423096,29.9523105621338,
-16.6702651977539,34.6003799438477,
-2.38343882560730,34.5363578796387,
33.8004264831543,41.1133499145508,
32.0558662414551,51.8761253356934,
-17.0521316528320,58.8330154418945,
-55.1553230285645,49.7782974243164,
-35.2675476074219,17.9935989379883,
22.4424076080322,-26.9103488922119,
53.1164016723633,-54.9699821472168,
28.2576560974121,-43.0546302795410,
-19.8509025573730,-2.57342147827148,
-36.8748893737793,25.0641136169434,
-10.9957180023193,11.5048809051514,
26.5198173522949,-25.2040176391602,
39.7168388366699,-35.4759750366211,
25.3549652099609,2.99592256546021,
6.63754463195801,53.2641716003418,
2.32116174697876,65.9719085693359,
-2.30470371246338,32.6972236633301,
-27.6177501678467,-7.83026313781738,
-62.9818916320801,-23.7743968963623,
-71.4768905639648,-21.4119720458984,
-41.3213195800781,-25.6917934417725,
-0.903756916522980,-35.0915603637695,
14.1350536346436,-32.2222213745117,
2.18133330345154,-11.6783657073975,
-3.05378317832947,1.89835739135742,
16.3622245788574,-8.23188877105713,
40.6032066345215,-23.6624832153320,
43.1597518920898,-13.3766136169434,
31.6283798217773,27.8826560974121,
26.9155845642090,66.5740509033203,
33.1805152893066,67.1374816894531,
30.9896850585938,31.4737243652344,
17.7087936401367,-3.02883887290955,
13.3773984909058,-15.4520425796509,
27.8192310333252,-9.20067691802979,
41.5433502197266,-0.300626456737518,
24.5467777252197,9.80021381378174,
-13.1764888763428,27.6553249359131,
-37.6765480041504,37.8998451232910,
-30.8246307373047,19.6738605499268,
-6.47622585296631,-22.5365848541260,
17.6828441619873,-49.8941116333008,
42.1377067565918,-35.9836463928223,
62.6155281066895,-1.10060286521912,
59.7709503173828,18.4121532440186,
32.6348571777344,18.0862388610840,
9.47396659851074,26.3458290100098,
12.9959316253662,56.8718948364258,
23.6100807189941,79.3174057006836,
-0.0658786296844482,65.7066955566406,
-54.3969268798828,22.4420204162598,
-84.9182510375977,-20.9054965972900,
-54.5454025268555,-42.7425079345703,
11.9387941360474,-47.9082527160645,
55.9666442871094,-45.6204986572266,
56.0726585388184,-38.2767601013184,
24.9244651794434,-28.4745388031006,
-13.7045745849609,-21.1033649444580,
-36.1064338684082,-19.5534801483154,
-21.8202896118164,-20.9348621368408,
25.6490859985352,-25.4592552185059,
66.2148437500000,-33.2313346862793,
51.2458724975586,-27.0702438354492,
-9.56179332733154,2.51223468780518,
-61.3919563293457,32.2970962524414,
-62.4867706298828,26.0984153747559,
-32.7644195556641,-17.9309692382813,
-8.76580905914307,-57.4665679931641,
12.9947080612183,-52.1781616210938,
48.8501052856445,-20.0623970031738,
78.7640686035156,-3.88219451904297,
76.0434112548828,-10.6918907165527,
47.7974891662598,-10.0149946212769,
29.2750549316406,8.91064453125000,
30.9964122772217,16.3475494384766,
22.4587097167969,-0.914060950279236,
-13.7738399505615,-11.8864765167236,
-43.6394996643066,10.1521739959717,
-41.9024467468262,39.4106216430664,
-31.6908054351807,30.3613586425781,
-43.8179626464844,-16.3110160827637,
-57.4434242248535,-47.7870368957520,
-23.5731048583984,-35.2699394226074,
41.8704261779785,1.24926984310150,
66.9550857543945,26.7906932830811,
17.6394367218018,39.9474029541016,
-44.6931800842285,52.4965820312500,
-49.4470977783203,54.5207519531250,
-13.8061504364014,34.5251350402832,
-8.37450790405273,7.07043313980103,
-51.8283691406250,-0.410608470439911,
-76.4263076782227,5.21746349334717,
-30.4279365539551,-2.97310018539429,
46.4532508850098,-26.8867568969727,
74.1101150512695,-39.5907554626465,
34.6983718872070,-21.1474323272705,
-12.1959123611450,13.4921455383301,
-16.2952289581299,36.8081359863281,
8.80656909942627,41.8748741149902,
15.5502767562866,42.2440948486328,
-9.12794017791748,42.7557220458984,
-39.3697319030762,38.4012565612793,
-43.8393020629883,32.9370956420898,
-28.6525096893311,18.4456062316895,
-13.1915569305420,-15.6416921615601,
-7.23132276535034,-59.0759696960449,
-11.6806030273438,-67.6720886230469,
-20.4253253936768,-21.7813720703125,
-25.9646167755127,34.2538108825684,
-15.6153688430786,40.5055503845215,
11.1985445022583,-0.569127321243286,
37.0577812194824,-24.6920204162598,
37.9004516601563,-0.867484092712402,
10.4172105789185,25.4141998291016,
-13.6829338073730,3.53608393669128,
-13.2190980911255,-32.5708923339844,
7.27627038955689,-17.4482460021973,
25.9869174957275,41.3976440429688,
33.7624320983887,71.1232223510742,
32.9939765930176,43.5876846313477,
24.6803989410400,7.96178531646729,
2.92811489105225,6.35434532165527,
-22.6609554290772,13.2457656860352,
-31.2276096343994,-14.3163824081421,
-12.2443218231201,-53.7867050170898,
17.7721138000488,-50.9877853393555,
36.0497512817383,1.23890495300293,
33.0932655334473,46.8205909729004,
15.9919233322144,51.4863243103027,
-10.1455974578857,40.1664009094238,
-41.7866249084473,37.0418815612793,
-65.0915145874023,33.6576919555664,
-64.9176025390625,20.7289524078369,
-43.3273696899414,17.3526859283447,
-16.1619033813477,32.3438987731934,
-3.46780681610107,29.2196369171143,
-7.09573650360107,-15.4589204788208,
-15.9804687500000,-63.3178939819336,
-18.5797920227051,-58.1110153198242,
-15.0459232330322,-10.9147481918335,
-13.3237380981445,2.24960064888001,
-17.1518344879150,-44.7018928527832,
-22.6529331207275,-83.2674942016602,
-18.8218612670898,-46.3689270019531,
-7.08902168273926,24.8501777648926,
-2.56875395774841,40.5322761535645,
-11.4586162567139,-15.8579330444336,
-14.3681859970093,-71.9316329956055,
10.1475276947021,-59.7132873535156,
51.6000289916992,1.37962460517883,
69.9523315429688,46.9363403320313,
46.4603500366211,41.8782310485840,
6.24859905242920,2.21608328819275,
-11.3927202224731,-42.2581291198731,
-3.59660768508911,-69.8149490356445,
1.77163136005402,-69.2238311767578,
-9.92757415771484,-39.4571609497070,
-23.0558795928955,-10.9990348815918,
-22.3587703704834,-10.6689119338989,
-20.3414192199707,-28.3338947296143,
-31.3411254882813,-28.0567436218262,
-46.3536224365234,0.415618896484375,
-39.6532096862793,37.7064361572266,
-6.85530948638916,53.8192863464356,
21.4210128784180,41.7391510009766,
20.1688690185547,16.8034687042236,
-5.16883850097656,-5.19914913177490,
-27.3183040618897,-14.7640600204468,
-28.9195156097412,-4.45785045623779,
-14.1728191375732,16.0697097778320,
1.60679244995117,13.6263246536255,
12.1241474151611,-20.1346263885498,
16.6260337829590,-52.2805633544922,
9.48910713195801,-41.0261077880859,
-9.13041210174561,-2.45353126525879,
-31.6647682189941,9.88760185241699,
-37.2822723388672,-21.7703151702881,
-7.14125585556030,-56.8305168151856,
50.4293365478516,-47.8208694458008,
93.0959854125977,-4.68672657012939,
77.9139480590820,25.8469905853272,
11.5845518112183,25.8043613433838,
-50.3969917297363,16.5042781829834,
-57.9435882568359,5.31715202331543,
-18.6904277801514,-18.8889007568359,
15.9095287322998,-50.4526290893555,
18.5284080505371,-59.5988769531250,
16.0982589721680,-35.2690391540527,
39.4016304016113,-10.0470409393311,
73.3031234741211,-13.2750854492188,
76.4316177368164,-19.0982646942139,
46.7369461059570,13.5722494125366,
19.8106479644775,71.1634292602539,
19.6803531646729,92.6378936767578,
30.5321922302246,49.4671936035156,
24.9760475158691,-7.94402027130127,
9.46167087554932,-16.7937355041504,
2.35997438430786,15.2661190032959,
2.15039682388306,37.6647720336914,
-1.37600541114807,28.0574150085449,
-8.35637283325195,16.2306041717529,
-5.60599851608276,25.2857570648193,
4.84867429733276,37.3777084350586,
3.22026324272156,20.9695892333984,
-8.29685401916504,-13.5695152282715,
-3.34137368202209,-29.6452178955078,
25.5346202850342,-9.39649868011475,
51.6566848754883,24.6090087890625,
46.9182319641113,43.0347709655762,
13.2181653976440,44.2922210693359,
-26.5630950927734,38.0771713256836,
-55.9961242675781,22.3360099792480,
-68.3162612915039,-7.53888845443726,
-56.5408401489258,-42.9260635375977,
-17.1203308105469,-57.1820449829102,
23.7039756774902,-32.3953208923340,
33.7885322570801,20.9228343963623,
14.0812778472900,67.5395202636719,
-1.53854656219482,84.2791900634766,
2.95448398590088,71.6794967651367,
7.67477941513062,45.0917968750000,
-6.16110515594482,18.9741325378418,
-24.2265930175781,-2.54448890686035,
-26.3956470489502,-21.6879062652588,
-21.5100593566895,-36.1659049987793,
-28.9949645996094,-39.3627357482910,
-43.4891242980957,-33.4401054382324,
-32.7635917663574,-26.8532390594482,
7.53988361358643,-24.1437568664551,
41.9019660949707,-11.0089216232300,
43.2143821716309,18.4248676300049,
24.8896522521973,48.5476646423340,
20.4006729125977,52.4250221252441,
26.8136539459229,25.4370555877686,
23.4967651367188,1.74373543262482,
7.66692209243774,11.7507209777832,
-6.32061815261841,41.2595062255859,
-10.4387140274048,51.9930343627930,
-12.3054018020630,31.7405605316162,
-13.3454523086548,8.14754486083984,
1.50153958797455,-0.163269668817520,
33.8162002563477,-1.50028288364410,
56.7928695678711,-6.68602323532105,
51.4489402770996,-0.502208113670349,
32.2283744812012,28.9556808471680,
23.4773979187012,60.7103729248047,
10.3785209655762,56.7792778015137,
-30.6817512512207,22.9510059356689,
-74.4748916625977,-0.211496055126190,
-72.2754287719727,3.74427556991577,
-12.6526832580566,6.37322235107422,
48.8120689392090,-11.8287220001221,
62.1914100646973,-21.6510505676270,
40.3813095092773,6.13683128356934,
29.1585884094238,45.8119697570801,
35.6773872375488,45.0609703063965,
29.1414337158203,2.71118378639221,
1.25941383838654,-31.4190444946289,
-22.5852146148682,-26.7871723175049,
-32.7308082580566,-12.0618305206299,
-45.0106239318848,-23.3265743255615,
-55.5660552978516,-47.0531883239746,
-34.6681327819824,-45.9322204589844,
22.7181015014648,-22.6036415100098,
70.9650573730469,-13.3200120925903,
67.1090698242188,-29.4805088043213,
28.5876960754395,-44.0159759521484,
3.68593573570251,-31.3762397766113,
7.64595031738281,-4.99209308624268,
12.7438945770264,10.4825086593628,
9.61094951629639,12.2911157608032,
17.2440376281738,12.3613262176514,
29.7802257537842,16.1570091247559,
15.5727310180664,16.6148910522461,
-28.4671268463135,11.5359516143799,
-46.3681907653809,10.9702587127686,
-5.96977853775024,11.9939384460449,
50.4538269042969,-2.40038776397705,
56.1254730224609,-32.7659568786621,
10.4015560150146,-57.2550659179688,
-23.8027267456055,-51.9456443786621,
-6.90199756622314,-14.7471408843994,
27.3702163696289,30.2073421478272,
24.0046520233154,52.9859542846680,
-10.8050775527954,37.2328491210938,
-36.9448280334473,-3.33277964591980,
-34.5194702148438,-39.6710319519043,
-15.2536954879761,-44.8350639343262,
3.36542892456055,-19.7356529235840,
2.79818916320801,1.84159612655640,
-25.9832420349121,-4.44964981079102,
-65.5862960815430,-24.1293334960938,
-74.4863433837891,-20.9271011352539,
-36.7450180053711,9.10036468505859,
7.00925350189209,33.0641746520996,
5.14066028594971,28.9858932495117,
-29.8429584503174,13.5175952911377,
-29.6179332733154,10.6813459396362,
25.7757110595703,13.7666263580322,
66.4980850219727,-2.76654815673828,
37.0112380981445,-33.1954116821289,
-15.7538614273071,-38.0294151306152,
-14.5353908538818,-5.17722177505493,
31.5332336425781,33.6699371337891,
52.8636665344238,43.8278808593750,
29.7284450531006,28.9451332092285,
18.6508216857910,15.1025600433350,
48.7541618347168,3.71602344512939,
63.5372276306152,-12.4725303649902,
13.8114166259766,-19.0573177337647,
-46.7165298461914,0.375976949930191,
-38.1360969543457,28.9508762359619,
24.2045001983643,27.8445510864258,
51.3150482177734,-8.35375499725342,
20.7930202484131,-36.2655563354492,
-2.55701613426209,-19.1433258056641,
15.6981039047241,19.2822036743164,
20.2081146240234,35.5903549194336,
-24.1589622497559,21.3930053710938,
-64.4067001342773,-0.694564402103424,
-30.1666793823242,-20.6320838928223,
41.4106330871582,-36.3842849731445,
52.2671203613281,-33.9838180541992,
-18.9250431060791,-8.74478149414063,
-79.8309783935547,15.0782279968262,
-64.0839309692383,-0.352548837661743,
-13.4644641876221,-41.7296142578125,
-0.0701367259025574,-54.8621597290039,
-19.2510547637939,-16.3212299346924,
-19.4416866302490,22.8334064483643,
10.2640085220337,10.1504468917847,
37.8156509399414,-34.0436820983887,
44.0976142883301,-48.0936470031738,
47.4632644653320,-21.8328723907471,
61.6908912658691,-0.664276957511902,
74.5957107543945,-10.0935678482056,
70.9998474121094,-22.4965744018555,
63.0196876525879,-1.87112581729889,
61.5259666442871,37.5756301879883,
47.9428520202637,63.0115165710449,
6.65665245056152,64.2267303466797,
-39.9505195617676,52.0787925720215,
-62.4370079040527,27.7150173187256,
-59.7002143859863,-16.2625732421875,
-44.6922264099121,-62.8556709289551,
-25.3505058288574,-73.9841461181641,
2.37265110015869,-38.0372543334961,
28.4738292694092,5.21545124053955,
35.9728622436523,18.8436336517334,
27.4073619842529,4.52470827102661,
29.1271858215332,-9.51395893096924,
49.7724723815918,-2.55609893798828,
60.5368423461914,28.1374950408936,
35.6947822570801,65.6130218505859,
1.54880475997925,88.3232269287109,
-3.13569617271423,75.4457015991211,
19.9587745666504,32.2059020996094,
28.5816497802734,-6.21908283233643,
3.53883457183838,-7.33669376373291,
-29.8582592010498,14.9074172973633,
-38.8492164611816,23.4567565917969,
-20.5789051055908,10.0213155746460,
0.935225784778595,8.57304859161377,
16.0574512481689,32.9651947021484,
23.9183692932129,49.2379646301270,
21.7979087829590,29.3355121612549,
5.53317356109619,-3.48214149475098,
-8.39863204956055,-1.03310894966125,
-1.57472109794617,41.5629081726074,
13.0199632644653,76.2360916137695,
6.98388862609863,68.4119110107422,
-15.9971294403076,36.1849288940430,
-28.5141429901123,5.38399505615234,
-15.8592271804810,-17.7295818328857,
0.521088123321533,-34.2414512634277,
-0.0569618195295334,-24.8952960968018,
-5.88029718399048,16.7258834838867,
5.23761129379273,50.3573989868164,
20.7470455169678,31.3165893554688,
15.8117446899414,-22.0502872467041,
4.86928415298462,-50.3071441650391,
20.8078899383545,-27.5972709655762,
54.9598464965820,3.68621611595154,
54.7796211242676,0.586363911628723,
4.65918540954590,-21.4568614959717,
-37.4122657775879,-16.7607975006104,
-15.3486003875732,17.0176239013672,
43.4361801147461,36.1384162902832,
63.6329650878906,22.0634269714355,
24.5226669311523,-7.26332950592041,
-16.1023864746094,-27.5776424407959,
-2.76364064216614,-31.1400356292725,
40.3337135314941,-20.4034824371338,
51.5564727783203,9.76149368286133,
15.3306045532227,48.7161445617676,
-30.5207595825195,64.3996429443359,
-49.2366714477539,42.0946464538574,
-33.3296241760254,6.65744256973267,
0.129644870758057,-6.18919467926025,
29.0565338134766,3.29313135147095,
34.3527374267578,4.41351890563965,
17.4046134948730,-2.98316836357117,
1.70843636989594,8.43951988220215,
1.33587145805359,42.2659149169922,
3.18654394149780,54.5347747802734,
-15.3536262512207,12.6137952804565,
-41.1263427734375,-55.9258041381836,
-30.8247337341309,-82.5455093383789,
14.5666065216064,-44.1969146728516,
36.8136672973633,14.0560340881348,
3.20866203308105,36.4200172424316,
-40.5595512390137,14.7916393280029,
-28.2381191253662,-16.9829406738281,
35.9289283752441,-28.7209701538086,
83.2856292724609,-19.7878513336182,
73.2994918823242,1.93959522247314,
42.4992256164551,27.8637714385986,
30.6403560638428,45.3227958679199,
24.9244937896729,41.1267318725586,
-3.36368203163147,17.9534263610840,
-38.8756332397461,0.813579559326172,
-36.4141120910645,12.0824670791626,
3.97545194625855,41.0795135498047,
29.7842941284180,56.6894378662109,
5.26684236526489,41.5004882812500,
-37.6228637695313,16.6366214752197,
-51.9654006958008,6.71612405776978,
-31.2263889312744,12.9759492874146,
-10.5078983306885,12.1191663742065,
-17.8789577484131,-3.81358051300049,
-39.4615898132324,-14.6214323043823,
-45.0386581420898,-3.14765596389771,
-24.6568794250488,17.3592033386230,
0.806733012199402,26.1106586456299,
10.5521535873413,20.9952831268311,
0.805975079536438,14.1640567779541,
-10.4665470123291,9.57178115844727,
-10.7275648117065,-6.12140226364136,
-5.78306341171265,-27.5065975189209,
-10.8294458389282,-32.1001319885254,
-32.4151802062988,-13.7620172500610,
-53.6878318786621,2.17627286911011,
-53.2740707397461,-9.81958866119385,
-27.9660282135010,-34.1255455017090,
14.3375673294067,-39.4996604919434,
50.4756317138672,-23.7794399261475,
59.9094734191895,-11.9858236312866,
37.8012886047363,-13.6878376007080,
6.73728895187378,-7.08746480941773,
-5.24941110610962,15.6915607452393,
6.73945856094360,27.4374008178711,
16.6458740234375,2.03072071075439,
3.86174488067627,-40.5153732299805,
-11.5546360015869,-54.6108016967773,
0.358607649803162,-29.1455993652344,
34.8644828796387,2.55061626434326,
44.8378448486328,7.26869583129883,
1.00171566009521,-4.33744716644287,
-63.1102256774902,-2.91664814949036,
-87.3131713867188,9.25743865966797,
-55.9023704528809,9.55010700225830,
-8.10692405700684,-12.8787069320679,
7.19394397735596,-41.5716171264648,
-9.78320503234863,-48.8404464721680,
-15.3239841461182,-35.4019012451172,
10.9256820678711,-17.3835964202881,
48.9323463439941,-2.00070333480835,
62.5287628173828,21.6479740142822,
39.6539039611816,55.9336585998535,
-1.92983317375183,72.6170883178711,
-38.2712631225586,44.6091613769531,
-54.9671134948731,-16.7329978942871,
-42.9705009460449,-58.5589103698731,
-5.73368453979492,-36.3727874755859,
29.9254550933838,26.8252716064453,
25.0886249542236,67.9287261962891,
-17.0969181060791,48.3890647888184,
-50.1401977539063,-7.43256378173828,
-25.2783451080322,-49.7799873352051,
34.9358177185059,-55.3866729736328,
64.4293365478516,-39.2874832153320,
31.9897994995117,-20.1501293182373,
-20.0429801940918,2.35197210311890,
-31.2966995239258,24.9309787750244,
0.725360274314880,35.4952125549316,
30.4878387451172,21.5955486297607,
27.9531822204590,-9.60688018798828,
11.0513877868652,-32.6200752258301,
-0.215358436107636,-23.8646049499512,
-10.4886894226074,14.4126720428467,
-30.9796581268311,51.0581970214844,
-50.3114013671875,52.6389503479004,
-49.3391494750977,22.4679718017578,
-35.8738670349121,-2.43635106086731,
-34.3234710693359,10.0336704254150,
-44.0872993469238,40.2414627075195,
-35.9157638549805,37.4720458984375,
0.0160169601440430,-4.50878286361694,
33.9134674072266,-38.1134033203125,
29.6567420959473,-27.1178970336914,
-1.70741486549377,-5.45283126831055,
-16.4835968017578,-18.4631633758545,
0.165848478674889,-53.7135200500488,
15.5457048416138,-53.1489028930664,
2.09340643882751,0.274763107299805,
-30.4362983703613,51.8922691345215,
-47.6738014221191,51.8422698974609,
-39.0844573974609,21.7955036163330,
-25.2191410064697,5.73745679855347,
-20.2675189971924,1.03747713565826,
-10.9322738647461,-19.5015964508057,
19.6493186950684,-46.0179901123047,
54.1099166870117,-36.0983505249023,
57.8493156433106,4.61837625503540,
17.6184082031250,15.7073144912720,
-33.1403541564941,-32.5234832763672,
-41.6236114501953,-88.4426345825195,
11.2023086547852,-86.8347702026367,
75.8296966552734,-31.9668502807617,
86.9087142944336,15.0030975341797,
33.8165321350098,21.6454601287842,
-28.6749572753906,13.8129730224609,
-39.4001693725586,20.6069507598877,
-4.44173049926758,27.8350276947022,
18.3119239807129,17.2804203033447,
-0.218071579933167,-0.105387777090073,
-23.5410575866699,-6.05219841003418,
-6.99898099899292,-5.22274303436279,
34.9780883789063,-14.1137733459473,
51.2721672058106,-28.5113353729248,
29.8252944946289,-33.8868064880371,
11.9000797271729,-25.1577835083008,
32.7608032226563,-13.5226535797119,
64.0479202270508,-2.97957539558411,
52.1530113220215,12.1930332183838,
-7.31526947021484,33.5951347351074,
-62.5025062561035,41.3556289672852,
-68.6943817138672,31.2290058135986,
-32.7997207641602,23.7940940856934,
0.537529349327087,33.4148216247559,
3.25192475318909,50.1270599365234,
-16.1800060272217,52.3923454284668,
-37.0449981689453,37.8325462341309,
-46.7760086059570,17.2619228363037,
-44.4727630615234,-1.80315732955933,
-31.1835842132568,-19.2120208740234,
-13.4754343032837,-30.5450801849365,
1.18455123901367,-27.4662265777588,
10.0507335662842,-16.6735668182373,
15.0738487243652,-16.5787277221680,
18.4228076934814,-30.0386829376221,
12.6102209091187,-33.0523719787598,
-8.25463294982910,-7.91760540008545,
-32.3966636657715,29.6913776397705,
-37.9995384216309,44.9353141784668,
-22.6870708465576,25.5015258789063,
-5.21052312850952,-8.33628845214844,
-5.29655647277832,-29.7886524200439,
-13.6715679168701,-32.4914131164551,
-3.31512212753296,-21.8169040679932,
25.7647323608398,-7.85160064697266,
44.6073913574219,4.86766958236694,
33.3630447387695,13.3345918655396,
5.07743740081787,15.0324916839600,
-15.6914453506470,12.5731182098389,
-25.4896869659424,15.5332603454590,
-35.4343948364258,24.3356342315674,
-48.1920127868652,31.7787837982178,
-50.6491241455078,26.9560031890869,
-37.7999458312988,2.86003494262695,
-19.1436824798584,-31.3823471069336,
0.373521089553833,-47.2202568054199,
22.6247940063477,-24.6657085418701,
39.1098709106445,15.3798980712891,
27.8193416595459,31.6751289367676,
-8.14142990112305,10.3284797668457,
-36.3467445373535,-11.9855976104736,
-33.8189582824707,7.87943935394287,
-21.6825847625732,50.7595558166504,
-28.2935218811035,53.4038162231445,
-42.0386657714844,-7.29434156417847,
-28.8071174621582,-70.9202041625977,
11.5836944580078,-64.4851150512695,
31.6065158843994,0.784429430961609,
8.73126125335693,46.2520484924316,
-24.0972499847412,30.4890041351318,
-21.1394042968750,-7.90418195724487,
4.48886823654175,-13.9603128433228,
10.8161439895630,11.1420736312866,
-12.9027881622314,19.6842346191406,
-38.4867286682129,0.124564051628113,
-41.6216468811035,-15.2497425079346,
-36.7154426574707,-3.97473025321960,
-34.7796592712402,15.5065183639526,
-23.3650321960449,21.3324165344238,
4.46589183807373,18.3871135711670,
28.8784885406494,16.7654037475586,
20.2754077911377,8.74419784545898,
-18.7770309448242,-11.4022340774536,
-54.5687370300293,-20.1844539642334,
-60.2036476135254,3.06997108459473,
-48.0730438232422,26.5194339752197,
-42.0032043457031,4.52837896347046,
-39.1693038940430,-55.8986625671387,
-15.9259490966797,-85.6134948730469,
38.5208892822266,-49.6920585632324,
91.0993728637695,-0.952967286109924,
90.3383331298828,-1.40527403354645,
30.1457157135010,-33.4286079406738,
-31.1133956909180,-31.9760818481445,
-37.9613838195801,13.0330429077148,
-1.62749552726746,40.1375083923340,
14.0319089889526,12.7841749191284,
-10.6997165679932,-24.1874675750732,
-31.9232234954834,-12.8902750015259,
-10.2842445373535,34.0098533630371,
25.3426628112793,55.1529426574707,
19.2154598236084,34.5831604003906,
-26.5606727600098,14.3910665512085,
-53.8585052490234,18.1412353515625,
-33.9743576049805,19.7654342651367,
0.128064334392548,-4.53624439239502,
14.6056404113770,-31.6196804046631,
14.0566930770874,-31.0772628784180,
11.3111534118652,-0.0121986865997314,
-1.88015604019165,27.7561855316162,
-35.5421829223633,26.5432033538818,
-51.2216682434082,-3.25848674774170,
-10.9239559173584,-42.6141242980957,
57.1180534362793,-64.4334945678711,
86.6772766113281,-40.4027137756348,
54.9819755554199,23.1523017883301,
7.22384595870972,68.7547760009766,
-6.31706523895264,44.3848991394043,
8.22032356262207,-22.5606288909912,
9.46678352355957,-50.4196510314941,
-10.7925338745117,-15.5651884078980,
-30.4303321838379,18.7013645172119,
-33.0212326049805,-7.76581382751465,
-19.5539169311523,-65.6879577636719,
9.87026214599609,-77.9927291870117,
41.1613121032715,-30.2271766662598,
46.8987922668457,11.0687131881714,
15.2650165557861,-1.55087077617645,
-18.9160766601563,-28.3535861968994,
-11.7353038787842,-17.0238857269287,
22.3091793060303,26.1019344329834,
28.3252754211426,52.2121238708496,
-12.0260400772095,36.6599540710449,
-45.2608489990234,6.46997165679932,
-14.1407871246338,-13.1717309951782,
50.7983589172363,-23.1650104522705,
81.2177047729492,-22.5074214935303,
64.2414474487305,-7.17530536651611,
49.3443603515625,14.8027305603027,
61.2560424804688,18.7266025543213,
69.8993682861328,-1.23634457588196,
46.9749946594238,-10.5121688842773,
15.0133514404297,27.8286781311035,
5.45565223693848,85.3321990966797,
3.27944207191467,97.9674453735352,
-18.2675571441650,43.4444122314453,
-50.2550735473633,-32.1710090637207,
-54.7701034545898,-64.9247283935547,
-25.8682785034180,-41.9053649902344,
-6.38145112991333,-5.86663818359375,
-21.9195270538330,0.408363938331604,
-46.1055755615234,-21.1372528076172,
-43.2017173767090,-40.9812736511231,
-20.4289588928223,-36.5005073547363,
-4.30185317993164,-14.2349328994751,
-4.53578805923462,0.983935713768005,
-10.0366497039795,-9.26413536071777,
-8.62192344665527,-34.2930107116699,
1.87942981719971,-43.3980407714844,
20.0875453948975,-17.8007869720459,
42.5576744079590,22.7392902374268,
45.8727340698242,45.5573005676270,
12.9812469482422,40.9755172729492,
-38.5916213989258,16.2592391967773,
-61.4963569641113,-11.2752952575684,
-33.7020187377930,-36.8469848632813,
9.92875480651856,-53.1795501708984,
28.5295944213867,-46.8970489501953,
21.6735382080078,-21.0347480773926,
21.9777069091797,-1.78506231307983,
40.2840995788574,-12.1776103973389,
51.4179306030273,-34.6147651672363,
31.8478603363037,-40.5945243835449,
-4.19955539703369,-28.4213790893555,
-17.6035976409912,-25.2906246185303,
2.86352014541626,-41.5468940734863,
36.1642570495606,-48.2766799926758,
56.1668891906738,-21.8435821533203,
51.9934844970703,24.5640144348145,
32.4791755676270,58.1516113281250,
6.49864339828491,66.7478256225586,
-14.6253118515015,61.3147659301758,
-22.5187435150147,47.3599319458008,
-17.4010791778564,20.6214332580566,
-8.45280742645264,-5.61267185211182,
-5.17407751083374,-2.92303657531738,
-6.67719173431397,31.5859718322754,
-10.2240591049194,59.1347541809082,
-22.6448535919189,48.9406547546387,
-49.9845199584961,13.6580972671509,
-76.8820877075195,-13.6528577804565,
-71.6693954467773,-21.5935611724854,
-24.9979915618897,-20.2384033203125,
28.1309947967529,-18.0897178649902,
47.9971237182617,-15.7305669784546,
30.7738170623779,-19.6536846160889,
16.1624164581299,-37.1270179748535,
29.2964820861816,-51.7339859008789,
52.2911605834961,-27.3698902130127,
45.4549446105957,28.0911407470703,
3.05303716659546,65.9822998046875,
-40.2680778503418,53.9266319274902,
-49.7644386291504,21.1293582916260,
-24.8420066833496,9.88672065734863,
7.47236347198486,17.9513454437256,
23.0239772796631,9.59488105773926,
23.9778213500977,-16.0307540893555,
27.1583461761475,-23.9983463287354,
41.0103225708008,-0.522726535797119,
55.6195755004883,18.6823215484619,
49.3064575195313,7.92495536804199,
26.1202239990234,-3.88159227371216,
6.38359546661377,20.9381713867188,
10.6777048110962,59.8914299011231,
31.0517768859863,60.4736251831055,
41.2066917419434,14.8512868881226,
28.3556041717529,-22.6850109100342,
10.4819993972778,-19.1469001770020,
1.18353581428528,-4.30098056793213,
-3.46356892585754,-19.2295284271240,
-12.8589668273926,-54.4341430664063,
-26.3853797912598,-61.8510437011719,
-35.3028869628906,-28.8643474578857,
-37.7322196960449,7.16004991531372,
-28.2868499755859,13.1528062820435,
4.40006637573242,2.27810859680176,
52.2444877624512,-3.07885336875916,
78.9448318481445,-4.82356166839600,
50.9964256286621,-13.9537696838379,
-6.48468542098999,-26.5059051513672,
-30.6981086730957,-29.6132087707520,
1.28718149662018,-22.3223342895508,
40.3680381774902,-16.2674446105957,
37.5156021118164,-18.1627368927002,
10.7289428710938,-20.1212406158447,
0.369325816631317,-14.5223026275635,
4.53605604171753,-5.33576250076294,
-6.07056999206543,9.43280315399170,
-26.8895359039307,28.3971729278564,
-22.6625652313232,33.5370712280273,
8.67696094512940,1.29515337944031,
20.6258125305176,-47.0153770446777,
-12.0752782821655,-58.7086753845215,
-41.2496299743652,-16.8654041290283,
-23.2355384826660,30.0333652496338,
10.3538265228271,28.0280971527100,
3.06473851203918,-12.6731777191162,
-33.3002624511719,-36.7873878479004,
-35.8651084899902,-22.6066226959229,
5.45761871337891,-9.59286117553711,
26.1202392578125,-26.4713134765625,
-6.47025728225708,-47.5183486938477,
-38.4054450988770,-41.1991577148438,
-4.54426956176758,-20.4466037750244,
69.3397750854492,-10.5655307769775,
99.7670288085938,-7.16788530349731,
64.3077011108398,5.77378129959106,
24.4948253631592,14.6513824462891,
28.4900760650635,-1.11999201774597,
45.8905677795410,-22.6640586853027,
30.8544521331787,-9.39107990264893,
-4.92049312591553,27.3241310119629,
-17.9053001403809,32.9668273925781,
3.17692518234253,-11.7001190185547,
28.8441677093506,-47.4869461059570,
38.8645820617676,-20.7887706756592,
36.4369239807129,31.4790706634522,
26.9212779998779,40.8908424377441,
5.97974777221680,3.91279792785645,
-19.2659835815430,-23.5430850982666,
-24.0196552276611,-19.3615665435791,
-2.34705877304077,-12.9734725952148,
14.9901285171509,-22.8341083526611,
3.66989755630493,-19.5010032653809,
-12.8497838973999,15.5648612976074,
-6.05611801147461,51.1105804443359,
15.9785976409912,47.4576263427734,
14.8796958923340,23.1535072326660,
-21.2172088623047,20.8213691711426,
-57.4420051574707,39.8651351928711,
-55.8433685302734,37.5890769958496,
-22.9347171783447,3.24880409240723,
5.77658748626709,-25.1309185028076,
13.3496570587158,-21.5723838806152,
8.79604244232178,-3.92331933975220,
6.90597391128540,2.21209526062012,
6.67826175689697,-3.17252755165100,
3.08294773101807,-5.72638463973999,
2.16482472419739,-10.1426391601563,
8.21128845214844,-28.9394550323486,
19.0436077117920,-44.2710494995117,
25.7507953643799,-28.1186027526855,
27.0148906707764,17.6066761016846,
29.5556697845459,53.3112182617188,
35.0382614135742,50.4487304687500,
33.7947235107422,26.5175457000732,
17.4729938507080,17.2659721374512,
-3.99071407318115,27.4572391510010,
-10.9054498672485,33.1953392028809,
1.89206981658936,21.1320266723633,
17.3349876403809,4.93032026290894,
12.7401485443115,8.12393665313721,
-10.4954729080200,25.1433582305908,
-34.1534957885742,23.8839702606201,
-42.6395034790039,-10.8570575714111,
-40.0827827453613,-50.4112663269043,
-34.3138656616211,-55.2953681945801,
-20.8395442962647,-23.3316440582275,
6.84723997116089,7.54911041259766,
37.6534271240234,11.8300542831421,
52.2712821960449,5.74578714370728,
41.8541526794434,23.3992881774902,
19.3474540710449,62.6005516052246,
-1.57158792018890,77.8882675170898,
-15.2363557815552,43.9767456054688,
-25.9665832519531,-9.86339092254639,
-25.2593803405762,-32.6967811584473,
-2.62656354904175,-14.3746557235718,
32.2797431945801,8.61515903472900,
50.4527816772461,3.59327626228333,
33.8938484191895,-16.2132587432861,
-0.869093179702759,-15.7010288238525,
-17.2093639373779,3.19997525215149,
-1.10547637939453,7.51498174667358,
22.4722805023193,-8.15713024139404,
23.4254264831543,-10.9723415374756,
7.70229768753052,24.9127006530762,
0.603668570518494,67.7147903442383,
4.55464839935303,65.7403640747070,
-3.98847532272339,20.8210582733154,
-35.2746887207031,-11.6312503814697,
-58.5924415588379,1.12951576709747,
-41.1603507995606,24.4841632843018,
-0.902451574802399,15.3363866806030,
12.8838281631470,-11.4787502288818,
-13.7997837066650,-9.52062225341797,
-33.7528533935547,21.7934741973877,
-7.47497272491455,36.2492485046387,
42.7515983581543,10.5047569274902,
58.8133926391602,-23.9413318634033,
27.0979404449463,-30.5219764709473,
-9.66504859924316,-15.8131704330444,
-15.8468799591064,-5.39065217971802,
-5.94712209701538,-6.83142089843750,
-9.48580837249756,-11.3815088272095,
-22.8167304992676,-21.1499462127686,
-21.3498077392578,-35.9081497192383,
2.04563593864441,-33.3560333251953,
23.5291671752930,10.6253261566162,
25.3888244628906,62.2657737731934,
16.1966972351074,61.6019515991211,
12.6261062622070,4.92802000045776,
13.8473682403564,-42.7128639221191,
12.2601480484009,-32.1691055297852,
8.95423507690430,7.42321300506592,
6.70413160324097,24.6129074096680,
8.33190917968750,17.4453258514404,
14.3159990310669,22.8686008453369,
11.5245914459229,43.7371253967285,
-11.6466932296753,37.9682655334473,
-47.3927650451660,1.09024822711945,
-66.3250122070313,-20.5680389404297,
-40.5155982971191,1.05998766422272,
14.2421607971191,24.4550838470459,
41.9343414306641,4.49618053436279,
16.9121208190918,-39.4281806945801,
-22.9003696441650,-45.7371215820313,
-26.3072376251221,-3.86949324607849,
-2.02399778366089,34.3135681152344,
1.32807362079620,35.0724487304688,
-26.3967895507813,18.7867889404297,
-36.6500549316406,17.1514205932617,
0.731602430343628,19.9767093658447,
44.6141433715820,-4.11238288879395,
32.4547729492188,-47.4847106933594,
-27.2872200012207,-69.7667846679688,
-63.1287841796875,-54.4229621887207,
-27.4222297668457,-31.7874965667725,
43.7728462219238,-30.4446048736572,
79.3795471191406,-37.7503471374512,
50.7713890075684,-24.4323139190674,
-4.27674531936646,9.94927787780762,
-37.7934608459473,32.5622863769531,
-33.0689849853516,16.6821498870850,
-9.15901565551758,-18.0017337799072,
8.19747257232666,-28.6689167022705,
5.79417657852173,-5.11623287200928,
-5.96846342086792,26.1207523345947,
-15.1443290710449,32.7504577636719,
-23.5665702819824,12.4343185424805,
-37.4131393432617,-6.62605571746826,
-53.5185165405273,-6.66063022613525,
-54.5823326110840,-2.22332954406738,
-31.9286937713623,-16.8828926086426,
0.167083382606506,-37.1229133605957,
10.1192731857300,-32.8359756469727,
-11.6199645996094,6.24928331375122,
-39.8136062622070,41.2491455078125,
-50.7108573913574,29.7050209045410,
-36.2241935729981,-20.2259559631348,
-3.45479393005371,-50.2779884338379,
33.6088905334473,-21.5752887725830,
58.9165458679199,35.4032821655273,
52.8292922973633,55.4635963439941,
14.1627769470215,23.6473045349121,
-30.3687686920166,-15.8805561065674,
-51.4061393737793,-19.9694004058838,
-49.3297576904297,0.289799153804779,
-52.1298522949219,1.28847503662109,
-58.7340583801270,-28.4293041229248,
-38.6528434753418,-54.8268737792969,
20.2912635803223,-49.0733184814453,
68.5837707519531,-21.4336357116699,
51.5551528930664,2.62478303909302,
-19.1713275909424,10.4322195053101,
-71.3159942626953,8.57561683654785,
-65.0058670043945,6.37370824813843,
-28.2657890319824,10.7721834182739,
-9.61257934570313,30.1909828186035,
-9.59004783630371,59.1427536010742,
-0.713068068027496,68.1324539184570,
10.9365139007568,37.4174499511719,
-2.34046697616577,-11.0442790985107,
-42.4835357666016,-31.9314136505127,
-67.6742172241211,-7.55404901504517,
-50.7528228759766,28.5205917358398,
-17.3877487182617,33.2227058410645,
-7.88623666763306,6.64486789703369,
-24.1137523651123,-18.2627029418945,
-41.9331245422363,-21.9623107910156,
-47.0948486328125,-12.9193429946899,
-42.2206382751465,-5.64351558685303,
-33.0199012756348,-1.85825979709625,
-13.3511743545532,1.81568646430969,
14.6469259262085,4.06090259552002,
26.5095863342285,3.85946083068848,
10.7796039581299,4.67227363586426,
-15.6388254165649,11.0904645919800,
-29.9243621826172,15.7716531753540,
-26.3112239837647,12.2495384216309,
-11.4346275329590,3.21925497055054,
3.31227207183838,0.641239881515503,
5.83593845367432,6.20000123977661,
-7.72408676147461,13.4224948883057,
-23.9216728210449,22.7184505462647,
-18.4305801391602,34.5604476928711,
10.8334722518921,36.1104469299316,
33.4764518737793,17.5166435241699,
19.6839523315430,-12.7947854995728,
-11.1682806015015,-21.9561252593994,
-17.5480079650879,5.07454204559326,
1.97030973434448,41.2238235473633,
3.94664192199707,48.8980941772461,
-26.3658142089844,27.2843952178955,
-43.9099197387695,8.72060871124268,
-13.3949508666992,9.97224998474121,
34.2307128906250,12.9277706146240,
37.0856094360352,1.44478321075439,
-7.10393190383911,-12.8995895385742,
-38.9517440795898,-12.9104394912720,
-25.6763534545898,-9.01303482055664,
-3.32017445564270,-24.9445285797119,
-9.80292415618897,-56.3779029846191,
-23.6097316741943,-71.5019912719727,
-7.13290882110596,-51.9575309753418,
26.8322792053223,-14.1632337570190,
30.0725402832031,8.45061492919922,
-0.383213609457016,7.59946584701538,
-14.4052486419678,2.65263605117798,
13.4341030120850,9.28750228881836,
44.0671882629395,26.4225101470947,
31.7449111938477,46.6882667541504,
-12.1165895462036,53.9763717651367,
-37.0188217163086,45.7622985839844,
-27.7526378631592,30.3636760711670,
-14.8796596527100,20.0376605987549,
-20.9854316711426,11.8620109558105,
-23.3033943176270,-6.09658813476563,
1.73977613449097,-29.3308849334717,
38.4946250915527,-29.2417793273926,
49.8305778503418,4.89063787460327,
24.6263980865479,41.2188873291016,
-8.92910480499268,31.7042846679688,
-19.1412048339844,-16.5321388244629,
-4.41939115524292,-39.5911254882813,
16.6398983001709,1.64769792556763,
25.8133010864258,68.3438873291016,
14.7321739196777,89.7076034545898,
-15.0654249191284,49.4100761413574,
-51.5242080688477,-5.46965551376343,
-67.7438583374023,-28.7635612487793,
-51.5032615661621,-19.1696014404297,
-23.4014644622803,-3.23144555091858,
-14.4207239151001,-1.11966311931610,
-27.0347881317139,-13.3331060409546,
-33.6848869323731,-31.5316734313965,
-12.1813716888428,-37.9766273498535,
19.5617046356201,-16.4656753540039,
19.1941471099854,20.5887393951416,
-20.3176250457764,38.3775711059570,
-57.7698135375977,23.4724483489990,
-51.1336059570313,7.20090341567993,
-2.80135297775269,12.4253759384155,
44.2155456542969,14.6702146530151,
51.4212036132813,-15.2403316497803,
26.9906177520752,-52.8557662963867,
10.0286188125610,-43.2104187011719,
21.8740921020508,19.9049568176270,
36.2407341003418,64.7305374145508,
12.8351974487305,38.0570793151856,
-43.1299476623535,-16.4304103851318,
-77.3075790405273,-21.8934288024902,
-50.0178070068359,23.6333503723145,
8.73080253601074,51.0631103515625,
30.4457778930664,23.9093093872070,
-5.00772857666016,-8.25060653686523,
-40.4050598144531,7.89122104644775,
-23.4785556793213,42.0846290588379,
23.0735969543457,33.0204315185547,
38.9052696228027,-19.5797367095947,
10.8407220840454,-52.7195053100586,
-9.96706485748291,-29.0616683959961,
19.0116119384766,10.3089752197266,
68.9310760498047,5.86214733123779,
84.0095214843750,-32.3662796020508,
47.6716499328613,-43.6146926879883,
-4.44355535507202,-7.86352109909058,
-36.9225997924805,29.1780891418457,
-43.5251617431641,16.8801307678223,
-35.9921760559082,-37.0874061584473,
-21.1790084838867,-71.9688186645508,
-2.48796129226685,-40.1619567871094,
9.67131233215332,32.0425834655762,
12.3488960266113,68.8193817138672,
12.5540390014648,28.7621555328369,
19.2781963348389,-45.8265113830566,
27.2111949920654,-69.3345870971680,
26.1638736724854,-9.03726196289063,
17.4583988189697,69.5876846313477,
13.7551326751709,75.5674667358398,
19.2346439361572,9.97665691375732,
21.7617683410645,-46.1020965576172,
10.5588741302490,-33.2701644897461,
-2.36425662040710,15.2474184036255,
-6.13985395431519,35.3516540527344,
-6.14951848983765,18.8870849609375,
-15.6454334259033,8.92061519622803,
-30.8815860748291,24.9162864685059,
-28.2292442321777,35.5170555114746,
4.03634405136108,11.5597953796387,
45.9226608276367,-20.6124477386475,
58.7320137023926,-24.1693420410156,
30.7062416076660,-4.67186784744263,
-12.5273532867432,-1.43793296813965,
-32.3240661621094,-28.2232189178467,
-21.5109920501709,-59.3384666442871,
0.328940749168396,-70.2790298461914,
9.56251621246338,-58.3281745910645,
6.34433841705322,-30.2941894531250,
12.9597616195679,-1.73746681213379,
39.7353897094727,7.90590858459473,
59.2657470703125,-9.29926681518555,
38.8357086181641,-32.1564750671387,
-11.3164482116699,-18.1588325500488,
-40.3574829101563,33.5140953063965,
-19.7955322265625,63.0107078552246,
20.2588272094727,28.5190849304199,
32.8391990661621,-30.3317794799805,
18.5408020019531,-33.3259010314941,
24.6128330230713,20.6212501525879,
54.6401176452637,51.9362106323242,
61.5974769592285,13.2622337341309,
16.8242683410645,-40.2139358520508,
-34.2125396728516,-31.6906452178955,
-35.6171760559082,25.9446887969971,
-1.97815930843353,43.5439987182617,
6.60712003707886,-6.13722562789917,
-20.9592838287354,-53.2043685913086,
-37.8584671020508,-28.9508323669434,
-18.2404747009277,37.0229568481445,
-0.722743391990662,62.2040023803711,
-17.0100593566895,19.3559589385986,
-41.3470916748047,-40.1958236694336,
-24.3282890319824,-63.2067413330078,
28.6336517333984,-49.2724189758301,
64.8533096313477,-23.3172187805176,
65.7601776123047,-0.0855447649955750,
56.3749046325684,13.6419057846069,
54.2944412231445,10.6919689178467,
46.1744117736816,-10.7010354995728,
26.1597919464111,-31.0646800994873,
11.3567771911621,-25.9781455993652,
13.6966381072998,-6.40841150283814,
17.9712810516357,2.82544398307800,
9.05041694641113,-1.10085105895996,
-6.02512884140015,0.740889549255371,
-16.2432384490967,15.5936422348022,
-28.7476234436035,26.6889839172363,
-54.2549896240234,13.8887214660645,
-65.7989120483398,-13.3447999954224,
-30.1201095581055,-21.4760494232178,
35.0054855346680,-1.07951140403748,
68.9002609252930,25.5559978485107,
46.4839210510254,33.2225074768066,
-0.295491933822632,13.8463973999023,
-24.8814449310303,-21.2003440856934,
-15.0237617492676,-53.6480064392090,
15.1752805709839,-65.9135055541992,
44.0334396362305,-50.7516555786133,
54.1649513244629,-19.8462657928467,
34.6824569702148,0.586017131805420,
-0.479624748229980,-5.57769393920898,
-7.91200399398804,-19.4794063568115,
33.5207328796387,-16.5374050140381,
78.3468017578125,0.516895949840546,
64.8260498046875,3.78425645828247,
6.32731628417969,-18.6218395233154,
-23.7547988891602,-37.6430740356445,
10.0180711746216,-27.1504478454590,
49.8950080871582,-5.01541280746460,
36.0029716491699,-2.80339288711548,
-7.74196720123291,-22.0032501220703,
-18.5724964141846,-27.4731082916260,
11.8551120758057,4.49675512313843,
23.6320266723633,41.1072654724121,
-14.0596103668213,36.4147949218750,
-52.3901252746582,-14.6060400009155,
-41.2597503662109,-66.1480789184570,
-0.772049188613892,-71.3432540893555,
9.70295333862305,-30.6982822418213,
-18.7028522491455,14.6072521209717,
-44.3091049194336,21.7065391540527,
-39.5948219299316,-11.8848991394043,
-15.6331663131714,-42.0282249450684,
7.81672573089600,-22.5401325225830,
19.7171993255615,36.9278488159180,
13.7035188674927,77.9633178710938,
-10.5581436157227,53.9330711364746,
-33.5615653991699,-14.5972318649292,
-22.7598571777344,-58.9111824035645,
18.0011310577393,-41.4387817382813,
39.8780326843262,5.82782888412476,
19.0966014862061,37.4826393127441,
-3.78092956542969,48.0141448974609,
9.44464874267578,52.0593185424805,
29.4204177856445,48.9071083068848,
6.76309156417847,27.9107856750488,
-42.1828842163086,-4.51347780227661,
-50.4874382019043,-18.9424381256104,
-2.64602923393250,-12.6194686889648,
38.6811637878418,-18.8751792907715,
22.7810897827148,-54.5697860717773,
-10.2880697250366,-79.6852340698242,
4.32226467132568,-53.6769447326660,
53.2186241149902,1.11978507041931,
66.4587707519531,21.5766181945801,
26.3258743286133,-14.4681243896484,
-11.2717666625977,-47.5588531494141,
-5.91313171386719,-27.7865200042725,
19.5817413330078,19.7259330749512,
29.7991390228272,35.5217590332031,
23.7248897552490,5.83669662475586,
16.2317447662354,-20.9560871124268,
6.38103437423706,-16.6960773468018,
-13.1524438858032,-5.68087244033814,
-26.9675960540772,-23.0568618774414,
-17.9680747985840,-53.6940650939941,
-6.89355468750000,-53.9889144897461,
-22.4779453277588,-17.9540863037109,
-43.5655174255371,15.0184478759766,
-23.0647697448730,9.00189208984375,
28.7382621765137,-24.2296829223633,
44.6114044189453,-50.0650138854981,
-1.12457728385925,-42.5565261840820,
-45.8591194152832,-8.29400634765625,
-29.0646533966064,25.4871215820313,
17.7745475769043,39.5250892639160,
14.8784608840942,36.6330261230469,
-43.5757789611816,30.5135059356689,
-74.5965347290039,27.4470310211182,
-23.9864273071289,18.7201709747314,
54.6312522888184,1.37457227706909,
75.0676498413086,-10.9574851989746,
31.6315994262695,-0.951613664627075,
-8.40039825439453,26.7711982727051,
-5.90668439865112,48.9609222412109,
13.4427366256714,52.7648582458496,
12.9864873886108,43.3508720397949,
-1.66320312023163,26.1672744750977,
-2.51285743713379,4.44842767715454,
13.1774864196777,-11.5369215011597,
23.8546638488770,-9.35639286041260,
15.3445158004761,2.51494622230530,
-5.53080844879150,2.26306009292603,
-26.4062976837158,-10.3095359802246,
-39.0098991394043,-7.03695774078369,
-32.7491874694824,24.9877758026123,
-8.06883811950684,53.3074150085449,
10.8163070678711,41.1081237792969,
4.12896537780762,11.5192165374756,
-13.7707366943359,18.7074241638184,
-15.3015918731689,61.7007980346680,
1.94636464118958,76.9891433715820,
5.83443498611450,29.7668247222900,
-22.7606925964355,-30.2222423553467,
-56.0574188232422,-40.9570808410645,
-51.2895812988281,-13.6974658966064,
-12.5724248886108,-10.4277048110962,
17.7805061340332,-46.3384284973145,
19.8231849670410,-68.3082199096680,
12.4855871200562,-45.4625930786133,
12.2939739227295,-15.0495691299438,
16.1183338165283,-26.9857864379883,
14.8676786422730,-63.7368278503418,
14.4395275115967,-66.2001419067383,
15.6848573684692,-21.2380561828613,
5.38661241531372,20.9795284271240,
-18.3952178955078,20.6567058563232,
-27.2145423889160,-7.50962686538696,
-1.96176171302795,-25.1690673828125,
32.1639099121094,-22.0345535278320,
30.5411567687988,-9.35185337066650,
-2.76137995719910,2.31854629516602,
-16.8243637084961,16.5524978637695,
8.97476482391357,37.7620391845703,
30.7022323608398,53.5401420593262,
7.87790966033936,56.5625457763672,
-36.8488998413086,48.2685890197754,
-48.9746093750000,30.5699748992920,
-17.3289871215820,6.96464443206787,
15.1611757278442,-9.27966690063477,
13.9972829818726,-12.0846738815308,
-9.74194717407227,-10.7277345657349,
-30.6526966094971,-12.9681291580200,
-42.1053199768066,-10.9257249832153,
-43.9644889831543,2.06840944290161,
-21.6018104553223,11.6068172454834,
27.1907634735107,-1.62310624122620,
67.1516723632813,-25.5098876953125,
61.0479850769043,-16.9077281951904,
17.4885940551758,34.9672050476074,
-18.9527072906494,75.7043304443359,
-20.7809257507324,50.8969154357910,
-5.67479801177979,-18.6529731750488,
-0.0119858086109161,-55.1616020202637,
-4.79534530639648,-27.2910003662109,
-5.95691967010498,21.3181381225586,
-5.08077955245972,41.2008361816406,
-10.5985946655273,36.7610626220703,
-10.5260782241821,34.3697586059570,
8.96372222900391,30.2038898468018,
34.1380729675293,2.98272728919983,
30.3450298309326,-32.1717529296875,
-9.02023124694824,-35.2932701110840,
-43.1612129211426,1.86879813671112,
-37.0747871398926,35.1707611083984,
-6.82644796371460,29.9229774475098,
5.16127443313599,0.705109834671021,
-15.3200979232788,-18.2485580444336,
-32.3257789611816,-20.8154697418213,
-22.3903541564941,-18.2268028259277,
-3.37223339080811,-5.04514598846436,
-4.18417692184448,20.1108856201172,
-22.4952373504639,41.1597061157227,
-24.4551486968994,36.9703979492188,
0.955896735191345,10.4006919860840,
31.3777618408203,-9.71800994873047,
38.9063949584961,-15.0477628707886,
22.8442382812500,-22.3486709594727,
4.14863014221191,-39.4803390502930,
-1.68846690654755,-48.4259452819824,
1.33991527557373,-35.2816658020020,
3.28384995460510,-14.8993377685547,
-2.15206217765808,-6.82188415527344,
-22.2061290740967,-2.03239893913269,
-51.3990554809570,10.2649688720703,
-71.4131698608398,15.9589557647705,
-60.6074638366699,-4.87066745758057,
-15.6528244018555,-43.1495513916016,
39.5840530395508,-57.1260375976563,
73.4252395629883,-26.8300647735596,
70.0452041625977,17.2249927520752,
40.1507186889648,33.6514587402344,
8.85816574096680,14.2716617584229,
-9.51866054534912,-13.6418819427490,
-7.43854999542236,-24.7348575592041,
2.72204899787903,-9.22148513793945,
4.60868549346924,25.6403942108154,
-10.6324605941772,59.2242126464844,
-31.8137741088867,59.7673263549805,
-37.5285987854004,19.2110614776611,
-18.8473014831543,-27.6927871704102,
11.0871524810791,-29.2718143463135,
26.4603080749512,17.7090835571289,
14.5323276519775,60.7011260986328,
-18.7700881958008,48.6113853454590,
-46.2420272827148,-6.52702045440674,
-45.5084495544434,-45.0965576171875,
-9.15851116180420,-33.8278579711914,
43.6925926208496,0.133635282516480,
77.5944290161133,14.7940864562988,
73.1993103027344,1.59969151020050,
43.2080574035645,-15.5615348815918,
17.0776557922363,-14.0810384750366,
9.22094535827637,0.156889140605927,
5.33642053604126,4.93030261993408,
-8.06841945648193,-8.78997039794922,
-21.9792156219482,-35.9591178894043,
-16.7926826477051,-51.9216003417969,
13.6618309020996,-40.2152137756348,
47.7852096557617,-7.96109390258789,
59.2821769714356,16.0846900939941,
45.3991508483887,8.25983428955078,
24.4359436035156,-20.7938823699951,
16.7193794250488,-34.5872344970703,
23.1604518890381,-16.7294406890869,
28.9194755554199,6.79289293289185,
24.4536895751953,5.24958992004395,
17.7504329681397,-19.2577419281006,
24.9506664276123,-26.1372776031494,
40.1337089538574,6.73812198638916,
40.0795364379883,54.5735206604004,
14.1911029815674,73.7060012817383,
-15.9190025329590,50.4137115478516,
-19.9277458190918,15.2978706359863,
1.38271808624268,-2.38381814956665,
22.6618747711182,2.10033082962036,
27.5021400451660,11.0056896209717,
23.4867591857910,17.5835037231445,
21.8052234649658,27.6669464111328,
13.3231801986694,40.7033538818359,
-12.3892621994019,46.6395378112793,
-37.8737640380859,41.7001609802246,
-39.3844833374023,34.0146217346191,
-21.1733551025391,36.3393554687500,
-6.50810718536377,42.7015686035156,
-6.80763387680054,38.9642028808594,
-8.81081485748291,20.0945549011230,
-6.70392513275147,-12.4996423721313,
-15.3778057098389,-49.5531234741211,
-32.0287704467773,-74.4860458374023,
-29.8224792480469,-69.4024200439453,
6.98747348785400,-28.1933689117432,
38.6911430358887,21.4831809997559,
15.8433732986450,40.3588676452637,
-43.1842918395996,14.6364488601685,
-60.9579124450684,-25.9478549957275,
-2.26605892181397,-37.2509231567383,
72.9421386718750,-7.63319349288940,
80.8533172607422,35.2253646850586,
19.4245891571045,56.2704887390137,
-37.8672332763672,39.9997329711914,
-41.1228408813477,0.772931039333344,
-10.3100214004517,-33.2243537902832,
10.7418804168701,-43.7633628845215,
19.9654998779297,-38.3760986328125,
42.5330734252930,-29.5145645141602,
70.9484634399414,-13.9274454116821,
71.7242889404297,16.7440700531006,
33.0046195983887,44.8307037353516,
-13.0688781738281,35.8826026916504,
-32.9895362854004,-15.8986396789551,
-26.9394416809082,-62.1328697204590,
-13.9506330490112,-49.4418029785156,
-8.73562908172607,9.58650970458984,
-13.5914640426636,54.0502433776856,
-19.8398437500000,55.2744827270508,
-18.3897895812988,40.5429534912109,
-3.34778642654419,33.3228530883789,
19.6442203521729,20.7714500427246,
21.9490756988525,-12.1265630722046,
-7.28466415405273,-37.6163902282715,
-40.9694061279297,-21.2119579315186,
-43.7492294311523,23.0635757446289,
-19.0401992797852,44.4171600341797,
-2.38778400421143,32.4140434265137,
-5.55993080139160,18.6303558349609,
-4.74176788330078,19.6688728332520,
18.3699512481689,16.2521419525147,
36.6495094299316,-5.19591665267944,
14.5819282531738,-13.5932588577271,
-26.4863262176514,14.7805967330933,
-33.3827056884766,43.0187683105469,
3.21915507316589,24.2813453674316,
29.9198513031006,-25.3386459350586,
2.08762788772583,-44.3742828369141,
-54.1548118591309,-8.14729499816895,
-75.1935729980469,32.5599098205566,
-46.0160980224609,20.7409458160400,
-13.5092554092407,-36.8715438842773,
-11.9173278808594,-80.3523559570313,
-26.2823486328125,-71.2086410522461,
-18.9737071990967,-24.7205429077148,
4.01029491424561,23.3569507598877,
6.95548915863037,47.4495849609375,
-20.0844631195068,39.9225425720215,
-38.3893775939941,15.1526556015015,
-16.0687465667725,-5.15971422195435,
24.6992969512939,-11.6936712265015,
41.6517105102539,-14.7026519775391,
21.1866703033447,-19.8785381317139,
-5.66355800628662,-14.2813615798950,
-6.20368719100952,8.90212821960449,
12.2063760757446,31.3693981170654,
13.7260551452637,20.2038669586182,
-14.6790657043457,-20.5649681091309,
-47.1945686340332,-41.0110855102539,
-55.5294647216797,-16.0963211059570,
-39.6689109802246,14.7473583221436,
-26.9086093902588,0.264491319656372,
-36.6979598999023,-48.7908706665039,
-48.4779319763184,-71.0442352294922,
-26.8918590545654,-43.7388305664063,
26.4549980163574,-11.6256761550903,
68.8832550048828,-13.6841020584106,
64.2674942016602,-26.2106494903564,
25.8816432952881,-4.23315525054932,
-8.53025817871094,40.5667419433594,
-23.2216968536377,46.4881362915039,
-30.2185382843018,-0.737783193588257,
-34.3134346008301,-43.0510444641113,
-24.6161708831787,-25.0347633361816,
-3.30741620063782,31.8859367370605,
4.16825962066650,59.8675117492676,
-17.2282123565674,35.8677787780762,
-39.1230087280273,-4.52771997451782,
-31.8432941436768,-26.1291122436523,
-3.98029041290283,-27.5056934356689,
19.2444725036621,-24.4127025604248,
34.4786376953125,-15.9195852279663,
51.4011993408203,-0.471685320138931,
52.4040946960449,0.174511313438416,
18.9402656555176,-26.8288955688477,
-20.8339405059814,-56.3115043640137,
-20.6923217773438,-51.7949638366699,
19.2933387756348,-17.6116905212402,
38.0383300781250,9.05225563049316,
3.49672126770020,8.57443809509277,
-27.2180976867676,-6.40876770019531,
6.16987562179565,-16.8917922973633,
68.9204559326172,-23.3393859863281,
74.1847000122070,-26.0466747283936,
17.7820816040039,-8.59518623352051,
-21.9643859863281,34.1236686706543,
-6.66620731353760,64.5392532348633,
12.0907726287842,50.6669082641602,
-12.7003469467163,10.3557357788086,
-43.9624099731445,-6.63918590545654,
-20.5426959991455,6.42616033554077,
32.5144157409668,10.4674482345581,
42.0063209533691,-14.4663343429565,
-7.19518089294434,-34.4417915344238,
-52.9299125671387,-16.7848110198975,
-54.1491355895996,17.3926086425781,
-41.9119148254395,20.0226135253906,
-45.1224822998047,-11.5265579223633,
-33.3468055725098,-31.0921535491943,
18.2120723724365,-16.1045055389404,
64.6471481323242,4.29696226119995,
47.0160598754883,-4.34861040115356,
-17.6682014465332,-32.1939315795898,
-56.7625122070313,-48.1069831848145,
-30.7937259674072,-43.0964508056641,
21.5260734558105,-30.5346202850342,
45.3622474670410,-22.6097106933594,
33.1518859863281,-13.3322324752808,
13.3647804260254,1.84171807765961,
-4.01077842712402,16.2950134277344,
-17.4925422668457,24.3420410156250,
-20.6615676879883,27.0120658874512,
-13.6298637390137,27.7526569366455,
-11.1024141311646,18.3627109527588,
-18.1734981536865,0.407599568367004,
-16.8316268920898,-13.6271476745605,
4.82544898986816,-21.0815067291260,
21.8565845489502,-30.7885856628418,
9.44300842285156,-45.3394126892090,
-19.0390205383301,-50.9019470214844,
-25.9608325958252,-30.3526916503906,
-1.74763655662537,5.58756780624390,
10.5341176986694,27.1456775665283,
-22.5216102600098,22.0019912719727,
-69.6333618164063,5.16942501068115,
-84.7991561889648,-7.71434831619263,
-57.7654457092285,-26.8590621948242,
-14.3762569427490,-59.1338233947754,
28.2733631134033,-75.4630355834961,
62.9609718322754,-45.6174011230469,
72.6843338012695,17.8829936981201,
51.1470794677734,59.3994064331055,
24.2881736755371,46.5379295349121,
30.7261009216309,11.1047639846802,
60.9379043579102,0.732351303100586,
57.9116287231445,22.1388549804688,
-0.322640419006348,36.2654304504395,
-55.5689468383789,21.3929862976074,
-41.5753517150879,-8.33043479919434,
20.3875560760498,-29.4599609375000,
54.2732849121094,-39.9037246704102,
37.6194686889648,-36.3939247131348,
19.9056129455566,-10.2369480133057,
29.5535144805908,34.9146461486816,
31.9965019226074,66.7287902832031,
-9.88584899902344,50.9515991210938,
-60.1480178833008,-4.16874504089356,
-57.6300163269043,-57.0240211486816,
-7.35342359542847,-68.2890930175781,
28.6201019287109,-37.3992080688477,
15.3763093948364,10.4070978164673,
-8.24691486358643,49.1106338500977,
-6.56814146041870,56.9924316406250,
4.30558633804321,31.6479396820068,
-5.49559783935547,0.681676745414734,
-24.2135353088379,-2.38007211685181,
-26.2494277954102,21.9995746612549,
-11.5875997543335,39.7871055603027,
2.45585441589355,27.4601268768311,
6.42145586013794,3.98553776741028,
7.72698307037354,-2.57990646362305,
-1.21751391887665,5.36315822601318,
-25.3793907165527,2.27638959884644,
-41.3178710937500,-19.1731567382813,
-12.8124675750732,-30.0122718811035,
45.3317375183106,-20.4723205566406,
70.4167709350586,-11.8306274414063,
40.7072792053223,-19.6957588195801,
5.90837860107422,-31.1687870025635,
13.0223817825317,-20.2085514068604,
33.9510383605957,7.50373554229736,
12.8604688644409,22.4864788055420,
-42.3411712646484,19.3272609710693,
-63.0214157104492,13.4898405075073,
-16.2029094696045,13.6048021316528,
44.1862144470215,6.96299648284912,
56.0310440063477,-14.4089145660400,
30.5108623504639,-29.4350738525391,
21.5250511169434,-3.90023875236511,
40.6292953491211,52.8783111572266,
48.7950859069824,92.4284667968750,
20.6926879882813,73.2501373291016,
-19.3459815979004,10.7375011444092,
-35.1893234252930,-38.4588127136231,
-25.9007778167725,-29.2476387023926,
-8.79592800140381,20.8127193450928,
6.62016010284424,49.1396141052246,
19.4832630157471,18.0577430725098,
20.8997325897217,-35.2220611572266,
-4.10336685180664,-46.2044830322266,
-41.6885337829590,-4.48159694671631,
-56.4420623779297,30.0568256378174,
-35.3651275634766,5.25793266296387,
-10.8472423553467,-55.1965408325195,
-8.94162559509277,-86.2722702026367,
-20.4390945434570,-65.6330032348633,
-12.0500440597534,-36.9353027343750,
23.2661094665527,-34.5247650146484,
52.9184570312500,-35.4079399108887,
44.4879417419434,-17.5134563446045,
7.76177406311035,3.00775837898254,
-20.6575183868408,-6.41552209854126,
-15.7396125793457,-36.0651512145996,
20.0956230163574,-42.6121749877930,
61.7450447082520,-14.6102228164673,
79.1481857299805,12.6556186676025,
60.1861152648926,19.0911846160889,
22.2137451171875,18.8738098144531,
2.60773777961731,26.3356895446777,
16.7777462005615,20.1036834716797,
34.7995834350586,-15.2494668960571,
22.6818370819092,-48.9022598266602,
-16.4723262786865,-31.4385356903076,
-41.3848838806152,25.2060451507568,
-26.8870563507080,60.2645149230957,
4.47690296173096,39.6653976440430,
18.3296451568604,-5.25639915466309,
13.4227638244629,-22.2044410705566,
7.70784902572632,1.55727744102478,
5.06563520431519,37.7845687866211,
-6.36696195602417,58.8482170104981,
-29.6859321594238,52.7579193115234,
-45.8958892822266,22.6729335784912,
-36.1685485839844,-23.8557586669922,
-11.1832056045532,-61.9027137756348,
11.5750312805176,-69.1116485595703,
24.0628547668457,-53.0831489562988,
27.9722747802734,-38.3075294494629,
22.2744808197022,-29.7649517059326,
6.19407176971436,-11.9394254684448,
-11.4402818679810,19.3929309844971,
-12.5766458511353,45.3054504394531,
-4.01460218429565,47.3487815856934,
-5.73178958892822,27.1804256439209,
-25.7981243133545,0.220034480094910,
-40.9280776977539,-24.8898410797119,
-23.8800029754639,-40.6493110656738,
14.3627319335938,-30.9410858154297,
35.0214385986328,10.3612527847290,
16.8878040313721,49.8939056396484,
-13.6297073364258,50.2143363952637,
-14.2694311141968,13.1562032699585,
17.0578498840332,-12.5065860748291,
43.3506355285645,7.04933166503906,
30.8600883483887,46.2970657348633,
-14.5537109375000,57.9035110473633,
-56.8041954040527,31.8011856079102,
-70.9115066528320,-1.41490745544434,
-60.5120429992676,-13.8747482299805,
-41.3206214904785,-9.00940322875977,
-24.0336933135986,-4.64090442657471,
-4.23078966140747,0.365765124559402,
19.4201221466064,12.3914461135864,
36.4376068115234,28.5336418151855,
37.0040359497070,39.9185256958008,
18.7263031005859,42.7861938476563,
-4.95370197296143,46.2792854309082,
-16.3482856750488,50.2843780517578,
-12.8830299377441,43.0469360351563,
-4.10149383544922,17.3677082061768,
-0.982426702976227,-17.6985893249512,
-5.19778633117676,-45.7125053405762,
-8.84963417053223,-58.6681098937988,
1.16499841213226,-57.9795188903809,
29.8136196136475,-46.1292610168457,
63.0441017150879,-20.0719470977783,
75.0049285888672,14.7372045516968,
51.3969345092773,35.6810722351074,
3.71954488754272,23.0507602691650,
-32.8448257446289,-12.4290723800659,
-36.7806854248047,-38.2765350341797,
-13.8540000915527,-37.0366287231445,
16.5612277984619,-21.7861957550049,
38.4747657775879,-13.0862178802490,
48.8347511291504,-6.07687854766846,
41.9194679260254,15.7351512908936,
17.0449085235596,45.6627655029297,
-11.8143997192383,46.2956390380859,
-20.5248279571533,8.47395992279053,
1.62054491043091,-26.9807014465332,
37.8066215515137,-15.0943021774292,
55.2008590698242,33.7891426086426,
38.1321907043457,58.9643554687500,
-1.16799879074097,31.2754554748535,
-35.4151458740234,-14.0602989196777,
-46.6652793884277,-22.4412117004395,
-36.3096275329590,2.75896453857422,
-14.9639806747437,12.7547168731689,
13.9077749252319,-15.1418809890747,
43.1484947204590,-44.4832496643066,
56.6356315612793,-29.1299686431885,
37.8949203491211,22.7508773803711,
-7.30711460113525,62.4059638977051,
-44.1215591430664,57.9207229614258,
-47.9784011840820,29.6703186035156,
-29.8388652801514,12.1103200912476,
-19.1302223205566,8.33022975921631,
-26.0515155792236,4.85212659835815,
-31.6206092834473,0.0341543331742287,
-22.6342926025391,6.93654346466064,
-14.1268224716187,21.9194374084473,
-21.1202716827393,24.2061405181885,
-36.8307533264160,4.75955200195313,
-38.4738311767578,-6.90254163742065,
-22.2410697937012,11.1475296020508,
-3.07792520523071,35.0974311828613,
3.18759560585022,19.9512825012207,
0.829684317111969,-29.9052982330322,
5.39337062835693,-59.6909675598145,
17.5942783355713,-29.6664676666260,
34.4772148132324,27.8779411315918,
46.0131568908691,47.2207374572754,
45.5632705688477,18.0996131896973,
33.7551078796387,-16.4625988006592,
13.2260608673096,-22.1425399780273,
-8.98705005645752,-16.6979770660400,
-22.0406150817871,-30.8413543701172,
-17.6414966583252,-58.1403427124023,
-1.26523339748383,-64.3713760375977,
8.08952999114990,-40.4874000549316,
-5.43899726867676,-18.4096946716309,
-31.8663234710693,-22.2080459594727,
-34.2318763732910,-41.6057586669922,
9.03069877624512,-46.6182250976563,
67.0610961914063,-23.8817119598389,
86.8246078491211,16.4339771270752,
53.7904586791992,44.2518234252930,
10.3445510864258,35.2704315185547,
-3.33836722373962,-1.71664404869080,
3.82189536094666,-31.3684730529785,
-2.37054491043091,-27.4264144897461,
-25.0323543548584,-1.29983472824097,
-35.7002487182617,5.65142631530762,
-19.3432102203369,-17.7566299438477,
0.302318602800369,-30.0374870300293,
0.366638481616974,0.747670173645020,
-4.47799062728882,45.3209381103516,
6.43323802947998,50.8004226684570,
26.6868019104004,19.4731235504150,
34.8964271545410,6.62722015380859,
28.6403675079346,33.7015151977539,
25.1082344055176,56.5002212524414,
25.8687057495117,32.7264671325684,
13.0171318054199,-9.16027259826660,
-9.03278923034668,-11.8458843231201,
-9.49568271636963,23.5119628906250,
24.5029182434082,43.1067047119141,
56.3632659912109,17.5985603332520,
42.0369148254395,-13.5491199493408,
-3.75181770324707,-10.3134508132935,
-23.8691997528076,12.7065324783325,
7.52755928039551,18.5542793273926,
45.0547637939453,-2.39879345893860,
37.9627532958984,-25.3899021148682,
-1.81686580181122,-31.1847476959229,
-22.2936820983887,-19.2827529907227,
-5.26728534698486,1.49984860420227,
16.0410461425781,21.3280181884766,
2.98147034645081,24.5913524627686,
-33.5083618164063,7.82950115203857,
-55.2435150146484,-4.62995147705078,
-49.0321693420410,11.3194398880005,
-37.4035034179688,37.4134101867676,
-37.6405525207520,24.3311080932617,
-36.1902809143066,-33.5731163024902,
-12.2168378829956,-74.8910827636719,
27.1845169067383,-42.2338562011719,
51.0625953674316,34.2312698364258,
34.2850532531738,73.7428970336914,
-6.04286289215088,37.7966156005859,
-28.8749122619629,-26.8360214233398,
-11.2617559432983,-47.1827354431152,
26.9149723052979,-12.9273252487183,
44.7600212097168,20.3738594055176,
24.0310592651367,8.93491363525391,
-11.2003316879272,-35.6534652709961,
-22.6407432556152,-65.4311218261719,
-7.60666799545288,-55.2412452697754,
4.52295446395874,-28.5474281311035,
-1.62820458412170,-25.7731475830078,
-8.51816463470459,-52.0306320190430,
10.6941661834717,-68.4305953979492,
41.5287590026856,-33.1819801330566,
43.8745841979981,35.1596527099609,
2.50077033042908,73.4033660888672,
-42.8842887878418,44.0612297058106,
-45.3429336547852,-18.1061592102051,
-7.97595357894898,-44.2918624877930,
26.1722450256348,-7.49444389343262,
28.4952926635742,45.9598770141602,
16.9417877197266,57.3052673339844,
22.6660919189453,25.0636234283447,
39.8897132873535,-11.7522001266480,
40.2649726867676,-22.2182025909424,
14.8196554183960,-7.76947736740112,
-13.4973831176758,12.8121995925903,
-23.5356121063232,33.6838188171387,
-21.4424304962158,47.7621040344238,
-29.2107334136963,36.5271530151367,
-47.1265678405762,-8.61926078796387,
-46.4440002441406,-59.0463218688965,
-8.14188480377197,-76.7608261108398,
36.5561027526856,-54.0376014709473,
44.6547164916992,-19.6953296661377,
8.94833564758301,-2.99766492843628,
-29.2778625488281,7.61635780334473,
-27.5219631195068,31.0112781524658,
2.00260257720947,54.6240692138672,
14.8915805816650,44.0987930297852,
5.39464473724365,-1.06620764732361,
7.54006767272949,-35.9873199462891,
34.1240119934082,-20.7798557281494,
48.2566642761231,23.2371406555176,
20.2527122497559,46.2895774841309,
-16.4910621643066,28.1458339691162,
-5.46348285675049,-1.22923827171326,
44.9401626586914,-7.51173114776611,
63.0825347900391,2.40968370437622,
13.7395000457764,4.99249267578125,
-44.2723579406738,-4.77712917327881,
-41.9032440185547,-16.7277774810791,
8.45230770111084,-25.7322044372559,
32.6874313354492,-38.5868835449219,
-1.40220546722412,-49.5593338012695,
-46.0873794555664,-41.4514122009277,
-48.2050247192383,-14.8485698699951,
-23.3922595977783,0.566428840160370,
-13.7132015228271,-18.4109249114990,
-26.9719696044922,-56.4415092468262,
-28.4071712493897,-73.8495178222656,
0.589978039264679,-50.3118820190430,
37.1126174926758,-5.08793067932129,
42.8283233642578,23.4647789001465,
15.9171905517578,18.5899333953857,
-13.0225543975830,-8.12942504882813,
-14.8271932601929,-33.7042274475098,
6.97562026977539,-43.5875625610352,
29.3493003845215,-38.1979179382324,
30.4818229675293,-25.7841434478760,
12.0695276260376,-14.8961286544800,
2.42357492446899,-2.88803505897522,
23.4489917755127,9.74756717681885,
55.3451690673828,19.7654285430908,
63.4796371459961,20.4341468811035,
36.7954216003418,15.9591197967529,
4.75405120849609,13.7048654556274,
2.38247418403626,12.0124721527100,
29.4697456359863,8.36659145355225,
51.9509658813477,0.351760238409042,
47.3484573364258,-0.829098820686340,
28.3354682922363,6.72407817840576,
14.3907527923584,8.84386348724365,
13.9061698913574,-6.18272113800049,
24.1577606201172,-22.7917079925537,
38.3751068115234,-16.4659404754639,
42.3148002624512,17.0679416656494,
18.1459140777588,46.7335968017578,
-32.1502265930176,48.2166633605957,
-74.9392089843750,29.0644969940186,
-75.1688079833984,13.6325445175171,
-39.5525817871094,6.21069955825806,
-12.2537574768066,-7.97967195510864,
-14.4060020446777,-32.5175628662109,
-22.4312038421631,-49.6421508789063,
-6.86062145233154,-40.3635673522949,
22.5365619659424,-17.9693069458008,
29.2482299804688,-12.0236444473267,
10.1797199249268,-33.3868064880371,
-5.84494638442993,-57.9641036987305,
3.77420020103455,-53.4899330139160,
22.1231307983398,-13.8503551483154,
24.3226337432861,33.8344497680664,
17.6047191619873,52.0624237060547,
26.2773342132568,29.2893161773682,
42.8740692138672,-3.86735773086548,
38.3620147705078,-8.77981948852539,
1.87920427322388,12.6256589889526,
-33.8003845214844,22.6054096221924,
-33.0803260803223,-5.23061466217041,
-5.48352241516113,-47.1101303100586,
19.2541961669922,-62.1923522949219,
28.8964920043945,-42.9202957153320,
34.4048194885254,-22.8959751129150,
39.5667495727539,-19.7502212524414,
28.9156303405762,-15.9651460647583,
-3.13780069351196,2.23805856704712,
-30.4161872863770,15.1890506744385,
-23.9417953491211,9.40292167663574,
4.79360914230347,3.88637685775757,
21.0391159057617,24.7966365814209,
7.25063610076904,55.4317207336426,
-24.6181011199951,56.3809127807617,
-46.9649772644043,25.0973358154297,
-47.9395599365234,0.872574567794800,
-25.3937339782715,3.62154221534729,
6.54596328735352,4.82457923889160,
26.8888549804688,-16.9201240539551,
19.9476337432861,-35.9374198913574,
-3.91458249092102,-18.3482189178467,
-15.5977096557617,15.1097412109375,
-6.59865379333496,18.3051776885986,
-2.95486187934876,-10.6768808364868,
-29.3015937805176,-24.3653373718262,
-63.6724319458008,-6.41561412811279,
-60.8378562927246,7.58121681213379,
-12.9495925903320,-14.9441061019897,
36.3109245300293,-45.7560882568359,
40.9692916870117,-35.4219360351563,
1.21803712844849,9.82605743408203,
-41.7206497192383,36.4495506286621,
-55.3501243591309,12.8144445419312,
-42.5793151855469,-26.4960002899170,
-26.8859634399414,-38.0050163269043,
-24.6637172698975,-17.0838279724121,
-30.1944770812988,7.17224788665772,
-30.3854293823242,13.6646623611450,
-17.2774696350098,2.26284098625183,
-0.329824745655060,-22.6268539428711,
1.70975613594055,-52.0657157897949,
-6.99018001556397,-70.9516448974609,
-5.44546079635620,-63.0140876770020,
14.5148124694824,-29.9486122131348,
33.1053962707520,4.55443429946899,
30.4422626495361,21.8933200836182,
12.2522735595703,27.8782749176025,
0.134513825178146,33.0389404296875,
-1.73251044750214,28.7242240905762,
-14.4840402603149,4.77348804473877,
-36.7417221069336,-28.6867446899414,
-36.0766334533691,-43.9885139465332,
4.59035968780518,-24.3987159729004,
48.8243637084961,15.9336080551147,
39.1630363464356,46.9664039611816,
-20.2965316772461,52.6633529663086,
-65.3946304321289,34.5261917114258,
-48.0308303833008,8.60397529602051,
10.0821065902710,-9.34552478790283,
48.2938880920410,-7.57208299636841,
38.4011383056641,14.0029859542847,
8.75071144104004,29.5353317260742,
1.06822764873505,19.4748191833496,
26.9152221679688,-6.94079208374023,
57.5983619689941,-23.5655288696289,
57.6847648620606,-14.3807373046875,
15.1660404205322,6.20360612869263,
-42.9100952148438,13.9879360198975,
-61.7349319458008,1.82608437538147,
-20.7199192047119,-16.2968482971191,
39.2648468017578,-19.8026504516602,
52.5020370483398,1.42823016643524,
10.0262250900269,43.7530250549316,
-31.0139102935791,77.4067459106445,
-24.9067192077637,66.6329650878906,
9.48554801940918,10.1668024063110,
23.1228179931641,-40.2562789916992,
10.2949724197388,-32.6445770263672,
7.53374147415161,20.0880546569824,
23.9176521301270,52.4819793701172,
23.3419647216797,29.0210094451904,
-11.8424463272095,-17.4057559967041,
-38.5336723327637,-33.8172492980957,
-14.8582963943481,-13.9147968292236,
41.8577690124512,4.70402383804321,
70.0077972412109,3.81259465217590,
48.3446273803711,3.23259282112122,
14.3934917449951,14.5716810226440,
5.24254131317139,23.1640300750732,
17.4427871704102,18.6977100372314,
27.2824783325195,11.3271074295044,
25.4778137207031,11.1166534423828,
17.5175991058350,8.03943920135498,
-3.51985597610474,-3.00055789947510,
-31.6736316680908,-6.49347066879273,
-36.5203971862793,5.21556377410889,
-3.16460371017456,12.7011890411377,
41.0193290710449,-5.35816287994385,
55.2727050781250,-30.7057571411133,
42.7955017089844,-18.1831150054932,
39.7363891601563,29.2915153503418,
49.0496635437012,53.9705734252930,
38.6770248413086,29.3922767639160,
-2.89748764038086,-7.91128349304199,
-30.8931674957275,-12.0838012695313,
-9.30226707458496,9.30965805053711,
24.3766040802002,20.5761184692383,
6.09899520874023,14.6302642822266,
-55.1019477844238,13.2557067871094,
-81.6890716552734,15.6619615554810,
-36.2299690246582,-1.75169897079468,
33.3647422790527,-29.1999340057373,
59.3335914611816,-23.0325202941895,
29.0344657897949,23.9019718170166,
-18.1617813110352,51.5667800903320,
-47.7095642089844,11.5577983856201,
-45.5205726623535,-55.5277595520020,
-14.7097377777100,-71.6162414550781,
34.2933158874512,-27.1249160766602,
69.9436340332031,14.7384414672852,
72.6562805175781,13.2663431167603,
57.9638061523438,-0.723257362842560,
56.2707939147949,17.0985813140869,
56.9529342651367,50.0184745788574,
22.9846172332764,48.8973388671875,
-35.0500183105469,9.43585491180420,
-58.9073410034180,-24.7162933349609,
-18.7491416931152,-25.4985313415527,
43.9149856567383,-12.4867124557495,
70.0347290039063,-6.74402952194214,
54.9857139587402,0.624816775321960,
41.4037780761719,20.4736766815186,
44.0564727783203,31.5147724151611,
38.5882568359375,13.8897590637207,
18.8641757965088,-19.9709739685059,
7.38607597351074,-30.4389152526855,
13.0473136901855,-1.82993519306183,
12.4987182617188,29.6711158752441,
-9.12486743927002,27.9405384063721,
-16.6529293060303,0.795955181121826,
14.5336208343506,-13.1745634078980,
55.2052154541016,4.52079677581787,
47.7784729003906,35.3012046813965,
-5.80339384078980,51.4247322082520,
-45.1760101318359,39.6717987060547,
-29.0812034606934,18.9211864471436,
11.5919237136841,17.8373451232910,
17.2958831787109,39.7920188903809,
-15.5804300308228,62.5854339599609,
-36.5521049499512,60.6740684509277,
-12.2173690795898,31.7798347473145,
32.2508430480957,-0.656630516052246,
53.2633895874023,-14.7949504852295,
30.4494514465332,-15.6075162887573,
-14.6868171691895,-15.7961997985840,
-45.0776062011719,-7.24397039413452,
-42.2559242248535,20.9184398651123,
-23.8697280883789,44.0910186767578,
-16.6450080871582,26.2537307739258,
-25.3578910827637,-29.5604133605957,
-26.7778968811035,-60.4391403198242,
-5.05916166305542,-18.9455585479736,
17.4500694274902,55.8259124755859,
-0.166483402252197,77.9891357421875,
-50.1617240905762,23.4881362915039,
-66.3793106079102,-38.4072036743164,
-16.5487232208252,-38.4356231689453,
45.2389183044434,7.99187517166138,
52.1359939575195,30.8815250396729,
11.2663345336914,10.5094718933105,
-8.15169620513916,-7.53723096847534,
21.3654708862305,8.52185916900635,
43.9226112365723,33.3200645446777,
14.7633800506592,22.8915748596191,
-26.3441982269287,-23.2006492614746,
-19.2673988342285,-60.1636581420898,
20.0330810546875,-56.9659881591797,
23.8671722412109,-18.9919395446777,
-12.3980331420898,24.9864807128906,
-24.4932556152344,46.8196868896484,
15.5754070281982,37.4142684936523,
45.4533958435059,6.55960988998413,
7.69477033615112,-11.0562295913696,
-57.6181716918945,-3.70903944969177,
-71.5778350830078,2.61825919151306,
-24.9110450744629,-17.9165954589844,
15.1194496154785,-44.5567512512207,
9.06257915496826,-36.5640983581543,
-5.65118551254273,5.17544460296631,
7.95828294754028,30.2486324310303,
25.7705554962158,4.07717561721802,
13.6398944854736,-39.4155960083008,
-9.91594409942627,-45.2623939514160,
-5.41579961776733,-14.4573879241943,
19.0167312622070,10.3467054367065,
27.7991466522217,15.7431783676147,
12.5665931701660,25.4453792572022,
2.63706016540527,50.2717704772949,
8.43532752990723,63.5139045715332,
5.44673681259155,50.3359718322754,
-20.0461940765381,32.7178688049316,
-40.6852607727051,32.2599220275879,
-25.7160625457764,31.4778976440430,
0.946877777576447,2.27330112457275,
1.14747667312622,-41.1155624389648,
-24.4856910705566,-56.3254470825195,
-42.1193389892578,-27.2418537139893,
-37.0008392333984,9.87502098083496,
-20.3549346923828,19.9811611175537,
0.658993124961853,7.83352184295654,
27.2850570678711,-5.39017724990845,
55.8162574768066,-15.0343589782715,
64.6120834350586,-16.3925628662109,
44.4668540954590,-2.57653665542603,
14.1350564956665,24.6609439849854,
-6.86873960494995,41.0375862121582,
-25.1016979217529,27.8894901275635,
-45.4638748168945,2.38193607330322,
-50.1235160827637,-6.90717220306397,
-29.0033874511719,-0.0623154044151306,
-10.6209630966187,-7.24096822738648,
-23.9824447631836,-33.2986488342285,
-46.6567230224609,-45.5519332885742,
-28.6899833679199,-25.9835834503174,
27.8757400512695,-5.26323127746582,
61.8580970764160,-12.7165069580078,
29.1577682495117,-30.7806320190430,
-28.4569950103760,-17.8262462615967,
-41.2511558532715,26.3245906829834,
-6.45960950851440,56.1811294555664,
17.9981422424316,47.2044868469238,
0.00294852256774902,21.9811210632324,
-24.9943046569824,9.05779743194580,
-18.7643947601318,-1.28069686889648,
9.54231357574463,-33.3999328613281,
23.4953517913818,-70.8817062377930,
16.8920783996582,-71.9107589721680,
6.09844827651978,-28.4766960144043,
-1.67473459243774,18.6235694885254,
-16.6712532043457,24.9007186889648,
-34.2219200134277,-5.18812227249146,
-33.2109718322754,-37.2028160095215,
-10.5057601928711,-41.1531639099121,
7.89613103866577,-21.4720897674561,
1.90189909934998,-4.12172365188599,
-10.3297529220581,-11.7402982711792,
-1.98175764083862,-39.9130668640137,
18.7173290252686,-59.8423309326172,
22.0525302886963,-44.1405639648438,
-0.498831510543823,4.53349733352661,
-23.3287429809570,47.0572662353516,
-24.4298343658447,49.1067886352539,
-11.5495424270630,16.3539352416992,
-9.26368808746338,-17.9455986022949,
-16.9022960662842,-37.3362846374512,
-8.92230415344238,-42.8419723510742,
20.9447727203369,-40.3528442382813,
43.2511901855469,-31.1030902862549,
30.0636463165283,-17.2714633941650,
-9.54290676116943,-8.41232681274414,
-35.8749618530273,-7.18404912948608,
-22.0468406677246,-4.70875263214111,
12.5983133316040,1.30460751056671,
27.6102447509766,1.82688903808594,
8.47525691986084,-7.27936649322510,
-12.2772283554077,-8.63436794281006,
-1.02843606472015,9.26197052001953,
35.6070365905762,29.4642028808594,
53.5477447509766,19.8784980773926,
21.2285385131836,-11.7406177520752,
-35.6112518310547,-27.6434421539307,
-53.8830146789551,-10.4118518829346,
-10.9284648895264,16.3497962951660,
47.0262451171875,22.7724018096924,
60.8803176879883,16.3746452331543,
26.0346221923828,20.2326354980469,
-12.4365015029907,30.4440269470215,
-18.6002578735352,17.3873195648193,
-2.40654540061951,-15.8439340591431,
15.6386308670044,-33.1375122070313,
37.3394927978516,-18.2064552307129,
66.2135009765625,0.596166610717773,
76.6657867431641,0.625753998756409,
45.2593879699707,1.49885690212250,
-5.46950435638428,31.1376018524170,
-21.0993309020996,66.1925888061523,
10.4242820739746,58.6389579772949,
41.7894058227539,11.6810493469238,
31.4957828521729,-15.1593828201294,
-2.10680842399597,7.31402587890625,
-19.6070575714111,32.0555801391602,
-10.4922637939453,7.65297508239746,
7.35418272018433,-43.4811820983887,
18.8625259399414,-57.7046890258789,
29.3062057495117,-24.1456813812256,
37.0473365783691,3.22581911087036,
29.7399063110352,-4.29753589630127,
10.7962398529053,-14.4619855880737,
-2.46354746818543,7.09297752380371,
-11.3713626861572,40.5399818420410,
-28.0085163116455,41.6692619323731,
-44.1597328186035,14.3741273880005,
-28.3123893737793,5.10855150222778,
11.9161615371704,25.7103557586670,
28.9510746002197,38.9375114440918,
2.40544843673706,14.8316402435303,
-27.5507984161377,-26.3265495300293,
-12.4770202636719,-47.5930023193359,
27.1253929138184,-36.4861373901367,
32.1409721374512,-7.70710659027100,
-1.76595449447632,22.3316917419434,
-18.9914226531982,40.2735443115234,
3.27826738357544,34.0596618652344,
20.3701858520508,4.12869596481323,
-7.96614837646484,-21.2975769042969,
-50.3412322998047,-15.8211889266968,
-52.8205223083496,5.19184064865112,
-23.4273853302002,-1.13199472427368,
-10.5191698074341,-38.1866836547852,
-23.9598999023438,-56.5022964477539,
-22.5502586364746,-21.0541915893555,
16.1635551452637,34.6157150268555,
55.6691017150879,46.8660812377930,
51.4610977172852,5.25658178329468,
14.3198165893555,-38.3086891174316,
-10.3515300750732,-34.7022476196289,
-2.66142034530640,1.77009856700897,
15.9084682464600,26.8290157318115,
19.3793792724609,21.0242385864258,
-1.50944459438324,2.53533983230591,
-37.6058235168457,-9.24358749389648,
-65.5712890625000,-20.8353652954102,
-58.1097831726074,-38.2471580505371,
-9.96150493621826,-50.4146652221680,
39.8470268249512,-40.6646308898926,
41.3783111572266,-11.5903644561768,
-9.48753738403320,15.4364557266235,
-56.9274177551270,20.6292762756348,
-45.2382812500000,5.85182285308838,
12.3268241882324,-7.32016992568970,
51.8944168090820,-8.93842411041260,
36.4207992553711,-8.42973613739014,
-0.797284841537476,-15.8265790939331,
-10.2240295410156,-29.0479412078857,
12.6572971343994,-26.7858657836914,
28.0542831420898,-2.96520161628723,
9.00228500366211,23.7575988769531,
-20.3325862884522,31.4640483856201,
-26.2610511779785,25.3305492401123,
-9.08922767639160,29.4398708343506,
0.101745963096619,47.0351409912109,
-19.5768795013428,51.1908531188965,
-45.5102348327637,27.4113025665283,
-50.6786613464356,-4.78013944625855,
-38.8134727478027,-11.7298192977905,
-29.8471050262451,8.33865737915039,
-33.7107391357422,22.5160026550293,
-38.1832275390625,11.1261606216431,
-26.9855995178223,-14.9130115509033,
-7.46160030364990,-34.0632896423340,
5.05456781387329,-44.0764923095703,
14.6053819656372,-49.3762702941895,
32.4179039001465,-42.3265686035156,
56.7582015991211,-13.3263235092163,
63.3336105346680,19.9449348449707,
30.4648838043213,26.0966949462891,
-27.0757827758789,3.04317188262939,
-61.3792800903320,-17.7646636962891,
-48.0550003051758,-6.50506782531738,
-14.2565670013428,23.6776866912842,
-9.49637413024902,37.6456451416016,
-39.1541557312012,20.2750530242920,
-57.7073860168457,-11.6604995727539,
-26.8413619995117,-32.8758621215820,
25.7416152954102,-38.3363113403320,
37.3211936950684,-30.8938827514648,
-10.0768623352051,-13.2282485961914,
-61.4094352722168,1.21033656597137,
-62.3151397705078,-0.480628907680512,
-22.1723194122314,-15.5433940887451,
6.25914525985718,-21.3107471466064,
-3.50437045097351,-3.26483798027039,
-28.5935115814209,23.8240432739258,
-38.6064262390137,28.0092754364014,
-32.6589431762695,1.80513429641724,
-21.3139343261719,-27.6005649566650,
-5.86562919616699,-34.2718582153320,
8.94607543945313,-13.9646854400635,
11.4395866394043,21.0061874389648,
-7.58089971542358,58.1546058654785,
-30.2643394470215,72.2300796508789,
-30.9341411590576,42.5449066162109,
-4.76384067535400,-18.8953971862793,
20.7991809844971,-61.2501640319824,
22.8813381195068,-41.4240570068359,
2.68862318992615,15.0027427673340,
-29.1331539154053,40.0523223876953,
-55.3677330017090,4.75215053558350,
-54.2458076477051,-41.6772575378418,
-19.1285934448242,-39.3491020202637,
22.1635265350342,7.94803810119629,
28.9092006683350,47.7892837524414,
-8.47984409332275,50.2813110351563,
-54.8142395019531,30.0580425262451,
-71.3221664428711,7.81227636337280,
-54.0724334716797,-16.6940841674805,
-26.0365715026855,-45.6710510253906,
1.56889152526855,-55.7104835510254,
27.7029476165772,-29.1455459594727,
38.7266120910645,6.39949417114258,
23.0022392272949,16.9423694610596,
6.16163110733032,4.33548259735107,
16.0695896148682,6.81775236129761,
38.3542137145996,36.0086708068848,
30.3313465118408,49.0964736938477,
-10.4314594268799,20.9510879516602,
-27.0077724456787,-20.8039646148682,
10.9769630432129,-27.0171279907227,
55.3667259216309,4.26042842864990,
38.4929275512695,22.0159587860107,
-26.0369567871094,-4.04952478408814,
-59.7859420776367,-44.5128021240234,
-32.4255371093750,-58.9029731750488,
-0.0614707469940186,-44.7713813781738,
-5.94468784332275,-33.0896186828613,
-21.3236045837402,-40.2592849731445,
5.03412485122681,-51.0435028076172,
57.2812347412109,-49.4858245849609,
71.2249450683594,-29.4928283691406,
34.4794616699219,7.33715105056763,
-2.47194218635559,50.4261016845703,
-3.10489201545715,79.6685485839844,
8.30730533599854,73.4260330200195,
-7.66994524002075,27.4737892150879,
-37.9347267150879,-27.9923534393311,
-37.6831283569336,-52.2733840942383,
-2.70539021492004,-31.9268951416016,
21.4231491088867,9.12819671630859,
12.9044342041016,31.2691268920898,
-1.95645773410797,14.5429096221924,
9.85341739654541,-22.5550231933594,
40.6310424804688,-38.0015792846680,
46.9860610961914,-15.4365615844727,
12.9800958633423,17.7017555236816,
-33.1466865539551,19.5439567565918,
-47.4548225402832,-10.3261451721191,
-22.3626861572266,-35.9687156677246,
11.5473089218140,-25.3290119171143,
25.1634788513184,5.33991813659668,
13.5640392303467,21.5452117919922,
-5.24917984008789,13.1626939773560,
-7.30314207077026,-0.430068403482437,
14.8746643066406,-7.11721181869507,
43.8962440490723,-10.6788711547852,
54.5580215454102,-10.4017534255981,
30.0164642333984,-0.297268390655518,
-17.9235706329346,18.6242866516113,
-49.7885780334473,23.6659564971924,
-34.7339820861816,-0.989586472511292,
20.6090202331543,-35.1710243225098,
68.0569686889648,-40.2378578186035,
72.0174179077148,-6.61499738693237,
35.7443847656250,36.0085334777832,
-0.679302275180817,51.1951560974121,
-1.37052154541016,32.4060554504395,
22.9067649841309,7.02166652679443,
37.8222961425781,6.11874532699585,
23.8895835876465,25.2864208221436,
-5.88268947601318,39.3928642272949,
-25.3117790222168,22.8929901123047,
-24.0657711029053,-21.3448772430420,
-10.3388824462891,-58.6342544555664,
8.72166633605957,-56.3932838439941,
36.9273109436035,-20.8779640197754,
71.2302093505859,7.90843105316162,
82.4414825439453,7.91694259643555,
43.9519500732422,-0.687701940536499,
-20.2297744750977,4.20079421997070,
-48.4143600463867,12.9717712402344,
-10.5380115509033,1.68731224536896,
52.1971092224121,-21.2190208435059,
66.9028015136719,-12.0896797180176,
24.3150081634522,41.1557540893555,
-16.7923374176025,81.2278823852539,
-10.8798503875732,60.6317596435547,
12.6691474914551,6.07882499694824,
2.26532053947449,-16.8959312438965,
-36.9531860351563,0.375625759363174,
-53.1371002197266,4.18800497055054,
-24.9453449249268,-24.2929191589355,
14.5233268737793,-33.7149467468262,
25.7853031158447,10.7568235397339,
9.90729618072510,63.8888359069824,
-7.55056810379028,56.7205505371094,
-23.6006278991699,-3.55816960334778,
-41.4722938537598,-42.3660774230957,
-45.6673622131348,-27.2104473114014,
-25.4035282135010,-2.26282358169556,
-0.393171429634094,-12.3418674468994,
-6.52379655838013,-39.9815673828125,
-34.1015167236328,-47.8214416503906,
-32.9767837524414,-33.4442596435547,
13.5973072052002,-15.8086662292480,
52.0009651184082,4.42534923553467,
31.7808742523193,27.5276546478272,
-24.3194942474365,38.2722434997559,
-46.1918334960938,20.2989406585693,
-12.0448293685913,-6.45583677291870,
20.2553310394287,-5.68291378021240,
-1.05634903907776,21.5249843597412,
-51.3115081787109,34.2985115051270,
-69.4464187622070,11.1028680801392,
-38.3726310729981,-18.4675006866455,
4.93457508087158,-26.5942077636719,
26.3177356719971,-23.3972148895264,
35.8121299743652,-26.3443279266357,
50.2509613037109,-28.2767238616943,
61.6463928222656,-13.6219511032105,
56.2298736572266,6.71858167648315,
38.9817352294922,6.05764961242676,
28.9886493682861,-18.5108261108398,
30.7025089263916,-34.0076560974121,
23.3819179534912,-22.3311443328857,
-0.141354322433472,1.70384192466736,
-18.4983615875244,12.4190549850464,
-13.4016389846802,8.21275997161865,
3.26367282867432,5.38835191726685,
4.27310609817505,3.69899582862854,
-19.4983367919922,-2.64658164978027,
-46.5572586059570,-4.85411691665649,
-48.1913414001465,6.78455829620361,
-29.2690429687500,23.9609794616699,
-21.7712917327881,24.1028709411621,
-41.1141242980957,-1.48073887825012,
-65.7660522460938,-25.5700244903564,
-57.6887741088867,-19.4031791687012,
-16.7774047851563,16.0156478881836,
18.7208003997803,48.4251022338867,
16.2382793426514,54.5684814453125,
-5.83970212936401,30.7677097320557,
-5.64042949676514,-12.7776775360107,
20.7350864410400,-58.5038146972656,
34.0417022705078,-77.8288650512695,
14.5387945175171,-49.0119628906250,
-7.65710258483887,8.84347343444824,
2.21890759468079,42.9718475341797,
32.3274154663086,18.9173374176025,
37.3320388793945,-37.1715736389160,
3.83618354797363,-64.6624984741211,
-30.6830444335938,-41.4739837646484,
-33.7335281372070,1.03882479667664,
-15.9235992431641,24.1284942626953,
-5.56425094604492,26.3927669525147,
-4.66371822357178,32.6331481933594,
2.19148063659668,46.7157211303711,
14.8265123367310,54.8972663879395,
12.3515615463257,43.1309585571289,
-10.1919727325439,19.0025749206543,
-26.3206901550293,-6.89541244506836,
-12.0814361572266,-28.0181388854980,
22.3703384399414,-35.4291534423828,
45.8112106323242,-21.1989059448242,
43.2695617675781,14.9872646331787,
24.9891872406006,54.2024307250977,
8.33561038970947,69.4028701782227,
-2.46120309829712,57.9598884582520,
-13.0455541610718,36.9971694946289,
-22.0075416564941,25.9336681365967,
-23.6025180816650,33.2383766174316,
-20.5110340118408,48.4080657958984,
-19.7019290924072,60.6128997802734,
-22.8116245269775,63.1990585327148,
-23.8001308441162,58.4858398437500,
-16.3384361267090,48.6460266113281,
-6.29111766815186,34.2166938781738,
-6.24329614639282,17.4897537231445,
-22.4363327026367,3.56230640411377,
-38.2992935180664,2.15157318115234,
-38.0048751831055,16.3395004272461,
-22.0444335937500,40.2805442810059,
-6.56942605972290,55.8995170593262,
-4.17421245574951,50.8429756164551,
-3.34863567352295,30.1074810028076,
11.9447603225708,7.97005224227905,
35.3932533264160,1.91220307350159,
42.1201972961426,15.9561872482300,
15.4389209747314,41.1490974426270,
-23.1767520904541,62.2327117919922,
-37.0079879760742,68.1897430419922,
-21.6670341491699,54.8915596008301,
-5.48173952102661,31.2449474334717,
-13.0652799606323,10.4049911499023,
-40.3405494689941,0.209508731961250,
-57.6275558471680,-7.24228906631470,
-49.9929008483887,-19.2180995941162,
-25.0853691101074,-28.4429798126221,
2.12871098518372,-23.0288944244385,
14.5728149414063,-6.80001640319824,
3.02961015701294,-2.22554945945740,
-29.4054336547852,-17.0736160278320,
-51.7608680725098,-33.1325035095215,
-33.2217407226563,-24.4571380615234,
8.83015823364258,1.02288556098938,
17.8426971435547,13.2220354080200,
-29.1106147766113,7.88701486587524,
-80.7573699951172,8.46350002288818,
-69.5852203369141,22.1671943664551,
2.68199634552002,26.2346839904785,
64.7536010742188,2.97162199020386,
69.1164169311523,-21.8001155853272,
38.4742279052734,-15.4352560043335,
12.9153337478638,9.92542743682861,
-10.5510349273682,15.2781305313110,
-40.5718650817871,-1.85608434677124,
-55.1289367675781,-7.17241621017456,
-27.7391910552979,14.2571353912354,
15.1990976333618,26.4677734375000,
17.1545524597168,-3.49054551124573,
-22.0214767456055,-47.2556152343750,
-34.7434425354004,-52.2172355651856,
11.7673454284668,-16.5472145080566,
58.9642715454102,15.5383100509644,
32.3524246215820,16.5404281616211,
-46.1660423278809,1.99519360065460,
-86.7289581298828,3.18144679069519,
-48.9502792358398,22.7279605865479,
2.49921393394470,39.4739227294922,
-2.18572664260864,31.5409698486328,
-44.9115066528320,1.03434038162231,
-56.8579864501953,-31.4018764495850,
-20.3478221893311,-35.6023674011231,
16.9499244689941,0.117747068405151,
17.4761352539063,41.9237556457520,
-0.416958600282669,45.7947235107422,
-3.08119177818298,8.72323703765869,
3.64539337158203,-23.7440757751465,
-5.95005989074707,-20.5266151428223,
-24.6369800567627,-7.60585832595825,
-15.6124753952026,-19.1625785827637,
24.6719264984131,-46.2956695556641,
53.3715629577637,-49.9867515563965,
37.4761962890625,-23.4467144012451,
0.544152021408081,-5.91851282119751,
-12.3601608276367,-24.2356224060059,
13.8492126464844,-53.1101112365723,
39.8302650451660,-49.2726936340332,
38.8674316406250,-5.36964273452759,
26.1543865203857,44.6625747680664,
23.0342025756836,66.7601623535156,
26.2717895507813,51.5474319458008,
14.2826004028320,12.1715354919434,
-10.3354778289795,-25.8524246215820,
-24.2069664001465,-37.4558372497559,
-23.6073036193848,-19.6981983184814,
-29.1165332794189,5.08944511413574,
-51.2905044555664,12.7391633987427,
-68.1832580566406,2.54594230651855,
-46.0017509460449,-6.46049070358276,
11.5024738311768,-3.23259353637695,
63.4214248657227,5.07264709472656,
81.8072280883789,7.16684007644653,
69.1006774902344,12.9293212890625,
42.1035346984863,34.6050949096680,
7.77390956878662,57.6423187255859,
-35.4757423400879,54.1046752929688,
-71.8961029052734,19.7942790985107,
-68.2798538208008,-17.6344470977783,
-13.3724317550659,-27.6835403442383,
47.0053329467773,-10.4500341415405,
49.3223037719727,10.8256483078003,
-7.69601249694824,20.2664279937744,
-55.3820228576660,17.7312622070313,
-35.0630455017090,4.91190385818481,
23.5095634460449,-16.7078514099121,
41.4782562255859,-31.5408020019531,
-4.68919372558594,-16.3979835510254,
-46.7360458374023,14.9355497360230,
-26.2541465759277,23.2677135467529,
22.6753387451172,-11.4440050125122,
31.5043869018555,-50.8128814697266,
-3.29769659042358,-52.0145874023438,
-20.2161884307861,-28.2374095916748,
3.93974733352661,-23.3026847839355,
21.6890621185303,-43.6483917236328,
-7.49470996856689,-43.7499313354492,
-45.9737586975098,-2.62136125564575,
-37.3551940917969,34.5761413574219,
4.17989253997803,28.3245925903320,
24.1970291137695,10.0274267196655,
5.75346517562866,30.1745223999023,
-10.2331724166870,74.4948883056641,
5.36446666717529,76.9229202270508,
20.9182319641113,13.6112937927246,
4.87811660766602,-61.9705963134766,
-18.9791221618652,-89.1689224243164,
-10.5421590805054,-66.7359008789063,
22.7103595733643,-29.4907150268555,
41.7159538269043,4.88658380508423,
28.9796752929688,31.9954128265381,
5.11817693710327,36.4985885620117,
-2.81966495513916,6.89635658264160,
11.1614761352539,-25.3899116516113,
38.2059860229492,-17.1718158721924,
62.6519622802734,19.6442108154297,
62.1867332458496,30.8715953826904,
19.8888053894043,-0.665858268737793,
-36.9467506408691,-30.1701126098633,
-50.4146118164063,-14.1554117202759,
-5.45201444625855,28.7544841766357,
47.2838211059570,46.5822792053223,
53.5111999511719,23.5279483795166,
24.7443084716797,-2.38439440727234,
6.09861183166504,-0.858425736427307,
14.8001775741577,13.2439308166504,
19.7897968292236,20.2192115783691,
1.80486440658569,15.8566589355469,
-15.2317380905151,7.06893873214722,
-9.46166324615479,-2.99212956428528,
-1.48706340789795,-4.82692003250122,
-12.6843738555908,5.93959045410156,
-26.2243518829346,15.4086217880249,
-12.3949270248413,4.12265825271606,
20.1516380310059,-27.5658550262451,
31.2821483612061,-49.3227691650391,
22.2530117034912,-38.3765869140625,
34.1958236694336,-11.9080142974854,
76.6773376464844,3.54647564888001,
99.5986404418945,11.7300415039063,
57.9275741577148,36.4014091491699,
-18.6944847106934,58.9604492187500,
-49.7781028747559,40.3732070922852,
-13.7126388549805,-10.2598524093628,
31.5652980804443,-30.5165634155273,
25.7750053405762,10.0245418548584,
-19.3888206481934,58.3604698181152,
-53.2718963623047,45.0269966125488,
-48.0312042236328,-19.0142974853516,
-15.1325330734253,-61.4299392700195,
20.4065780639648,-44.6609878540039,
36.9011383056641,-3.10240983963013,
29.1073932647705,25.0596065521240,
9.18132972717285,48.9232521057129,
-2.92578244209290,78.7822265625000,
4.11946010589600,79.8190231323242,
12.3793334960938,29.0427207946777,
2.30802154541016,-34.4967079162598,
-21.3088645935059,-49.2101631164551,
-30.1243877410889,-12.0711002349854,
-27.1400260925293,19.3530197143555,
-32.5192222595215,13.9106397628784,
-42.6906433105469,-3.30566287040710,
-31.3713397979736,-3.45318460464478,
-1.55380678176880,-4.33423233032227,
6.94497632980347,-25.4736938476563,
-23.8522777557373,-35.5992851257324,
-49.8167304992676,-0.866464138031006,
-23.9556179046631,45.3133583068848,
27.6701507568359,40.2252426147461,
41.7667541503906,-18.3936614990234,
8.64485645294190,-59.7522315979004,
-7.72878265380859,-32.8714447021484,
27.2241134643555,24.2021903991699,
66.4198837280273,52.7155151367188,
48.6527519226074,42.3326034545898,
-12.7448387145996,29.1690616607666,
-54.9963035583496,20.8790016174316,
-52.7425880432129,-7.61028480529785,
-27.7924404144287,-47.9596138000488,
-5.37114048004150,-52.0614166259766,
12.8701944351196,-4.26322650909424,
26.0155086517334,43.8625450134277,
24.7083415985107,39.9668617248535,
11.1946029663086,-0.507806777954102,
10.7485055923462,-24.9916915893555,
33.3884620666504,-13.8010673522949,
53.4253273010254,6.70693349838257,
48.5064315795898,17.4405574798584,
34.5167465209961,33.0328788757324,
24.2342300415039,62.0552215576172,
4.70549631118774,78.1252670288086,
-27.8487930297852,58.3511085510254,
-41.3830337524414,24.2308502197266,
-12.8484935760498,8.94495010375977,
25.4871788024902,13.6084871292114,
17.3598690032959,16.6663074493408,
-31.6086483001709,9.43501567840576,
-47.6878547668457,5.25679016113281,
2.61002898216248,3.91138029098511,
58.1475524902344,-3.29257655143738,
50.5802459716797,-20.8296871185303,
6.38393974304199,-32.1025657653809,
0.657845735549927,-23.7370929718018,
39.1469993591309,-3.81400299072266,
55.4475212097168,17.2434043884277,
11.8101100921631,34.6328620910645,
-46.8378257751465,38.0592918395996,
-58.5486145019531,10.8700113296509,
-36.8284759521484,-37.5431861877441,
-30.8832263946533,-59.9044036865234,
-44.6151199340820,-30.9810943603516,
-42.1941299438477,23.6887855529785,
-15.4696102142334,56.4039955139160,
0.230267956852913,57.6817855834961,
-13.1254014968872,55.3563385009766,
-18.5599002838135,61.0830841064453,
10.1145792007446,51.9970245361328,
30.8148860931397,18.2683162689209,
-4.95962238311768,-13.9227132797241,
-73.6190185546875,-18.2973346710205,
-95.2122879028320,-14.6967811584473,
-34.3003845214844,-29.0820140838623,
51.2994003295898,-47.2033958435059,
74.2719345092773,-33.1543350219727,
25.9512557983398,11.0824460983276,
-24.6437797546387,36.5131874084473,
-23.4955234527588,13.3621997833252,
12.7241058349609,-29.8584308624268,
27.7261848449707,-47.2497749328613,
-2.44814276695251,-27.2775135040283,
-44.6895675659180,-1.32533299922943,
-49.3107490539551,6.76103162765503,
-7.88883304595947,0.385254621505737,
39.7511558532715,-13.3684120178223,
51.6627960205078,-30.9813575744629,
33.6278228759766,-46.8193092346191,
19.5798454284668,-46.7323532104492,
23.4442424774170,-26.1788482666016,
30.7439975738525,-2.00082039833069,
18.9327888488770,5.17536878585815,
0.476427614688873,-2.00992059707642,
6.26306629180908,-9.44617366790772,
33.5523223876953,-8.09437179565430,
51.3775749206543,-3.84184670448303,
41.7729110717773,-0.640403270721436,
15.6569185256958,14.3108158111572,
-7.16031265258789,42.9987602233887,
-21.3644371032715,59.7807617187500,
-25.3517093658447,43.2936820983887,
-7.20076704025269,6.00711679458618,
31.4603729248047,-10.9693927764893,
53.9600143432617,13.4977893829346,
26.7043628692627,51.5716972351074,
-30.0523891448975,59.6323661804199,
-54.5812339782715,27.1134300231934,
-20.3875923156738,-16.5525321960449,
28.2370643615723,-39.0683746337891,
30.4793338775635,-30.5581665039063,
-8.27907276153565,0.0423364639282227,
-38.2515449523926,31.4065990447998,
-32.3173027038574,39.5817146301270,
-12.2658672332764,15.5545444488525,
-2.69547128677368,-22.5628013610840,
-7.42307853698731,-43.4143295288086,
-14.4312324523926,-34.5905799865723,
-23.6394615173340,-18.2969741821289,
-33.2775993347168,-12.0023546218872,
-25.6036128997803,-14.9243774414063,
5.63017320632935,-11.9907560348511,
34.8439903259277,-9.79537677764893,
35.6516876220703,-19.7520675659180,
22.4161376953125,-33.7477874755859,
30.7048950195313,-25.3527565002441,
58.0025787353516,5.29544544219971,
62.1589698791504,27.8545608520508,
29.1583404541016,18.4699878692627,
1.71679282188416,-8.40980720520020,
19.8966941833496,-16.3697471618652,
59.7969169616699,9.42551994323731,
56.1306838989258,54.7778587341309,
-1.63280403614044,85.3709106445313,
-53.8854179382324,75.3924560546875,
-52.1104812622070,29.8958683013916,
-17.7711791992188,-24.9383926391602,
0.721715211868286,-55.7490272521973,
-4.16911077499390,-56.3505058288574,
0.475544333457947,-46.5530166625977,
27.8535366058350,-44.2389221191406,
50.8680801391602,-37.6132125854492,
45.9294357299805,-13.9305782318115,
21.3288993835449,14.3396863937378,
-3.14496660232544,26.1858634948730,
-23.9222259521484,27.1742057800293,
-41.2376785278320,35.9452705383301,
-40.4032974243164,44.9452896118164,
-15.0268821716309,26.9537620544434,
13.4900846481323,-18.5469207763672,
17.4403190612793,-56.2643814086914,
10.1478166580200,-54.3245506286621,
23.0586891174316,-30.0479316711426,
52.5093727111816,-14.3043069839478,
57.1615791320801,-6.06482410430908,
17.1968498229980,14.9562034606934,
-29.6348457336426,40.8569068908691,
-33.1078567504883,44.1103057861328,
-3.67637681961060,28.5501384735107,
5.19054460525513,22.7150382995605,
-24.6047477722168,29.1460132598877,
-52.9141044616699,12.0349979400635,
-41.1024436950684,-30.0372161865234,
-0.0896995067596436,-44.4360122680664,
28.0783710479736,10.3528423309326,
25.4008388519287,78.9336547851563,
6.22683763504028,69.8389205932617,
-3.07979440689087,-16.3064022064209,
10.4436244964600,-75.0338058471680,
34.3700675964356,-34.0118408203125,
41.4280052185059,48.8737640380859,
13.6605777740479,69.3223800659180,
-34.9819641113281,11.4948387145996,
-62.6312599182129,-43.5337524414063,
-42.3292770385742,-38.7300453186035,
3.20422291755676,-5.73264360427856,
28.3438816070557,7.00653076171875,
22.5554199218750,8.25369930267334,
6.88245296478272,34.9523353576660,
-4.71661186218262,73.9435653686523,
-13.0322427749634,68.8159561157227,
-15.7683410644531,6.53527402877808,
-2.22869396209717,-47.1009750366211,
22.5519447326660,-31.1904621124268,
25.6969070434570,22.3184432983398,
-8.91728210449219,37.9893455505371,
-47.7127304077148,-11.5929260253906,
-46.7056045532227,-73.8774871826172,
-9.20221996307373,-82.3138198852539,
24.6781425476074,-38.6701507568359,
30.2021179199219,-0.146419167518616,
25.8810405731201,2.33272457122803,
32.6006011962891,-6.00436830520630,
37.5785408020020,2.75007629394531,
20.3175239562988,20.5287437438965,
-6.76720333099365,17.3809585571289,
-12.4099693298340,-7.75916481018066,
12.6192483901978,-18.2636108398438,
33.9486961364746,12.0857925415039,
22.1773185729980,52.6230010986328,
-11.3447980880737,53.4301109313965,
-31.1337089538574,15.8649158477783,
-18.8773174285889,-11.0455589294434,
8.83616828918457,0.251171886920929,
32.6013984680176,21.6910533905029,
51.1296234130859,17.4777870178223,
60.8534126281738,-0.426891684532166,
50.6554718017578,13.7963237762451,
13.3548278808594,56.0446090698242,
-29.7701358795166,71.0829772949219,
-46.3483848571777,30.1899414062500,
-35.9778671264648,-20.1454467773438,
-27.8409729003906,-22.9849205017090,
-41.3176307678223,7.26023387908936,
-52.0447387695313,11.4472389221191,
-30.6333312988281,-21.0133800506592,
12.6862306594849,-36.4009017944336,
42.6434020996094,-2.49531984329224,
36.6112289428711,32.8204917907715,
7.66890716552734,13.0803337097168,
-18.8423995971680,-40.4346199035645,
-31.9427127838135,-51.8307342529297,
-32.2449417114258,0.671896457672119,
-21.1918334960938,57.6941795349121,
-1.65402925014496,60.0217742919922,
16.8947563171387,21.7861766815186,
22.4165306091309,-3.01960992813110,
10.8690919876099,0.938492000102997,
-13.3500928878784,4.98889017105103,
-36.3111495971680,-0.826633810997009,
-34.7987556457520,1.61931490898132,
-4.26121425628662,19.5516510009766,
33.4001121520996,31.3291664123535,
45.0736045837402,13.8335084915161,
28.8351058959961,-14.0736885070801,
12.0991992950439,-13.9706916809082,
12.3875560760498,17.6200370788574,
7.35281181335449,42.6975593566895,
-25.4633445739746,30.4774608612061,
-66.9576873779297,-10.8207950592041,
-70.7899780273438,-49.5787048339844,
-26.5455207824707,-59.9506835937500,
24.5515003204346,-42.7511253356934,
40.2869796752930,-21.4603710174561,
24.5858249664307,-11.5969343185425,
9.73824310302734,-14.6916465759277,
13.1555881500244,-10.9233684539795,
23.7571144104004,15.6989698410034,
28.1988391876221,53.0487594604492,
23.1759796142578,67.3572082519531,
13.8436698913574,42.5469436645508,
6.54512023925781,4.41924810409546,
3.72879981994629,-10.1850481033325,
11.9946308135986,3.89965486526489,
31.5890865325928,15.3189926147461,
54.4933280944824,3.33521366119385,
63.9514007568359,-16.3625507354736,
48.3573989868164,-15.0468425750732,
10.3371963500977,1.62396144866943,
-29.1228218078613,-1.26700520515442,
-39.7425651550293,-33.8091583251953,
-16.6746597290039,-65.2827682495117,
9.42729854583740,-57.8322143554688,
2.75432276725769,-18.1218738555908,
-36.1742782592773,9.82430362701416,
-66.4934768676758,2.25201630592346,
-54.3245697021484,-14.3501520156860,
-10.4376621246338,-5.27989101409912,
25.4881343841553,24.7838764190674,
30.0938396453857,41.0028915405273,
18.1556911468506,27.8551235198975,
20.3343906402588,5.97102022171021,
43.7805175781250,-0.848744332790375,
62.9918479919434,3.86827945709229,
51.3788642883301,2.01269435882568,
9.84042739868164,-4.33264255523682,
-24.6081352233887,-3.01890563964844,
-21.0897655487061,0.828103542327881,
10.3440675735474,-9.05253791809082,
32.4655647277832,-28.7203750610352,
20.2576274871826,-33.7547111511231,
-4.28330707550049,-9.80537605285645,
-6.91545057296753,18.6863059997559,
15.1116313934326,28.3934631347656,
31.8617267608643,25.4831600189209,
22.5714149475098,34.4488830566406,
-3.85230636596680,49.3113594055176,
-18.8475284576416,37.8956832885742,
-16.5379562377930,-10.7601604461670,
-6.44309806823731,-55.7603797912598,
-1.62027394771576,-50.0716323852539,
-0.857102632522583,-0.984177589416504,
-6.16183233261108,34.2813415527344,
-14.8996887207031,12.2705106735230,
-21.2665405273438,-47.1538658142090,
-12.5855045318604,-88.5926132202148,
15.4366416931152,-79.8255767822266,
44.5003089904785,-35.6232490539551,
45.8061485290527,13.0914211273193,
14.5440502166748,45.1529846191406,
-21.3282890319824,58.1938972473145,
-25.5420970916748,49.8474388122559,
6.31614112854004,23.0810222625732,
46.1069793701172,-5.08975982666016,
62.4505729675293,-12.0451755523682,
57.0840072631836,-0.449889302253723,
49.4666137695313,5.06455326080322,
48.6372489929199,-9.65728092193604,
41.7753677368164,-28.0666923522949,
22.9544181823730,-25.6691036224365,
6.96600198745728,-9.70429515838623,
9.75220966339111,-10.1141910552979,
23.5154342651367,-32.6734733581543,
30.9242591857910,-46.7261695861816,
27.3165683746338,-30.0782814025879,
20.0990200042725,4.67128276824951,
11.4226531982422,23.2904129028320,
-8.62383651733398,21.8887634277344,
-34.5176925659180,22.7106227874756,
-47.7604522705078,28.8354530334473,
-39.7829856872559,25.4312114715576,
-26.1149063110352,5.22557687759399,
-24.6220264434814,-5.84094619750977,
-26.6020755767822,7.82760047912598,
-19.4946823120117,25.9833602905273,
-7.78084754943848,21.2275810241699,
-8.18257427215576,-1.39177346229553,
-16.2203273773193,-13.4075469970703,
-13.6481266021729,-6.12413072586060,
3.87848043441772,-2.27015590667725,
13.4051675796509,-18.4382438659668,
0.519608139991760,-37.2005615234375,
-19.7310619354248,-35.2838745117188,
-22.8954219818115,-18.3907318115234,
-14.0651464462280,-10.1687278747559,
-12.4829473495483,-22.0989360809326,
-20.3424663543701,-43.2646942138672,
-16.6122112274170,-54.4078712463379,
7.30497646331787,-46.3896903991699,
25.8557758331299,-19.1330299377441,
15.5058975219727,10.4503793716431,
-6.71710014343262,23.4189796447754,
-10.5571184158325,14.9853200912476,
11.0293712615967,3.18041229248047,
30.8802852630615,13.6594057083130,
28.2398586273193,41.7199974060059,
18.4526062011719,54.0504570007324,
29.9799575805664,30.7966403961182,
58.3061523437500,-10.7468328475952,
63.9074897766113,-33.0422821044922,
25.6405048370361,-22.7582378387451,
-28.2831764221191,3.67106008529663,
-48.3872184753418,17.0143108367920,
-17.7346343994141,6.32519006729126,
20.0962200164795,-19.7467651367188,
15.7020549774170,-42.9117774963379,
-31.7726783752441,-48.8437156677246,
-71.7103424072266,-29.5566844940186,
-63.0249443054199,4.00630187988281,
-20.0324592590332,30.8005828857422,
11.1301069259644,30.9080734252930,
9.93237781524658,5.36358547210693,
-1.74269104003906,-21.9460582733154,
7.70171737670898,-32.7311172485352,
31.4603652954102,-31.4176864624023,
41.1243133544922,-31.3946418762207,
25.1105594635010,-39.8145523071289,
8.76177024841309,-43.3595924377441,
14.6948432922363,-28.0830574035645,
38.6135749816895,-5.22336387634277,
54.7463684082031,8.00933742523193,
46.8817939758301,5.27849674224854,
24.2449321746826,0.697113215923309,
2.39305758476257,7.33995771408081,
-9.13975334167481,20.2078418731689,
-6.97273492813110,17.2900657653809,
6.66645860671997,-11.4164438247681,
25.1435375213623,-48.3195877075195,
37.3079833984375,-57.5348777770996,
35.6125450134277,-25.3909511566162,
27.4017028808594,22.3516349792480,
24.4828872680664,41.7145118713379,
27.4403610229492,18.1448040008545,
33.8208236694336,-13.6850872039795,
43.6734352111816,-10.8268384933472,
48.9841461181641,27.5676345825195,
38.3493804931641,58.3265037536621,
12.4296302795410,56.1343803405762,
-7.70351266860962,35.9681282043457,
-3.84598946571350,23.2609615325928,
15.8040494918823,21.0552005767822,
25.5180950164795,14.9515542984009,
19.5608882904053,4.68914890289307,
21.2160835266113,4.87368774414063,
36.7623443603516,14.0005283355713,
34.0122756958008,14.4029579162598,
-9.00058364868164,7.58976459503174,
-55.3867225646973,13.4924802780151,
-54.8254547119141,32.5439033508301,
-10.4792003631592,33.1938629150391,
16.9945430755615,-2.96310997009277,
-9.27022743225098,-39.4607734680176,
-59.2170982360840,-32.2272109985352,
-80.6285858154297,4.09618759155273,
-64.7936935424805,13.3536167144775,
-32.8598403930664,-20.4945983886719,
3.25088310241699,-50.4894828796387,
44.8448867797852,-28.0030822753906,
68.8343582153320,20.1404476165772,
45.0377807617188,39.1092262268066,
-9.81392478942871,18.8618164062500,
-36.3127517700195,2.26057958602905,
-6.65813636779785,12.6690807342529,
36.5341262817383,27.9188861846924,
43.0507354736328,23.3182582855225,
14.0626649856567,7.33834886550903,
-13.6228322982788,2.12176895141602,
-19.3416328430176,4.87897205352783,
-22.0811710357666,3.05880236625671,
-35.6726913452148,2.91987991333008,
-47.8429183959961,14.5344657897949,
-47.1653442382813,26.0815448760986,
-43.2646827697754,8.50956535339356,
-38.4057731628418,-36.0270004272461,
-26.5597686767578,-64.9529418945313,
-8.76957988739014,-54.9222755432129,
-0.922151982784271,-31.6685981750488,
-1.99861705303192,-25.9183712005615,
10.9582767486572,-32.8881072998047,
37.7579536437988,-24.2817745208740,
46.6771888732910,5.24018764495850,
11.6460075378418,27.9040088653564,
-37.5149002075195,20.9181747436523,
-46.6586914062500,-8.10223197937012,
-13.1963834762573,-33.9997596740723,
14.0882740020752,-45.4328727722168,
9.28487396240234,-37.8797912597656,
2.21435928344727,-13.5355186462402,
19.2350387573242,5.72331285476685,
36.7461700439453,-6.36858701705933,
29.6262760162354,-44.3319206237793,
15.8856086730957,-61.7077331542969,
27.8996772766113,-28.7790279388428,
48.4244766235352,24.1052436828613,
29.2831554412842,44.8679656982422,
-32.3489227294922,22.7590408325195,
-77.4141845703125,-2.94559764862061,
-64.8247070312500,-10.2516059875488,
-23.9441528320313,-23.9542388916016,
-1.45274150371552,-60.6379203796387,
4.76310968399048,-84.1077804565430,
22.8662223815918,-55.5023498535156,
40.9281311035156,4.79427814483643,
32.2135391235352,39.6223373413086,
7.64887142181397,26.6612415313721,
7.62051057815552,-0.479199618101120,
34.7956085205078,-10.8159866333008,
40.9913253784180,-12.5831193923950,
3.17039036750793,-19.9688720703125,
-36.9483833312988,-23.2109680175781,
-28.7985630035400,-10.8468856811523,
7.81202220916748,4.08690118789673,
16.3232917785645,-1.52653360366821,
-12.8012485504150,-21.7734146118164,
-32.3969879150391,-22.9926033020020,
-22.4585170745850,-2.48022365570068,
-13.4561367034912,14.4122018814087,
-29.3905506134033,11.3334989547730,
-49.1687927246094,2.26342391967773,
-40.2884597778320,1.75965428352356,
-11.4247827529907,14.7276687622070,
8.53796195983887,31.7114315032959,
9.26345729827881,39.4755325317383,
7.92267131805420,31.2642440795898,
8.55928516387940,2.81133031845093,
-0.315344333648682,-28.7931900024414,
-14.9719190597534,-32.3857345581055,
-14.0282602310181,-7.82793760299683,
3.24867868423462,2.27745723724365,
9.33772182464600,-33.9528503417969,
-0.349534302949905,-79.8454589843750,
0.909240722656250,-71.9858551025391,
23.2385311126709,-10.1592626571655,
42.5364265441895,31.4370708465576,
34.7339324951172,3.94517803192139,
16.6637516021729,-46.9641418457031,
21.6807632446289,-42.1877746582031,
43.7214698791504,22.2446842193604,
42.5677108764648,71.7795867919922,
8.83731937408447,53.3383255004883,
-19.6014289855957,2.39595603942871,
-18.1200389862061,-19.0205135345459,
-2.49763441085815,-3.78241872787476,
6.16256713867188,9.32072448730469,
18.8641662597656,2.60767006874084,
41.1601409912109,-3.87761735916138,
43.4926338195801,6.66800785064697,
-0.215503692626953,22.1738834381104,
-56.8799514770508,21.5048198699951,
-63.4584159851074,4.59088134765625,
-11.7103414535522,-16.4503116607666,
39.9548034667969,-26.1797542572022,
41.3557777404785,-16.7929286956787,
15.3181219100952,11.9473161697388,
9.93005752563477,37.9557952880859,
29.7438278198242,26.1648807525635,
42.7337684631348,-21.0036888122559,
41.8631401062012,-50.8864440917969,
41.2930145263672,-24.8885269165039,
39.4572219848633,32.7928886413574,
19.8875923156738,59.3604850769043,
-16.3440952301025,34.7821235656738,
-40.0434722900391,3.25227069854736,
-31.6903190612793,4.32806777954102,
-9.51882743835449,23.0998668670654,
3.42792797088623,20.6149330139160,
11.0906972885132,-0.451551258563995,
22.0832042694092,-5.08376836776733,
25.4129428863525,15.9222965240479,
7.14606475830078,28.6875381469727,
-10.9859533309937,7.98833227157593,
-0.780304908752441,-22.8931446075439,
28.5551319122314,-24.3667373657227,
30.2845516204834,6.28352737426758,
-7.59723567962647,34.0342140197754,
-42.5592803955078,30.1521358489990,
-29.9267692565918,3.89609670639038,
9.91950225830078,-10.6450929641724,
23.0651264190674,5.14948701858521,
-2.53050994873047,31.3752460479736,
-19.7571430206299,43.7347335815430,
9.92421150207520,36.9302940368652,
55.1247329711914,26.5722618103027,
57.6081619262695,28.2512779235840,
10.9961385726929,34.8749923706055,
-32.1160469055176,25.8687515258789,
-22.6019229888916,1.22745943069458,
26.2576522827148,-16.3191833496094,
61.0500373840332,-13.8281421661377,
51.7632827758789,-4.18311643600464,
20.2735118865967,-0.938093245029450,
3.20961189270020,1.58468556404114,
3.30570435523987,22.9534931182861,
-0.770931184291840,60.6528358459473,
-16.0844688415527,77.7288131713867,
-23.7512550354004,54.8245811462402,
-5.98300790786743,19.7290954589844,
24.0057296752930,15.5258579254150,
29.9925651550293,39.0605659484863,
-1.49350810050964,49.3307800292969,
-41.2037734985352,17.2048435211182,
-52.9714546203613,-26.1140518188477,
-36.3758277893066,-30.9651546478272,
-16.5696258544922,-1.51528859138489,
-11.3017911911011,8.49739646911621,
-10.7938776016235,-23.0638160705566,
1.11184859275818,-57.0152893066406,
13.9349079132080,-39.8639450073242,
15.0130891799927,17.1925735473633,
9.39262771606445,51.3269500732422,
12.2521896362305,35.6775894165039,
24.2313766479492,12.9193248748779,
23.6871814727783,27.4714050292969,
0.876783907413483,51.0983085632324,
-23.8141098022461,29.4499435424805,
-23.8464279174805,-32.6441993713379,
-0.703033685684204,-61.7632369995117,
16.3673858642578,-14.8586912155151,
8.96810150146484,56.8021049499512,
-13.1737775802612,65.0519256591797,
-22.8785781860352,-1.45587706565857,
-4.99260759353638,-66.8682785034180,
24.0689067840576,-65.1661300659180,
36.9150810241699,-14.7910060882568,
16.4802742004395,19.6398258209229,
-26.1364707946777,8.74297523498535,
-55.7014122009277,-15.1011219024658,
-46.4353675842285,-14.3543930053711,
-9.07788276672363,0.344446003437042,
21.0819454193115,-6.11256790161133,
20.8031425476074,-39.2549743652344,
2.78246164321899,-63.9785842895508,
-7.39098072052002,-54.7723312377930,
-5.26096296310425,-21.0885124206543,
-12.1101522445679,4.69155883789063,
-35.4218101501465,6.56626796722412,
-45.4464302062988,-3.05740356445313,
-15.0939245223999,-12.9342641830444,
36.0958671569824,-25.4022903442383,
52.0909576416016,-31.5164470672607,
12.1523494720459,-15.8317403793335,
-38.0533256530762,16.4503479003906,
-42.4333534240723,31.8560199737549,
-7.73877620697022,3.61293935775757,
12.6412582397461,-36.9269027709961,
-1.43327486515045,-34.3556632995606,
-11.7138099670410,16.5449314117432,
13.8268985748291,55.6624259948731,
48.8644294738770,30.0145530700684,
43.4923324584961,-37.1435279846191,
1.90221166610718,-79.0269088745117,
-19.2695007324219,-64.1285781860352,
8.18733787536621,-28.2895927429199,
50.4830436706543,-11.3294963836670,
56.9673004150391,-16.2336044311523,
24.0884418487549,-21.5983810424805,
-10.3458175659180,-15.7000570297241,
-17.7950305938721,-1.53293025493622,
-4.83443975448608,18.3289031982422,
9.52059078216553,40.5431709289551,
23.5344810485840,48.1786155700684,
39.9669036865234,28.3406734466553,
52.5806884765625,-4.28020477294922,
46.1432342529297,-19.0108947753906,
17.7397384643555,-4.06126785278320,
-15.1528930664063,16.4102954864502,
-21.5981807708740,18.3120841979980,
9.10669612884522,13.1935853958130,
47.1866836547852,25.9868736267090,
51.1401367187500,47.5353813171387,
15.4367218017578,49.9142570495606,
-23.9151458740234,16.9206104278564,
-30.0017261505127,-19.5596504211426,
-7.45207643508911,-23.3418788909912,
7.79276561737061,1.00544476509094,
2.68919348716736,16.8176555633545,
-6.75058937072754,7.00139379501343,
-8.21107578277588,-11.2182769775391,
-14.0675573348999,-17.3207740783691,
-32.8743667602539,-12.3686800003052,
-46.7486801147461,-9.75743198394775,
-42.3078422546387,-13.1885290145874,
-29.3365459442139,-22.5706882476807,
-28.7895088195801,-42.6782722473145,
-29.8297271728516,-67.2397232055664,
-8.09837913513184,-69.1907119750977,
30.8372364044189,-26.9429607391357,
52.1240234375000,30.6631317138672,
37.7640419006348,50.4487304687500,
7.97234916687012,20.3880271911621,
-6.07846593856812,-10.5735979080200,
-6.93016004562378,-4.45433759689331,
-13.2807712554932,12.9086904525757,
-24.5991001129150,-4.77703952789307,
-23.5458736419678,-49.1433715820313,
-9.69078254699707,-68.0471267700195,
9.04190921783447,-38.6925888061523,
29.1997356414795,2.26065063476563,
53.6174812316895,17.1665878295898,
64.7934875488281,13.5188694000244,
41.8028144836426,21.1315803527832,
-4.95685720443726,33.7715072631836,
-28.4250106811523,28.5228500366211,
-4.20444393157959,2.72525167465210,
28.5689201354980,-12.4800338745117,
15.4650392532349,-3.00562715530396,
-35.4743194580078,15.3494758605957,
-61.9460144042969,20.1970443725586,
-38.6184425354004,1.05142688751221,
-9.93373870849609,-25.7889881134033,
-22.1029167175293,-37.7475700378418,
-57.7222671508789,-24.3274345397949,
-64.4689407348633,2.15921235084534,
-33.9629974365234,11.3543443679810,
-7.38708543777466,-15.5181236267090,
-7.79174041748047,-55.7093544006348,
-8.09403705596924,-70.1760940551758,
13.8129329681396,-53.4797401428223,
35.7934341430664,-36.2795524597168,
22.2769927978516,-37.3878860473633,
-12.2815103530884,-36.1232719421387,
-25.8535156250000,-17.2990036010742,
-9.34329223632813,-3.57074260711670,
5.95122051239014,-21.6841945648193,
3.53073453903198,-56.0522537231445,
-0.215880468487740,-62.5671844482422,
13.4075546264648,-27.2102260589600,
32.0588188171387,15.9956293106079,
30.7142066955566,33.7199440002441,
14.2526741027832,30.7977733612061,
4.18343019485474,22.3766231536865,
-1.86420226097107,9.24123191833496,
-9.07415771484375,-6.97772121429443,
-8.58596611022949,-10.0569982528687,
10.8075361251831,7.45065546035767,
34.4855766296387,18.3866691589355,
39.1088790893555,0.499985158443451,
31.4380264282227,-21.6529655456543,
37.6637115478516,-6.34802436828613,
53.2088470458984,36.6282730102539,
36.0112609863281,55.0391960144043,
-24.9824981689453,23.5161552429199,
-68.7706756591797,-16.1696109771729,
-38.4074935913086,-15.9458818435669,
24.6654319763184,16.9679050445557,
28.5886707305908,31.5049266815186,
-40.5265617370606,9.90337467193604,
-95.7225036621094,-20.4113960266113,
-69.6707458496094,-28.4136981964111,
-2.78529214859009,-10.4711923599243,
19.5561828613281,23.2494392395020,
-12.3962564468384,53.1367492675781,
-32.9719848632813,54.9676666259766,
-9.72305774688721,23.7508602142334,
19.2544746398926,-6.30099296569824,
14.0700445175171,0.712125658988953,
-4.73421525955200,37.2021713256836,
-4.76947116851807,55.9910316467285,
2.71801972389221,36.7068290710449,
-12.2648849487305,10.0069837570190,
-34.4414062500000,13.3706884384155,
-22.5667839050293,29.7523269653320,
16.5873737335205,24.2987327575684,
31.9642410278320,5.32612752914429,
1.57198619842529,9.76268959045410,
-31.6096019744873,33.2534675598145,
-19.6623878479004,36.6480636596680,
23.5548381805420,12.0548334121704,
43.7497940063477,-1.50379192829132,
25.7890300750732,22.5218868255615,
0.0747718811035156,54.6557388305664,
-10.8144187927246,56.2247467041016,
-9.53227806091309,36.2363739013672,
-0.854196190834045,28.3369274139404,
17.6298332214355,34.5914077758789,
39.6497764587402,26.6342849731445,
45.2561454772949,-1.80553722381592,
23.8659629821777,-19.0700969696045,
-2.61925792694092,-15.5634946823120,
-10.3429431915283,-18.0512409210205,
-2.68067121505737,-33.4041671752930,
6.10430526733398,-33.2475738525391,
18.9622917175293,1.41737675666809,
40.9997978210449,36.9623489379883,
47.4922752380371,31.8000068664551,
19.1611499786377,-9.83052158355713,
-20.4301967620850,-43.4037513732910,
-25.7819366455078,-49.0908279418945,
7.34986400604248,-43.0307159423828,
29.9168262481689,-34.5663375854492,
11.2776126861572,-7.54227924346924,
-11.3780117034912,33.0764389038086,
9.14638710021973,51.5818328857422,
53.8453788757324,30.3919277191162,
59.3683700561523,8.80845737457275,
12.1292037963867,30.5747528076172,
-28.6509895324707,76.2954788208008,
-20.3970108032227,92.7878494262695,
8.23402976989746,63.1259498596191,
2.64773178100586,25.7130966186523,
-34.9914093017578,17.8855533599854,
-53.4209594726563,31.6401462554932,
-32.8108177185059,32.3315887451172,
-3.22888660430908,10.4961662292480,
3.00626516342163,-13.9622287750244,
-6.71214246749878,-23.4829387664795,
-8.83382320404053,-12.6672534942627,
-9.95295429229736,5.59179639816284,
-27.6878757476807,9.91835880279541,
-48.8883056640625,-14.6827087402344,
-43.0514602661133,-45.4443893432617,
-12.5868425369263,-40.0521278381348,
1.61593294143677,3.48493099212647,
-21.3010139465332,38.2412261962891,
-56.1762504577637,22.2216453552246,
-56.0697937011719,-20.5839500427246,
-9.98185157775879,-31.4420223236084,
41.9354667663574,4.20371961593628,
58.1540641784668,30.2744560241699,
33.5140838623047,10.0534505844116,
-5.75532674789429,-21.5930233001709,
-30.5522480010986,-17.9014873504639,
-32.1096992492676,6.01538705825806,
-19.5645942687988,-1.48773169517517,
-10.9917449951172,-44.8313674926758,
-8.42105960845947,-63.0595054626465,
-5.35729265213013,-19.3708305358887,
-2.02410864830017,41.3535652160645,
-13.2827863693237,53.4940109252930,
-36.4285278320313,21.2445354461670,
-47.2421989440918,1.65163624286652,
-25.6301174163818,20.0332183837891,
14.6627321243286,35.0406761169434,
36.6304130554199,9.93879985809326,
29.3315544128418,-26.8069114685059,
18.0948810577393,-27.9369335174561,
18.3822917938232,2.25090169906616,
6.62242412567139,18.4587612152100,
-31.4395408630371,-0.384581089019775,
-66.4151229858398,-27.4772644042969,
-61.8539199829102,-30.5625057220459,
-30.9107532501221,-12.7128190994263,
-17.6939010620117,0.545178771018982,
-31.5992908477783,0.880692243576050,
-36.1704559326172,-4.89780807495117,
-11.6533937454224,-12.6315841674805,
8.25353145599365,-18.4980869293213,
-11.3143796920776,-10.7089157104492,
-46.1246566772461,6.47891950607300,
-53.8589477539063,12.0081415176392,
-35.0360488891602,-6.52506208419800,
-30.8193626403809,-26.7633781433105,
-50.0604782104492,-18.9291324615479,
-48.5237884521484,11.7165908813477,
-2.96415805816650,27.7595062255859,
45.6781692504883,16.6278057098389,
45.7088699340820,9.61262893676758,
9.81330204010010,31.4590358734131,
-9.43809604644775,61.3651237487793,
11.3834619522095,64.4036254882813,
33.6652259826660,40.5635261535645,
16.2957668304443,21.5051536560059,
-22.3258476257324,17.4239978790283,
-30.3930263519287,7.97252178192139,
4.84219264984131,-16.4617881774902,
44.8744659423828,-34.3734359741211,
46.1490592956543,-24.1368293762207,
9.87796783447266,4.49934291839600,
-25.1937847137451,15.4869184494019,
-23.6478805541992,-6.78004360198975,
4.89749288558960,-38.2851448059082,
20.9936885833740,-44.9076652526856,
-0.830557703971863,-16.8701019287109,
-37.6474647521973,21.9704971313477,
-44.2822113037109,33.2340545654297,
0.713681697845459,1.61252188682556,
56.3330841064453,-40.1748161315918,
65.1943359375000,-41.4509811401367,
18.4106998443604,2.51399683952332,
-30.7735309600830,39.6707878112793,
-39.0976295471191,22.4914970397949,
-19.0798587799072,-27.1460018157959,
-13.3540325164795,-43.7849731445313,
-28.7376785278320,-3.47414922714233,
-34.0810661315918,41.2755050659180,
-11.9797315597534,29.1432971954346,
7.97989463806152,-22.0679283142090,
-0.225053668022156,-48.4902496337891,
-20.0975704193115,-29.5436744689941,
-12.1666069030762,-7.75837326049805,
25.2840385437012,-14.3345289230347,
55.5753364562988,-33.5907440185547,
52.0926322937012,-34.5281867980957,
32.7959060668945,-24.8512039184570,
25.9514579772949,-29.7447929382324,
38.5732688903809,-37.8898811340332,
58.7714729309082,-19.0084171295166,
64.2682037353516,20.7681598663330,
39.8807029724121,40.2202033996582,
-3.44845557212830,28.1800308227539,
-36.7841186523438,22.0851364135742,
-39.7513694763184,45.0107002258301,
-25.9367847442627,62.6271095275879,
-32.7939186096191,38.8254852294922,
-61.9064559936523,4.29354381561279,
-69.2101440429688,11.1664943695068,
-30.7368545532227,50.6139755249023,
8.69333267211914,57.5934982299805,
-2.68200469017029,7.46577453613281,
-41.9432373046875,-42.1138648986816,
-47.7674369812012,-31.3814907073975,
-7.17285442352295,13.1934413909912,
17.3180809020996,23.2299003601074,
-7.64304590225220,-13.1616859436035,
-39.6710281372070,-41.1030044555664,
-23.0329322814941,-26.4999618530273,
13.0204620361328,1.80161142349243,
3.87404918670654,5.33772945404053,
-54.6186408996582,-15.9836807250977,
-92.1742630004883,-31.8681774139404,
-66.3283843994141,-31.3911113739014,
-20.5383758544922,-25.6367435455322,
-12.3362569808960,-24.3100204467773,
-31.9941787719727,-21.4047183990479,
-30.3716049194336,-17.0336742401123,
6.82871627807617,-17.2774600982666,
49.0165367126465,-15.6575498580933,
68.1260147094727,-0.735444784164429,
64.2541122436523,13.8394031524658,
56.2204742431641,11.9009571075439,
50.7194976806641,1.26123797893524,
47.9078407287598,5.98124933242798,
50.5446662902832,28.5058555603027,
53.1689109802246,39.1973800659180,
41.1244773864746,14.5327529907227,
18.3647632598877,-21.2755870819092,
2.94884228706360,-32.5275459289551,
-3.44523406028748,-21.2461681365967,
-23.9720020294189,-17.1892890930176,
-57.4646606445313,-19.9085121154785,
-72.9179992675781,-4.15438842773438,
-46.8621673583984,31.1203441619873,
-7.87512683868408,43.3388023376465,
-4.97879791259766,8.54923248291016,
-36.1097412109375,-35.2906532287598,
-46.0404281616211,-35.8740501403809,
-12.1603345870972,3.72077918052673,
26.7018070220947,27.7803897857666,
20.1778697967529,5.92317008972168,
-16.7172698974609,-32.3044281005859,
-36.8513793945313,-43.9050903320313,
-26.5649013519287,-28.3511962890625,
-19.5199356079102,-15.0807485580444,
-30.4263210296631,-13.0903263092041,
-33.1983375549316,-5.52458143234253,
-5.19159555435181,13.3428173065186,
27.2646255493164,29.4008674621582,
24.1213703155518,27.0249214172363,
-15.6626071929932,10.3036880493164,
-49.3561630249023,-7.53909301757813,
-38.8055000305176,-19.7812805175781,
0.476476907730103,-28.0371932983398,
33.0930709838867,-32.5443992614746,
43.1615486145020,-30.8029689788818,
34.2851562500000,-24.7780666351318,
22.4870090484619,-18.7733287811279,
14.9545001983643,-14.6507129669189,
5.17645168304443,-13.3311395645142,
-5.69794654846191,-18.7879600524902,
-5.44463729858398,-26.6066837310791,
10.9773874282837,-24.0564346313477,
27.4211044311523,-7.66942548751831,
12.9350566864014,10.0483503341675,
-33.1208877563477,12.8494434356689,
-69.7280502319336,1.36144649982452,
-45.8382682800293,-5.38502073287964,
27.4135627746582,4.35530281066895,
72.4892883300781,20.6874771118164,
32.5672683715820,27.5613460540772,
-52.3625183105469,21.7401161193848,
-92.3157043457031,9.51936054229736,
-44.9319610595703,-7.83567762374878,
33.2988967895508,-28.2153167724609,
63.2031250000000,-31.9673099517822,
35.7057533264160,-0.514697492122650,
-1.08872544765472,52.2611198425293,
-15.8909454345703,79.0409011840820,
-23.7608432769775,45.8229751586914,
-36.0070915222168,-25.9342155456543,
-31.0441761016846,-78.0461807250977,
9.90970706939697,-70.5206222534180,
56.3395576477051,-18.4154720306397,
55.4602088928223,30.6339225769043,
8.01930522918701,41.3414154052734,
-23.1490077972412,14.8065958023071,
2.76686930656433,-15.8614273071289,
50.3559417724609,-19.0380344390869,
52.6632080078125,11.3840675354004,
-3.59652256965637,45.9440536499023,
-60.8983230590820,54.3151245117188,
-63.5515441894531,34.7191886901856,
-28.5209693908691,15.8186244964600,
-9.79204654693604,15.4324502944946,
-28.9101924896240,21.5532913208008,
-52.2665328979492,13.4726867675781,
-38.4555282592773,-12.8170957565308,
5.86333894729614,-31.3107643127441,
36.9628181457520,-25.7726993560791,
26.8839035034180,-8.76007652282715,
-4.37200880050659,0.183303043246269,
-17.6554508209229,-10.8561258316040,
-5.39473438262939,-31.9444370269775,
11.9471340179443,-45.3860359191895,
18.7544574737549,-43.7647171020508,
20.6588497161865,-31.3141307830811,
30.3050918579102,-17.2458114624023,
37.7279357910156,-12.5691833496094,
20.5941848754883,-15.9057855606079,
-14.6583528518677,-15.5289077758789,
-36.0797920227051,4.19599103927612,
-22.8082237243652,33.3431701660156,
5.28454589843750,45.5020065307617,
17.8930702209473,27.6853694915772,
9.06945896148682,6.23342418670654,
-4.80704784393311,16.6518535614014,
-16.0375728607178,54.1402168273926,
-27.3565292358398,72.3786163330078,
-28.3069744110107,43.9579086303711,
-6.22041082382202,1.22121596336365,
31.4106388092041,-4.05901765823364,
51.6985130310059,23.9762229919434,
38.0239639282227,34.3231391906738,
15.6561021804810,11.0627384185791,
13.0820140838623,-7.65294408798218,
17.1670379638672,13.0434837341309,
3.43193292617798,48.6080780029297,
-17.1804828643799,50.8088989257813,
-12.6693086624146,19.2474098205566,
14.3216371536255,-0.957711756229401,
29.0769882202148,9.05284118652344,
16.9096794128418,28.4123325347900,
7.76501941680908,33.0258255004883,
21.3822746276855,30.7126007080078,
27.8895797729492,27.2686614990234,
-5.11865663528442,9.34563636779785,
-45.5817413330078,-25.7060947418213,
-36.6910171508789,-41.1316184997559,
12.6395568847656,-11.1029663085938,
30.6820526123047,33.3585395812988,
-13.3398094177246,40.1567077636719,
-60.5669441223145,6.20037841796875,
-48.1457557678223,-22.0772380828857,
1.43724787235260,-7.37071895599365,
18.5081291198730,30.2038440704346,
-12.2562789916992,50.5600090026856,
-39.8424072265625,47.3789863586426,
-32.1758346557617,39.0954208374023,
-16.7066040039063,30.9178066253662,
-23.7410182952881,15.6422567367554,
-30.9807262420654,-4.57793903350830,
-7.82562255859375,-22.1657676696777,
25.3350830078125,-29.5470333099365,
23.9246196746826,-22.9955577850342,
-10.3742904663086,-0.823321938514710,
-26.9300346374512,27.2632732391357,
-0.183172821998596,32.0006027221680,
36.7476615905762,-0.827433347702026,
41.2164878845215,-46.7789459228516,
14.6091918945313,-59.8463516235352,
-6.21445655822754,-31.3452434539795,
-1.33119201660156,-6.16458463668823,
13.0392560958862,-20.3374462127686,
17.0593776702881,-46.1101608276367,
12.0376205444336,-35.8773574829102,
4.30719041824341,12.6158781051636,
-5.76788902282715,41.3502464294434,
-17.4559020996094,12.5364522933960,
-21.5582485198975,-46.1863136291504,
-11.5458698272705,-73.6138000488281,
8.89306163787842,-47.1614990234375,
19.6883640289307,0.787886321544647,
5.09626579284668,30.6059207916260,
-24.0648231506348,35.5588569641113,
-37.6444854736328,29.8846073150635,
-20.4464912414551,26.6089076995850,
13.3995847702026,22.1409778594971,
28.0605201721191,17.7599601745605,
3.57379889488220,20.0364818572998,
-29.6177368164063,28.8086414337158,
-26.6676406860352,38.8902015686035,
13.2855491638184,41.0492591857910,
42.5104255676270,32.1709938049316,
21.8642406463623,21.2393360137939,
-28.9624786376953,20.7031650543213,
-55.8791122436523,24.4017200469971,
-42.4005775451660,18.1691398620605,
-24.8080978393555,-4.66252660751343,
-36.4117431640625,-34.7643470764160,
-47.5801582336426,-51.2600517272949,
-14.0352249145508,-52.6697158813477,
48.0322608947754,-54.3703727722168,
69.3839874267578,-59.0949630737305,
19.3322467803955,-49.9029273986816,
-44.6686019897461,-14.6186809539795,
-48.6011009216309,19.7038097381592,
0.274645328521729,23.1460990905762,
28.9667644500732,9.45756340026856,
4.15008258819580,14.5785226821899,
-29.5636100769043,45.2228393554688,
-24.3647117614746,64.1760482788086,
-3.90577125549316,44.5342636108398,
-19.4654998779297,4.93287277221680,
-62.8352394104004,-20.1441898345947,
-72.9540634155273,-31.1641559600830,
-29.4703540802002,-43.8103141784668,
21.8619441986084,-46.9497146606445,
28.8107719421387,-21.4318866729736,
-2.99179840087891,10.1306285858154,
-33.0582466125488,-0.731497347354889,
-37.8884620666504,-45.1350479125977,
-22.6863422393799,-57.9387512207031,
1.25245630741119,-3.92072534561157,
21.6945438385010,53.8036231994629,
16.7985286712647,44.7285079956055,
-18.5587882995605,-12.8592586517334,
-47.0377311706543,-37.8615493774414,
-34.3403701782227,-3.79747653007507,
0.580157458782196,33.0819511413574,
12.0184068679810,18.7992668151855,
-7.23492765426636,-15.2744455337524,
-20.1009693145752,-17.7472724914551,
-11.9999074935913,5.50897693634033,
-10.0505332946777,11.8581047058105,
-37.4014587402344,-9.41527938842773,
-54.6293373107910,-23.6000576019287,
-18.6796798706055,-10.1217451095581,
39.1148910522461,19.4831485748291,
47.4104309082031,45.0661773681641,
1.25087261199951,57.4423370361328,
-34.0704307556152,51.3396415710449,
-17.3379955291748,27.6502494812012,
15.4465065002441,3.54223251342773,
15.2752246856689,8.45762634277344,
-4.20780181884766,42.6416397094727,
-3.55475783348084,62.7016639709473,
13.5139513015747,44.0735969543457,
1.30173873901367,13.4785041809082,
-45.8789672851563,1.54310441017151,
-79.7799758911133,-3.72717308998108,
-66.3365554809570,-22.8284111022949,
-30.5611267089844,-42.7527999877930,
-10.9368648529053,-30.7341709136963,
-4.05361461639404,5.48962354660034,
14.2292194366455,17.3238754272461,
31.1684589385986,-10.9241523742676,
20.5536289215088,-30.5976276397705,
-13.1966438293457,-5.54277467727661,
-34.8750228881836,26.3010940551758,
-26.6230373382568,9.68276596069336,
-8.80683517456055,-40.8336105346680,
-13.0020322799683,-54.1958656311035,
-37.7943649291992,-13.0836009979248,
-53.2219848632813,16.9827175140381,
-40.2520446777344,-15.5381307601929,
-5.90886783599854,-71.0470809936523,
29.2729072570801,-73.6682662963867,
39.4265594482422,-17.4457073211670,
13.8923473358154,30.4171695709229,
-16.9293785095215,20.3450050354004,
-14.7729101181030,-16.9610691070557,
21.0487537384033,-21.4095630645752,
49.3808670043945,10.5094537734985,
40.9819793701172,37.8164634704590,
19.6609363555908,33.7020912170410,
24.3238391876221,10.4039745330811,
42.7799415588379,-4.66032028198242,
27.1454162597656,-5.28987360000610,
-24.5818939208984,-7.03029394149780,
-49.6748504638672,-26.5651569366455,
-5.12294292449951,-50.1731605529785,
56.9375457763672,-47.0126037597656,
61.4514083862305,-0.633214354515076,
8.50393390655518,57.1855964660645,
-27.6761951446533,76.5312728881836,
-4.56982564926148,36.2185707092285,
33.6889305114746,-14.4832286834717,
28.7587909698486,-12.8984012603760,
-7.78542947769165,32.7956199645996,
-18.3110771179199,55.2049407958984,
12.2826404571533,19.2891502380371,
42.5805625915527,-35.8142967224121,
34.8993835449219,-52.3881607055664,
4.04514598846436,-26.1486701965332,
-22.0812950134277,-2.97138118743897,
-40.1073951721191,-5.95246219635010,
-54.5203628540039,-19.7498207092285,
-51.2564620971680,-32.6421546936035,
-22.0946540832520,-52.9832420349121,
7.98483657836914,-74.1650543212891,
7.47539854049683,-64.4224090576172,
-20.7344455718994,-14.4679145812988,
-31.6805381774902,31.0340023040772,
-1.22663831710815,22.6030941009522,
39.2679290771484,-18.3855609893799,
46.0967636108398,-33.8762435913086,
20.7186412811279,-8.44948387145996,
-6.99504804611206,16.2835597991943,
-17.2590484619141,3.95186853408813,
-11.3019008636475,-28.4323997497559,
1.72423601150513,-38.9630775451660,
11.1658916473389,-21.1959743499756,
10.0538959503174,3.03260278701782,
0.117976859211922,22.7210407257080,
-0.946774184703827,36.4675331115723,
17.6085720062256,32.5303344726563,
37.8793563842773,6.53785514831543,
33.3809432983398,-16.9367141723633,
7.80231571197510,-5.49265575408936,
-2.59246826171875,28.0333938598633,
20.2694721221924,34.1919860839844,
44.9156112670898,-0.256621837615967,
41.9080657958984,-29.3697261810303,
21.9946384429932,-8.21291446685791,
12.4230051040649,34.9585342407227,
16.8564643859863,32.7711944580078,
15.0101442337036,-21.5654773712158,
0.0857468247413635,-62.8852043151856,
-14.2251958847046,-46.1159019470215,
-14.9796380996704,-4.36689996719360,
-4.75919771194458,9.00530719757080,
13.3477973937988,-7.80950164794922,
37.4001274108887,-9.08972454071045,
51.3458251953125,20.9767017364502,
27.6604652404785,51.0945701599121,
-26.3368778228760,53.7313804626465,
-62.8068809509277,41.5925140380859,
-51.1213874816895,35.7799568176270,
-17.8156356811523,33.0457878112793,
-5.09542655944824,14.7110710144043,
-14.3147382736206,-12.0476016998291,
-16.2687225341797,-22.5953674316406,
-3.38189244270325,-16.6122570037842,
-8.34333610534668,-13.0609807968140,
-37.9095115661621,-14.9294214248657,
-54.2016754150391,-8.56057643890381,
-27.3555507659912,15.1975536346436,
11.1087312698364,37.8925590515137,
3.11734747886658,32.6921386718750,
-45.5755577087402,5.11863994598389,
-72.1993560791016,-13.7063350677490,
-40.8577308654785,-2.38683748245239,
2.49774575233459,29.6966018676758,
-1.78636431694031,55.8579826354981,
-43.7485389709473,47.0081939697266,
-59.4267845153809,5.20525550842285,
-12.6539363861084,-40.0683250427246,
53.9666519165039,-48.5018959045410,
71.0679855346680,-16.9827346801758,
22.5471801757813,12.6475658416748,
-35.3837242126465,-1.66430544853210,
-47.4656333923340,-49.2197647094727,
-8.54800128936768,-75.7560043334961,
38.8392601013184,-47.7594718933106,
55.8849372863770,5.58889198303223,
42.3249816894531,28.9035530090332,
29.1113090515137,12.4378643035889,
28.1306571960449,-4.84551715850830,
18.6854820251465,5.05996370315552,
-5.74268770217896,33.0487976074219,
-20.3815021514893,51.5055160522461,
-0.666576385498047,46.6975440979004,
31.7421131134033,32.1707954406738,
24.4929275512695,17.1151294708252,
-35.6500244140625,6.53589487075806,
-84.7940063476563,1.95858287811279,
-59.5469055175781,-3.08582067489624,
9.14087104797363,-18.3123550415039,
41.9630355834961,-41.0911064147949,
11.9512834548950,-45.5188102722168,
-21.7862796783447,-9.34622001647949,
-3.92901301383972,42.0488433837891,
35.5253944396973,51.7955665588379,
30.7632369995117,3.73414492607117,
-14.9552564620972,-47.8033676147461,
-36.9561958312988,-41.7828674316406,
-4.71989059448242,16.5107746124268,
31.3427410125732,66.7235107421875,
16.2323303222656,67.0636062622070,
-24.3797683715820,35.6279182434082,
-24.0474128723145,11.2030096054077,
28.4060115814209,7.30399036407471,
75.8781051635742,9.29328536987305,
69.7226486206055,7.37575912475586,
28.8556594848633,1.71548712253571,
-5.81924629211426,-10.8621807098389,
-17.0907516479492,-30.4652976989746,
-17.2925968170166,-48.3959808349609,
-14.0786619186401,-55.0119132995606,
-6.16524505615234,-48.8730697631836,
0.231351703405380,-29.0770626068115,
-3.30664110183716,-0.356816053390503,
-4.88781070709229,21.2709484100342,
14.6332607269287,13.7317485809326,
42.1638450622559,-19.4635105133057,
40.4986267089844,-41.5899810791016,
2.05410194396973,-17.3426361083984,
-37.6907386779785,23.2956809997559,
-45.7171440124512,25.8289489746094,
-29.9842853546143,-16.9308471679688,
-21.5021362304688,-50.5896682739258,
-26.6836910247803,-37.4512405395508,
-18.6571598052979,-11.6656074523926,
8.49049282073975,-20.5416107177734,
30.1644954681397,-48.8306236267090,
26.4286975860596,-39.0863113403320,
11.4157257080078,19.5875968933105,
5.39243268966675,71.7919921875000,
9.23959827423096,67.6854171752930,
15.2845048904419,32.8082504272461,
20.2075634002686,21.7262763977051,
23.4005279541016,45.3958473205566,
15.0465993881226,66.3086166381836,
-6.48876428604126,59.6948699951172,
-24.8264369964600,33.1227073669434,
-22.0287303924561,1.52547264099121,
-0.890813469886780,-30.2186622619629,
11.9849376678467,-48.2543678283691,
9.22685623168945,-37.5157661437988,
0.726300716400147,-7.71195983886719,
-12.6593313217163,8.38185214996338,
-44.3802108764648,-7.78069972991943,
-80.1169586181641,-26.7215404510498,
-78.7840347290039,-15.6971416473389,
-27.8846054077148,14.4292888641357,
29.7290420532227,21.6293983459473,
45.4196434020996,5.27964830398560,
24.5626678466797,8.74034404754639,
7.49434185028076,42.9613647460938,
4.17688465118408,67.5262908935547,
-12.6813087463379,53.3065643310547,
-47.2831954956055,23.1056766510010,
-62.3646278381348,21.8954639434814,
-35.7279319763184,41.6200103759766,
-7.13858699798584,35.2004089355469,
-13.3848381042480,-4.38004922866821,
-32.1173744201660,-34.0092735290527,
-19.4994792938232,-20.8894424438477,
18.6711158752441,10.0608110427856,
37.0743522644043,28.1748695373535,
20.3334960937500,35.7670021057129,
4.17641925811768,44.4083671569824,
10.5752992630005,37.1344757080078,
18.1867370605469,4.08813667297363,
2.94651365280151,-21.3192405700684,
-13.7118320465088,-0.135932207107544,
-7.17750644683838,47.5693511962891,
-0.140355050563812,61.0137634277344,
-26.3238334655762,17.6650886535645,
-65.3969039916992,-29.8145503997803,
-63.8317871093750,-34.4628868103027,
-21.1498432159424,-15.9852190017700,
10.3530111312866,-22.9149570465088,
-1.00715970993042,-52.7443389892578,
-23.5848445892334,-65.8304443359375,
-20.6128826141357,-46.4158859252930,
-9.59627628326416,-12.0433349609375,
-25.9858398437500,14.6942205429077,
-54.0151748657227,28.5777053833008,
-41.9870376586914,27.2359313964844,
12.2746267318726,7.88478803634644,
52.3755226135254,-6.11470890045166,
43.8953971862793,12.0674057006836,
16.8592662811279,56.7148551940918,
10.3681745529175,80.9925765991211,
15.0663881301880,53.8814239501953,
0.274050951004028,11.8099784851074,
-25.5948867797852,3.59508800506592,
-27.0508899688721,24.7236442565918,
5.23587846755981,27.3360996246338,
31.1227188110352,-8.34039402008057,
25.6893138885498,-48.5980987548828,
7.74235534667969,-54.7625389099121,
8.40044593811035,-20.4303894042969,
20.4568576812744,19.3249702453613,
18.7973117828369,32.7809600830078,
5.43882083892822,10.0241613388062,
3.85829687118530,-33.6287117004395,
15.7737798690796,-62.9441795349121,
19.6624622344971,-49.5227584838867,
2.93169307708740,-1.82279264926910,
-16.8581409454346,40.1597862243652,
-14.8152208328247,44.7777481079102,
-0.634574115276337,33.2785644531250,
-3.86814117431641,36.5279426574707,
-34.7012519836426,46.8236274719238,
-68.5887374877930,29.2607975006104,
-77.7146987915039,-21.6179332733154,
-55.3948554992676,-66.1604003906250,
-12.2410840988159,-64.6546478271484,
30.3158111572266,-26.5835380554199,
53.9987907409668,0.232492983341217,
54.5599822998047,-2.54543805122376,
45.6956939697266,-16.6000576019287,
39.0204429626465,-19.8579235076904,
34.6886711120606,-8.09667778015137,
21.5712890625000,15.8460559844971,
-3.17283797264099,47.7949905395508,
-22.2809562683105,74.1704025268555,
-24.4701938629150,64.3233947753906,
-20.9680919647217,17.6398410797119,
-19.7980690002441,-24.1111621856689,
-10.4512062072754,-21.7773723602295,
13.1990880966187,13.4323663711548,
29.8915748596191,30.7612419128418,
15.8302345275879,0.410167932510376,
-14.5090808868408,-48.6324958801270,
-12.4699831008911,-64.3665008544922,
33.3382530212402,-36.8493995666504,
72.4312973022461,9.66281890869141,
60.0084075927734,41.1209411621094,
18.4026279449463,41.9318161010742,
12.3304138183594,20.5873699188232,
48.6194725036621,7.82301330566406,
66.7185974121094,23.9646434783936,
25.9241523742676,52.1016464233398,
-35.1791839599609,49.4257850646973,
-50.2853698730469,3.20453929901123,
-9.07894039154053,-41.8657531738281,
34.7073860168457,-37.0419540405273,
41.2913551330566,6.12221622467041,
22.0174598693848,25.0089511871338,
6.68843412399292,-10.2387981414795,
4.20109558105469,-54.6679344177246,
5.84672212600708,-57.0789375305176,
10.1555633544922,-22.9314689636230,
15.0616283416748,13.0205593109131,
9.08561801910400,34.8934288024902,
-11.4769535064697,48.9413223266602,
-16.1254291534424,52.2385902404785,
11.6415748596191,33.1554069519043,
47.8635444641113,7.87875890731812,
43.5955238342285,8.53110122680664,
-4.90952348709106,35.0433845520020,
-52.7458648681641,41.6607933044434,
-57.8256988525391,11.8894824981689,
-29.6564273834229,-13.9873142242432,
-5.00989341735840,6.03450012207031,
6.37415122985840,44.2441711425781,
12.5372905731201,44.1710929870606,
14.6465501785278,4.98890209197998,
10.2379245758057,-15.3819847106934,
15.3756132125855,7.12367105484009,
43.3551483154297,34.0608940124512,
70.7712173461914,25.8174209594727,
56.6386108398438,2.13569021224976,
-0.109302997589111,6.53420352935791,
-52.2366180419922,27.3856067657471,
-58.9637794494629,16.4720230102539,
-32.6448860168457,-34.2735671997070,
-11.7633047103882,-70.6797180175781,
-6.79547882080078,-54.3651733398438,
-1.31538009643555,-12.9562072753906,
5.09008502960205,4.22242879867554,
1.22014760971069,-14.0537109375000,
-5.72601985931397,-39.5818786621094,
1.83013713359833,-49.7429580688477,
18.2254810333252,-39.2713737487793,
15.0686235427856,-12.6982841491699,
-11.7011213302612,22.3697566986084,
-24.5946388244629,44.2681312561035,
3.46432971954346,35.0274276733398,
43.2998275756836,5.25400161743164,
51.1084671020508,-12.3281936645508,
25.4901084899902,-4.85856056213379,
12.8130159378052,4.87343454360962,
30.7258949279785,-2.72465801239014,
39.9090423583984,-8.22688198089600,
10.3992862701416,11.4349660873413,
-32.4906005859375,47.0302429199219,
-42.0142059326172,70.0768203735352,
-12.4130859375000,60.5695686340332,
15.4892597198486,27.5049400329590,
10.6310119628906,1.43405604362488,
-13.3079776763916,2.26826095581055,
-27.1153793334961,25.6407356262207,
-21.4331169128418,42.3606491088867,
-4.14400815963745,20.1914539337158,
19.9310455322266,-31.1343936920166,
42.4074249267578,-57.3941459655762,
44.4005889892578,-18.4855346679688,
23.7846164703369,44.8387985229492,
6.72966909408569,54.8104820251465,
11.6640110015869,4.52612638473511,
19.3489265441895,-33.3191757202148,
-2.16435265541077,-8.97132110595703,
-40.5264472961426,30.9721488952637,
-49.2636299133301,11.2086343765259,
-12.5175647735596,-53.6819648742676,
26.0186614990234,-72.6369476318359,
24.3601493835449,-9.06106758117676,
1.15300667285919,62.0562057495117,
0.333612650632858,62.0121269226074,
19.3753833770752,15.9781627655029,
17.1819038391113,-1.63848185539246,
-18.2542324066162,21.3426837921143,
-52.9046707153320,23.8788623809814,
-57.3575706481934,-21.5163955688477,
-46.5118942260742,-59.2040824890137,
-43.2684631347656,-40.9502334594727,
-43.8644447326660,1.61104953289032,
-30.0074539184570,6.63740301132202,
-5.13958787918091,-26.3194618225098,
9.67596149444580,-38.2570724487305,
3.10486412048340,-4.76149129867554,
-14.7634315490723,30.7413654327393,
-29.2820358276367,28.5778121948242,
-35.0654830932617,9.30241012573242,
-24.8705787658691,16.3925323486328,
2.80434226989746,38.6535797119141,
29.7268981933594,41.5136909484863,
36.9783096313477,12.9748353958130,
25.4436054229736,-13.6826763153076,
9.13778781890869,-17.2766075134277,
-6.58998489379883,-14.7188377380371,
-16.1911640167236,-22.4576396942139,
-15.7470264434814,-23.9772644042969,
-1.38918089866638,-1.20732104778290,
9.96913242340088,21.6457691192627,
0.708885610103607,13.0695266723633,
-19.9542980194092,-16.6001758575439,
-18.4813060760498,-25.0238113403320,
10.4642210006714,5.66628026962280,
27.1103992462158,46.1073684692383,
2.41828250885010,65.1965942382813,
-30.6462612152100,64.4655075073242,
-27.4665031433105,62.9538497924805,
0.0326757431030273,56.4950828552246,
-1.68127775192261,30.3021697998047,
-42.3252029418945,-2.53517842292786,
-74.4461364746094,-14.5758361816406,
-56.1581115722656,-5.53777599334717,
-11.0122756958008,-0.135857254266739,
10.7233886718750,-11.3385496139526,
4.12495040893555,-23.3918857574463,
-1.67897164821625,-24.1241168975830,
2.28958749771118,-19.6897125244141,
-1.05899000167847,-23.8252964019775,
-13.5310306549072,-33.7429428100586,
-6.12154102325439,-37.8320045471191,
27.0500698089600,-39.3471450805664,
50.1967544555664,-42.5428123474121,
35.0524902343750,-36.7412376403809,
8.53137397766113,-14.4908142089844,
10.3234968185425,6.09733200073242,
38.5709304809570,-0.659453868865967,
47.8054771423340,-20.6838207244873,
15.3732910156250,-20.4344882965088,
-31.3705520629883,1.07067751884460,
-44.9126319885254,4.28635311126709,
-18.4195518493652,-34.0203323364258,
22.0975131988525,-70.7785644531250,
50.2889442443848,-51.3471260070801,
49.5026664733887,12.7464914321899,
21.2735843658447,51.4855957031250,
-16.7288761138916,25.9878749847412,
-39.2416000366211,-26.1382713317871,
-34.5589714050293,-42.3928413391113,
-19.8854846954346,-15.1458330154419,
-18.9260540008545,16.8472976684570,
-29.6028137207031,26.2807140350342,
-35.1430549621582,23.8083305358887,
-28.9379291534424,24.4878120422363,
-26.5993976593018,19.9307365417480,
-36.0749931335449,-7.18711948394775,
-34.2164192199707,-48.3424263000488,
0.572943806648254,-61.9002304077148,
50.0738449096680,-27.7844543457031,
73.9126052856445,20.7598438262939,
55.3594970703125,30.8272857666016,
22.6503601074219,-7.96309757232666,
13.7648763656616,-51.9039802551270,
28.9174575805664,-48.0837364196777,
37.0182533264160,0.0634560585021973,
18.7394180297852,29.8083667755127,
-12.6274299621582,5.35555076599121,
-32.4322586059570,-36.3113632202148,
-31.7475852966309,-38.4092178344727,
-17.0381679534912,-3.78930020332336,
-0.305420458316803,9.05760002136231,
5.91848611831665,-27.1143760681152,
-2.07979655265808,-66.5585250854492,
-13.1461944580078,-48.4988479614258,
-9.06566143035889,12.0144100189209,
5.52492713928223,43.0465126037598,
8.44591140747070,18.8029098510742,
-9.64498519897461,-15.0222377777100,
-27.2680377960205,-16.7981796264648,
-12.2813529968262,-7.10920381546021,
20.8525295257568,-21.2587013244629,
28.7472171783447,-46.2757949829102,
-1.08292818069458,-41.8263282775879,
-29.4775371551514,-12.6113471984863,
-29.1789226531982,-2.56108713150024,
-13.1163196563721,-18.8605575561523,
-5.66723728179932,-17.6517562866211,
-3.92889070510864,22.3560390472412,
5.63553762435913,55.9553375244141,
7.79642009735107,39.6007347106934,
-18.2207145690918,-0.512427151203156,
-48.2163848876953,-6.21249008178711,
-35.7021141052246,18.6769485473633,
14.9824905395508,17.3194694519043,
44.1290397644043,-21.9605731964111,
21.9712066650391,-47.3301811218262,
-5.42851829528809,-22.4940528869629,
9.46697616577148,16.8065643310547,
36.8640022277832,18.9419670104980,
19.2071552276611,-10.5666484832764,
-36.0724983215332,-21.3947143554688,
-61.6667747497559,-2.40661430358887,
-28.7860298156738,5.05553388595581,
14.6443252563477,-18.5717391967773,
13.9512739181519,-44.8986053466797,
-17.5630779266357,-40.8706512451172,
-29.4482955932617,-11.7128858566284,
-10.5762958526611,20.6083106994629,
9.14078426361084,37.8451347351074,
12.7640285491943,34.2528114318848,
12.6600170135498,14.3591032028198,
11.9148836135864,-1.32721900939941,
-0.503426909446716,14.2145652770996,
-19.5973224639893,51.6893463134766,
-27.7109680175781,59.3865089416504,
-17.0919437408447,1.96378064155579,
0.588967978954315,-71.9664993286133,
14.6618499755859,-77.1566238403320,
24.1203937530518,-8.60005950927734,
26.7697830200195,49.0111007690430,
11.2510023117065,36.4486236572266,
-21.2640533447266,-7.39479351043701,
-36.9578475952148,-10.1892166137695,
-16.4564704895020,27.6998786926270,
9.30631637573242,43.0555915832520,
4.12665319442749,10.0926933288574,
-13.4750528335571,-28.9403095245361,
-3.95993661880493,-35.0773391723633,
29.4205493927002,-22.9464836120605,
36.8353996276856,-23.0098648071289,
2.55192565917969,-22.7941360473633,
-24.6510009765625,3.30283069610596,
-0.360507488250732,38.4270858764648,
46.0624961853027,40.0201492309570,
55.4020767211914,10.6483364105225,
27.4405803680420,-6.07736968994141,
15.1157922744751,10.1316699981689,
30.0600452423096,35.2620887756348,
31.2198657989502,30.4929294586182,
-4.15286636352539,-6.84834289550781,
-29.0927448272705,-47.5386734008789,
0.732904911041260,-64.3519515991211,
54.6866874694824,-49.4935684204102,
66.1922454833984,-8.89365196228027,
28.3120765686035,31.0381622314453,
-3.19652295112610,32.3381690979004,
8.85224914550781,-1.97675871849060,
35.6391105651856,-26.3774547576904,
36.4457664489746,-5.66487979888916,
23.9680175781250,36.2981262207031,
28.3588695526123,51.0677185058594,
39.0581398010254,34.8527145385742,
17.9826087951660,25.1907024383545,
-31.3443145751953,40.6786842346191,
-66.5869827270508,53.3182716369629,
-60.2499694824219,37.6602516174316,
-32.9349555969238,17.5395069122314,
-19.6610183715820,22.4651870727539,
-28.5750885009766,34.3532066345215,
-39.8894195556641,10.1754713058472,
-42.3814010620117,-41.0478248596191,
-37.0534896850586,-67.2918243408203,
-20.8092651367188,-41.2559165954590,
6.42347908020020,1.55282187461853,
29.6786994934082,19.3381023406982,
37.1307296752930,13.6812820434570,
36.4687957763672,6.78533029556274,
38.4211616516113,3.49615955352783,
41.3472328186035,-13.2205448150635,
35.2520408630371,-39.0847473144531,
27.5156326293945,-42.8521347045898,
33.1134223937988,-14.8711118698120,
42.9275398254395,23.0551528930664,
29.8445930480957,46.6317787170410,
-14.5735597610474,56.8896102905273,
-50.7641448974609,59.3151931762695,
-44.1114349365234,48.4290237426758,
-14.4468479156494,22.7735786437988,
-6.66322326660156,4.03623628616333,
-28.6217651367188,3.80400371551514,
-42.8181686401367,2.62444496154785,
-22.5446853637695,-27.5839710235596,
11.6968231201172,-73.5415725708008,
23.2744770050049,-84.9021072387695,
3.99785637855530,-43.8693733215332,
-23.7222976684570,5.18277311325073,
-40.3799133300781,6.03176307678223,
-38.3669815063477,-34.6224594116211,
-18.3372478485107,-57.1587524414063,
14.2914695739746,-29.7908878326416,
36.9223632812500,18.9687080383301,
26.6820030212402,35.9176712036133,
-14.6511383056641,9.31046390533447,
-48.1258010864258,-22.2183647155762,
-40.9502677917481,-23.0516262054443,
-4.23200321197510,3.59619688987732,
25.0704154968262,26.0996093750000,
21.3842144012451,24.7975120544434,
-6.47884178161621,9.12245655059815,
-25.7617969512939,6.84728288650513,
-22.1864051818848,24.8699283599854,
-7.03899002075195,44.2201461791992,
-0.608183324337006,32.4227485656738,
-6.61024761199951,-5.05286359786987,
-12.8901863098145,-32.0067329406738,
-8.30185031890869,-17.4901657104492,
-0.819311976432800,22.0915756225586,
-8.25306320190430,44.0393180847168,
-30.0175189971924,27.6306724548340,
-40.3328247070313,2.68029117584229,
-18.2309303283691,5.31074810028076,
18.7283916473389,25.6332817077637,
30.5311489105225,25.0158920288086,
5.93184137344360,-8.59547805786133,
-27.5174751281738,-45.8560752868652,
-38.2991943359375,-54.0233650207520,
-31.6365756988525,-42.0286521911621,
-32.9638481140137,-37.4082832336426,
-39.9665756225586,-48.8531074523926,
-25.5667724609375,-56.7982406616211,
16.4103660583496,-46.7939682006836,
51.6643943786621,-26.9276905059814,
46.4484481811523,-9.50886535644531,
12.9329757690430,4.29193115234375,
-8.88168430328369,14.2464609146118,
-2.25080299377441,13.3845443725586,
13.5666799545288,0.816654086112976,
18.5079383850098,-9.21184730529785,
14.8483161926270,-4.97494506835938,
8.93141365051270,5.49295473098755,
1.10262894630432,10.8233890533447,
-10.6956853866577,16.5982017517090,
-21.1092967987061,32.3791656494141,
-17.0567703247070,46.0412063598633,
-2.33756089210510,25.4037818908691,
9.97760391235352,-24.5268516540527,
17.1753559112549,-55.8821144104004,
20.6537189483643,-30.7017402648926,
19.5899467468262,20.6938114166260,
14.8956165313721,42.5050964355469,
11.4483184814453,19.0083904266357,
4.85451984405518,-6.08332109451294,
-8.98993492126465,0.608900964260101,
-23.0327568054199,25.0847892761230,
-15.3910150527954,34.4801635742188,
17.7729282379150,26.5355148315430,
40.7041664123535,23.0720176696777,
11.3604030609131,22.7890720367432,
-50.0550651550293,8.76915359497070,
-68.0789413452148,-16.7087917327881,
-5.71071243286133,-29.2514743804932,
78.0132293701172,-19.5214443206787,
94.5170516967773,-9.47442054748535,
39.8314895629883,-16.3235664367676,
-11.4061250686646,-33.0957870483398,
-5.89244747161865,-48.0085067749023,
27.8747825622559,-58.3541107177734,
32.9533805847168,-60.8336296081543,
1.34969711303711,-40.8620986938477,
-29.6864261627197,3.35164260864258,
-37.6656074523926,36.0977668762207,
-33.8279953002930,16.6390247344971,
-28.9546184539795,-37.6171531677246,
-17.6916389465332,-67.1282730102539,
0.238196134567261,-46.1193122863770,
13.0704250335693,-7.50704956054688,
20.2494487762451,7.41437387466431,
33.7053222656250,1.97495627403259,
51.0952758789063,4.12739562988281,
46.6364631652832,16.4727745056152,
12.5531558990479,17.6825866699219,
-25.8274173736572,2.69440793991089,
-31.7186546325684,-10.9866304397583,
-11.6054954528809,-13.0325431823730,
-5.68961954116821,-14.5038938522339,
-25.4175529479980,-16.5098114013672,
-40.1088714599609,-5.98330163955689,
-29.5545558929443,24.8290061950684,
-14.0922670364380,49.6949806213379,
-16.5628242492676,38.3822479248047,
-22.2864227294922,5.27666902542114,
1.06486105918884,-13.6752395629883,
45.7040023803711,0.0890755653381348,
66.1685638427734,31.9182071685791,
43.8659515380859,48.4408493041992,
14.6906433105469,33.5962066650391,
16.1032009124756,4.87511253356934,
31.3930988311768,-8.33312702178955,
17.3405475616455,3.03005790710449,
-23.9144191741943,18.1849632263184,
-46.7118415832520,4.58862972259522,
-28.7675933837891,-31.4020881652832,
4.68223190307617,-41.0666809082031,
20.5286273956299,5.28601646423340,
22.8809413909912,64.1148834228516,
26.9248542785645,61.2722549438477,
26.2522869110107,-4.23376750946045,
3.17111539840698,-54.7804603576660,
-27.2797832489014,-37.5704956054688,
-31.7655105590820,5.56499242782593,
-10.9442920684814,4.90926408767700,
0.946179151535034,-37.6089324951172,
-11.7261409759521,-51.6314201354981,
-18.3338127136230,-8.36942291259766,
0.215623617172241,41.7026786804199,
20.0227260589600,49.0826110839844,
10.7608823776245,32.1870155334473,
-17.0367279052734,29.3998451232910,
-31.4996986389160,30.0762367248535,
-22.4503421783447,5.00489521026611,
-13.3186607360840,-29.7713661193848,
-18.4575595855713,-23.0629787445068,
-20.9154052734375,29.2927227020264,
-12.7313156127930,69.5471420288086,
-5.62691116333008,62.4463233947754,
-11.9123573303223,37.3259658813477,
-20.6024093627930,37.9304466247559,
-25.7650032043457,55.9551277160645,
-30.1602287292480,49.8136253356934,
-31.4872074127197,19.6116924285889,
-21.1800251007080,6.35795259475708,
-4.19756221771240,19.7282047271729,
-7.45534706115723,19.0997791290283,
-37.7488059997559,-14.8968877792358,
-54.3720245361328,-49.8368797302246,
-17.4968547821045,-43.0181007385254,
50.8706092834473,-5.79526567459106,
84.2620544433594,19.7413482666016,
61.1836700439453,16.5563068389893,
28.8881206512451,9.96578025817871,
26.4315891265869,20.4674682617188,
26.6684722900391,34.6045761108398,
-10.7166070938110,31.9161529541016,
-67.5133590698242,19.5913505554199,
-81.4034118652344,6.46489381790161,
-33.0898628234863,-5.72095727920532,
26.7895622253418,-17.7149467468262,
41.0819015502930,-17.7269020080566,
10.6663169860840,-3.94650864601135,
-22.6313304901123,11.7311334609985,
-34.5155601501465,16.1092872619629,
-29.0288791656494,16.8122673034668,
-13.2796411514282,25.5449581146240,
9.09546661376953,38.0197296142578,
24.5223941802979,35.6077156066895,
16.7520847320557,13.2616367340088,
-1.90503668785095,-9.44539165496826,
-7.41245698928833,-25.3732204437256,
7.41082906723023,-44.5763511657715,
21.5534744262695,-63.5622825622559,
19.6957817077637,-60.0510063171387,
8.66319847106934,-30.3930664062500,
2.98599600791931,-2.02258372306824,
-5.81389856338501,-3.37241649627686,
-30.9084568023682,-24.1908111572266,
-51.4504280090332,-36.3451004028320,
-37.6406211853027,-36.6552848815918,
4.93643569946289,-37.7067985534668,
38.7588729858398,-32.5667839050293,
41.3770637512207,6.57138156890869,
27.5591545104980,67.0577850341797,
14.1410217285156,91.7141952514648,
-2.14085602760315,43.4530601501465,
-21.2999153137207,-30.3750972747803,
-20.1973953247070,-57.2124443054199,
13.0918025970459,-23.3234558105469,
43.6816177368164,18.2940502166748,
24.6968708038330,21.9087429046631,
-34.5479888916016,1.06313252449036,
-69.0680389404297,-11.5947637557983,
-40.0973854064941,-7.50102138519287,
15.8350830078125,-2.38960266113281,
39.8586311340332,3.75012564659119,
24.3600692749023,19.1248550415039,
5.21185159683228,38.4150619506836,
5.37944555282593,43.4000740051270,
9.28403377532959,34.4095268249512,
-3.85882520675659,34.1951828002930,
-23.1739616394043,49.0531616210938,
-29.3172149658203,56.4351501464844,
-17.4639930725098,40.0970687866211,
-0.137881249189377,12.4166297912598,
14.2584571838379,0.714099287986755,
28.5265750885010,9.99452400207520,
43.0889320373535,18.8268184661865,
51.0035247802734,13.0949039459229,
48.0289154052734,6.05642938613892,
34.3933677673340,16.3388347625732,
7.75335407257080,37.2734642028809,
-24.5783348083496,46.2650985717773,
-52.4458236694336,30.9675216674805,
-61.9903640747070,1.85451579093933,
-41.0541305541992,-22.1290473937988,
-0.489515781402588,-30.8486557006836,
34.7744483947754,-31.9763889312744,
42.8131065368652,-31.7381362915039,
25.3692340850830,-24.0665721893311,
2.16026353836060,0.672872900962830,
-6.40281724929810,33.0363655090332,
1.36998140811920,47.8368377685547,
4.98937606811523,25.0759029388428,
-7.47379589080811,-22.0005455017090,
-16.4860420227051,-51.1756401062012,
5.42086124420166,-35.8169746398926,
47.5723915100098,0.867075562477112,
66.0998229980469,13.9397525787354,
28.5509071350098,-2.43649244308472,
-32.6448936462402,-12.6732225418091,
-60.9468917846680,3.16644692420959,
-42.9221534729004,22.8638477325439,
-20.8906269073486,11.1569042205811,
-27.0132751464844,-22.5520935058594,
-31.1408061981201,-34.6928939819336,
5.80604648590088,-13.9403963088989,
57.7003326416016,0.107863426208496,
59.1959915161133,-13.9458189010620,
0.516800880432129,-26.8688488006592,
-50.9477310180664,-12.8762884140015,
-35.4553718566895,8.93056392669678,
26.5983390808105,6.34601449966431,
63.5227622985840,-3.75486183166504,
42.7999076843262,17.9454574584961,
-4.82264137268066,56.6936912536621,
-42.5132980346680,47.3335990905762,
-54.4981613159180,-18.9632644653320,
-41.8987770080566,-62.7655601501465,
-13.5745754241943,-22.8988513946533,
3.08395671844482,49.1779403686523,
-16.1137695312500,54.1203193664551,
-51.4063606262207,-11.1677436828613,
-50.3708343505859,-49.8809204101563,
-6.11498069763184,-11.8616380691528,
23.5800514221191,44.7975807189941,
-4.93516921997070,41.5273857116699,
-55.5341835021973,-2.59841132164001,
-54.3312377929688,-16.2522926330566,
0.310732364654541,12.9914722442627,
31.0638198852539,25.7738552093506,
-5.12938928604126,-17.6304512023926,
-53.2725372314453,-74.5538711547852,
-46.8677024841309,-80.2560729980469,
3.17716789245605,-31.2233619689941,
30.3450393676758,20.8784885406494,
3.01523876190186,40.6497688293457,
-39.9689483642578,28.7506217956543,
-55.0104331970215,0.934393644332886,
-42.7847709655762,-27.6870498657227,
-23.4256610870361,-54.1168594360352,
-5.23594474792481,-75.8018035888672,
15.4137859344482,-76.7876892089844,
25.0496025085449,-43.7933540344238,
17.5856742858887,14.9387207031250,
12.2536077499390,60.6850204467773,
24.9169311523438,55.2419700622559,
36.0124320983887,8.48818016052246,
18.5226860046387,-26.0885105133057,
-14.2499103546143,-15.3259572982788,
-19.0095043182373,9.86544799804688,
13.4268817901611,-3.08360528945923,
38.3023452758789,-39.7730674743652,
16.6834087371826,-44.7034530639648,
-25.2284946441650,2.96072149276733,
-37.1506538391113,56.4828834533691,
-19.4386024475098,61.2737274169922,
-20.6225070953369,20.9045581817627,
-54.0401992797852,-22.4279556274414,
-69.2693405151367,-40.5760574340820,
-26.2745628356934,-40.2374343872070,
38.3398590087891,-23.7839050292969,
57.9829597473145,5.17764568328857,
19.8513965606689,21.5134544372559,
-20.1626243591309,1.57150065898895,
-16.3231563568115,-40.9637870788574,
13.7540998458862,-50.0206604003906,
19.3087272644043,-1.71144485473633,
-7.21350383758545,52.6097373962402,
-26.3498134613037,52.4890480041504,
-8.24948120117188,5.43154239654541,
30.0575466156006,-23.3249950408936,
50.2331237792969,-1.76425838470459,
29.3800735473633,31.0059261322022,
-8.78194713592529,22.0937232971191,
-19.7903003692627,-20.9786224365234,
6.76186656951904,-42.9347648620606,
36.0539588928223,-17.8549480438232,
33.7326698303223,30.0130691528320,
6.18949365615845,59.2665214538574,
-6.50736522674561,54.1093597412109,
18.8224220275879,21.9080238342285,
47.4308891296387,-18.0744934082031,
37.5173034667969,-37.2673454284668,
3.80191946029663,-16.1377696990967,
-10.1778364181519,27.0389328002930,
0.306623816490173,50.5857048034668,
-8.51383399963379,31.5994052886963,
-51.0212211608887,-5.91471004486084,
-77.7309494018555,-15.9346628189087,
-40.7736396789551,5.19664955139160,
28.4566802978516,22.2994537353516,
49.2566680908203,17.2175426483154,
7.64105796813965,1.95102679729462,
-28.4677085876465,-9.11437606811523,
-3.73880958557129,-13.7140083312988,
45.9808807373047,-12.6288290023804,
49.2490653991699,-1.77262628078461,
-1.69870090484619,10.8979225158691,
-52.3948173522949,6.47190427780151,
-65.2256698608398,-14.2094774246216,
-54.2719001770020,-21.2624492645264,
-36.7069511413574,0.138423204421997,
-12.6946296691895,17.6009120941162,
16.0762615203857,-6.92147064208984,
28.0193328857422,-48.3947143554688,
9.25299739837647,-44.4084739685059,
-19.5425090789795,12.3093013763428,
-30.4001979827881,60.0851707458496,
-27.8174800872803,51.3492927551270,
-33.1716957092285,13.3401546478271,
-41.4628105163574,-6.48438119888306,
-29.2653770446777,-13.3338670730591,
-5.89813661575317,-38.6983337402344,
3.27991867065430,-68.3618698120117,
-0.979478120803833,-56.4679374694824,
7.06342935562134,-3.05350255966187,
34.7719078063965,27.1768417358398,
47.3092041015625,-0.628230810165405,
18.8750476837158,-34.9322395324707,
-19.8995151519775,-8.64306735992432,
-28.6640167236328,59.8643569946289,
-14.3622455596924,89.3198623657227,
-20.3340930938721,44.9283828735352,
-49.6548309326172,-22.4510974884033,
-58.9871253967285,-47.1725959777832,
-30.6627292633057,-17.7197189331055,
-4.00623178482056,22.0871334075928,
-17.5160789489746,34.1437568664551,
-50.5221862792969,16.6895141601563,
-51.1117172241211,-14.5459976196289,
-6.33036613464356,-39.9356117248535,
42.1704101562500,-46.6902236938477,
54.9087257385254,-32.9884529113770,
34.5404090881348,-15.7907409667969,
7.14922380447388,-5.02461957931519,
-5.12424278259277,8.37639331817627,
1.14753782749176,27.1165599822998,
24.9208354949951,35.6567649841309,
53.0905189514160,21.5557174682617,
59.2946243286133,0.426632463932037,
32.3413887023926,1.72384369373322,
-5.70708179473877,32.0679359436035,
-26.0438518524170,53.1636543273926,
-19.5152416229248,35.8430976867676,
1.12952530384064,2.43495941162109,
11.0407714843750,-9.13446331024170,
0.314927339553833,-1.53840041160584,
-16.7264900207520,-2.74284124374390,
-15.0778760910034,-15.1773424148560,
16.3782005310059,-7.50020837783814,
54.9253883361816,29.2508068084717,
55.6641082763672,53.2440795898438,
9.11577606201172,27.1062793731689,
-35.3716735839844,-17.4592552185059,
-25.4775238037109,-19.4052639007568,
18.4116516113281,23.4280223846436,
24.8255233764648,52.1936798095703,
-29.2154655456543,30.9827346801758,
-78.0972290039063,-3.03943324089050,
-57.5801467895508,-5.75657463073731,
9.88579082489014,2.23856043815613,
48.5207214355469,-22.5087718963623,
29.8752136230469,-64.2426681518555,
3.07508969306946,-61.5609016418457,
6.98697662353516,1.09356784820557,
16.2105579376221,59.4227828979492,
-2.32548785209656,53.2531394958496,
-28.2234172821045,0.172229766845703,
-20.7802085876465,-32.8081054687500,
12.2243509292603,-19.4191551208496,
21.8548545837402,8.86285018920898,
-6.14743757247925,22.5131206512451,
-29.3757514953613,26.1848411560059,
-17.8815498352051,32.0617980957031,
6.74762058258057,37.9111557006836,
11.2817516326904,38.3739089965820,
4.47424840927124,33.7476158142090,
15.9995145797730,29.4654560089111,
41.4115447998047,27.4848003387451,
41.0053863525391,21.6648311614990,
7.33445215225220,6.29229068756104,
-18.8362445831299,-16.9931259155273,
-11.8080854415894,-41.8807754516602,
5.75359392166138,-52.2987937927246,
-0.355574905872345,-35.8156356811523,
-28.7199382781982,-13.6219606399536,
-47.2351570129395,-14.7829141616821,
-39.9333839416504,-30.2491569519043,
-22.6235370635986,-18.7018241882324,
-8.18877410888672,28.4306278228760,
6.26830625534058,66.0626754760742,
17.7691230773926,53.1292190551758,
11.1026220321655,16.0622043609619,
-9.42208576202393,12.1672029495239,
-16.9500656127930,43.7371559143066,
-0.543809533119202,47.3205451965332,
10.5134325027466,-4.00032043457031,
-7.32073450088501,-56.9607276916504,
-29.8604946136475,-47.7090835571289,
-15.0615978240967,6.59731912612915,
31.1157665252686,34.0362358093262,
53.4487304687500,13.3091535568237,
18.7674465179443,-2.87939381599426,
-34.2099952697754,21.9431762695313,
-45.1524696350098,53.7209625244141,
-15.5186958312988,40.0468597412109,
8.73350334167481,-11.9639606475830,
-2.63972949981689,-48.2126541137695,
-31.3682842254639,-36.0474205017090,
-44.9624786376953,-3.38895034790039,
-29.0538558959961,2.66053104400635,
4.66734647750855,-22.3045845031738,
37.1616821289063,-45.1237678527832,
50.2940254211426,-35.9114265441895,
37.0467224121094,3.27023601531982,
16.5405464172363,44.2077941894531,
17.2642250061035,50.7579078674316,
36.2239952087402,20.2786827087402,
32.8891830444336,-7.57963609695435,
-11.9876604080200,-1.71121788024902,
-54.0403480529785,20.5331363677979,
-45.7989349365234,12.6469154357910,
-6.34505176544189,-32.4929656982422,
3.87283015251160,-67.9287948608398,
-31.4965629577637,-49.4466361999512,
-52.1416664123535,1.22630095481873,
-13.1090803146362,30.0098400115967,
45.0629806518555,25.6841831207275,
48.3091125488281,22.7437095642090,
-2.69080185890198,32.7071113586426,
-39.2369194030762,24.1465454101563,
-25.6184520721436,-15.6137571334839,
-1.19961369037628,-51.5522842407227,
-7.37613105773926,-44.8688316345215,
-21.8971462249756,-9.24026489257813,
-5.85466861724854,13.9374666213989,
28.0504760742188,14.1506900787354,
33.4921836853027,12.4733390808105,
-1.87185347080231,15.6935644149780,
-42.2654190063477,10.0767335891724,
-50.8155632019043,1.28101181983948,
-36.5179138183594,16.0084590911865,
-19.9240798950195,54.5060920715332,
-2.90288400650024,69.1736526489258,
13.9976835250855,38.7910118103027,
17.1416759490967,5.21242284774780,
6.44222068786621,10.9500761032105,
6.16469621658325,36.9927520751953,
23.3730888366699,31.2557945251465,
30.3685207366943,-6.08775234222412,
11.0690679550171,-20.0447750091553,
-8.80406951904297,13.3065223693848,
4.85306358337402,49.0051383972168,
31.8836765289307,37.1667976379395,
19.4273719787598,-1.37214815616608,
-35.8896865844727,-15.8124294281006,
-67.3649520874023,-6.46885204315186,
-30.4748516082764,-10.2226667404175,
31.0162582397461,-30.4547672271729,
50.5299987792969,-30.8675212860107,
21.3382186889648,2.62893271446228,
-7.99691390991211,34.4681320190430,
-12.4433431625366,34.1037864685059,
-6.23915147781372,15.6809873580933,
-0.537507832050324,14.1476383209229,
13.0490350723267,24.3705959320068,
32.2131462097168,21.3820018768311,
34.5627899169922,9.70101928710938,
14.5641832351685,12.3948020935059,
-3.24875879287720,20.1722450256348,
3.09063076972961,-2.93247509002686,
13.0875139236450,-49.2963867187500,
2.69696569442749,-59.8838386535645,
-15.1771011352539,-16.7361335754395,
-14.0143108367920,24.9592151641846,
-4.36876678466797,7.12928342819214,
-10.2865142822266,-39.0525894165039,
-24.9067668914795,-34.8710441589356,
-29.3465499877930,27.1342010498047,
-24.7905292510986,65.6153869628906,
-32.1953353881836,25.4397983551025,
-47.9577178955078,-39.7825202941895,
-38.4723434448242,-51.1157493591309,
-2.35104274749756,-3.89851665496826,
13.3033008575439,41.4614562988281,
-20.1937713623047,45.9431266784668,
-64.0119171142578,24.5238208770752,
-60.8136978149414,-2.55254411697388,
-21.4244346618652,-34.6688079833984,
-3.58060359954834,-62.0741462707520,
-16.7133426666260,-59.4138526916504,
-12.6253747940063,-18.7442722320557,
31.5211811065674,21.6734313964844,
69.8957901000977,28.2921237945557,
50.2210960388184,18.7006893157959,
-8.67797470092773,28.1116027832031,
-40.9667587280273,47.4122352600098,
-13.5753936767578,39.9217300415039,
36.4085502624512,6.52613353729248,
59.0610618591309,-14.2121162414551,
39.3950653076172,5.71726703643799,
2.47920584678650,41.0180664062500,
-22.4978008270264,50.2128143310547,
-20.7665386199951,30.9612674713135,
4.48431968688965,13.1838655471802,
27.7551326751709,4.37188911437988,
24.8809299468994,-6.83171129226685,
6.09444570541382,-21.7603015899658,
-5.63848352432251,-22.8586750030518,
-2.48637700080872,-8.41134643554688,
-1.12974834442139,-0.355186402797699,
-13.7410802841187,-4.26558780670166,
-33.2496719360352,1.38494515419006,
-39.8787498474121,34.8211784362793,
-33.1386299133301,70.9415512084961,
-25.2278099060059,72.5423355102539,
-16.0351505279541,33.6713943481445,
-2.23145294189453,-6.53912448883057,
-1.65273678302765,-20.3569431304932,
-29.0809288024902,-20.4514865875244,
-60.9654159545898,-26.9455471038818,
-51.9317092895508,-34.1341743469238,
6.99442291259766,-25.4141159057617,
62.1135444641113,0.556589484214783,
60.7672882080078,27.1719284057617,
21.1835250854492,43.5113220214844,
2.74041128158569,44.0969924926758,
21.3969306945801,32.2394180297852,
32.5602035522461,20.2177562713623,
11.5656738281250,23.5665206909180,
-8.65332031250000,43.1338958740234,
5.13829898834229,57.8354873657227,
20.9782600402832,43.6209640502930,
-7.18495559692383,5.87092161178589,
-58.0185012817383,-18.1593723297119,
-58.6020240783691,-14.5671195983887,
10.1726989746094,3.49359655380249,
70.4348449707031,18.5157546997070,
50.7798767089844,26.7261257171631,
-12.8249549865723,19.1116161346436,
-36.4684028625488,-13.2383651733398,
-4.67442035675049,-48.8232765197754,
18.9094562530518,-46.3918952941895,
-4.26062345504761,-1.49627733230591,
-38.1450424194336,32.2926712036133,
-37.5717277526856,7.68532943725586,
-14.1613311767578,-46.4777336120606,
-2.32165098190308,-51.8863677978516,
-2.37593102455139,3.18857860565186,
1.13864219188690,53.0501670837402,
-5.57205152511597,45.5130653381348,
-45.1677360534668,6.47660827636719,
-90.5131912231445,-18.3238582611084,
-79.7581329345703,-31.8897018432617,
-9.36954879760742,-52.4331588745117,
40.6617355346680,-61.8541336059570,
18.8081092834473,-33.4847908020020,
-29.7247657775879,5.54711580276489,
-38.1861228942871,-3.90205097198486,
-5.28435850143433,-56.0283889770508,
16.4852733612061,-72.5447006225586,
4.42478704452515,-10.3857040405273,
-14.5763502120972,71.7529602050781,
-20.0044555664063,85.5596694946289,
-25.7643108367920,32.7367744445801,
-28.7054386138916,-20.3973331451416,
-3.57633829116821,-42.1746368408203,
43.7623939514160,-45.1170997619629,
59.2543067932129,-35.5805206298828,
21.8420124053955,-5.04844236373901,
-13.6336994171143,36.0523376464844,
8.75516891479492,45.2888374328613,
51.6545829772949,10.7862043380737,
43.6703338623047,-21.2679901123047,
-18.0328998565674,-16.4401073455811,
-57.3961143493652,-0.400392293930054,
-31.7769527435303,-9.79914379119873,
13.0563087463379,-20.0867080688477,
12.5627079010010,15.2130908966064,
-20.4330940246582,69.5707855224609,
-36.3858299255371,64.7261962890625,
-30.5647926330566,-7.99960422515869,
-28.8081970214844,-66.6279067993164,
-32.2389259338379,-41.0185012817383,
-20.7301406860352,36.6450691223145,
-2.42807722091675,79.5894470214844,
-8.28680992126465,60.3403053283691,
-31.9624919891357,22.4293193817139,
-29.9215011596680,6.82741212844849,
10.8752431869507,4.06741428375244,
47.7375297546387,-3.75741481781006,
45.2364082336426,-11.4999361038208,
28.5060253143311,-12.2699146270752,
43.5031089782715,-12.9138936996460,
68.2215194702148,-9.43789386749268,
45.4882316589356,10.9404916763306,
-16.4471549987793,34.7484054565430,
-49.5289077758789,25.2992610931397,
-20.3868694305420,-17.7103786468506,
27.3687705993652,-45.7620162963867,
35.0917091369629,-21.5919322967529,
3.67407894134522,23.1388874053955,
-28.7420024871826,17.9313564300537,
-41.2070503234863,-37.8980865478516,
-39.8133354187012,-67.6214599609375,
-22.3231868743897,-30.1221179962158,
10.6814050674438,31.6412506103516,
26.2910175323486,55.1026191711426,
-9.89236164093018,39.7239532470703,
-70.9382629394531,21.3804454803467,
-79.9073181152344,11.2061548233032,
-16.5081939697266,-7.73948669433594,
50.3694076538086,-27.6072692871094,
53.4879455566406,-20.6966953277588,
11.2225351333618,7.34897613525391,
-13.5590000152588,9.81414794921875,
-2.49864935874939,-31.4605255126953,
4.89863204956055,-68.5406494140625,
-17.5301513671875,-50.7003746032715,
-37.0422096252441,-0.716581106185913,
-21.3444042205811,23.1584091186523,
13.4662075042725,6.90504550933838,
29.5328750610352,-11.1890220642090,
14.6030244827271,-11.9823837280273,
-12.8918313980103,-14.6219396591187,
-34.4414443969727,-35.7814331054688,
-35.8795242309570,-55.6697425842285,
-9.06122016906738,-47.8970451354981,
34.7155380249023,-29.5504779815674,
59.3552246093750,-30.0477924346924,
45.4702835083008,-41.4139595031738,
16.7477092742920,-32.7470397949219,
12.4971971511841,-1.96227240562439,
35.9284553527832,12.0532865524292,
51.3335151672363,-9.55268859863281,
37.1414489746094,-38.6779823303223,
16.4139080047607,-42.3343009948731,
14.9528865814209,-23.3345966339111,
18.9723110198975,-11.1038980484009,
3.14719843864441,-12.6394720077515,
-23.7679004669189,-12.1984958648682,
-32.7309799194336,-2.14865565299988,
-11.7001342773438,1.35627222061157,
14.4845657348633,-12.6365642547607,
18.8191375732422,-23.8807334899902,
-0.252802640199661,-10.2838010787964,
-20.4735107421875,19.6418895721436,
-23.3644332885742,38.7858772277832,
-3.21730113029480,34.0010604858398,
28.9271469116211,20.3559818267822,
50.2870063781738,15.9859199523926,
40.6109733581543,22.4634571075439,
7.17028379440308,19.0971088409424,
-13.2043371200562,-8.77510547637940,
4.93583059310913,-49.4584159851074,
45.6380348205566,-72.2682037353516,
65.0263214111328,-46.6917228698731,
43.5934638977051,18.9542884826660,
0.847926616668701,76.6161804199219,
-34.0259017944336,80.8204879760742,
-54.4611358642578,32.8401489257813,
-70.4352264404297,-22.6171379089355,
-77.7140579223633,-42.8348197937012,
-59.5401191711426,-30.0208396911621,
-14.0741300582886,-12.8745326995850,
28.0900859832764,-6.03712797164917,
33.3145141601563,2.69193840026855,
3.23333311080933,23.0009956359863,
-25.6685924530029,41.0178833007813,
-22.7589664459229,28.8712921142578,
3.75578069686890,-14.4018735885620,
23.9387626647949,-47.5974884033203,
22.8192329406738,-33.4085388183594,
13.9191551208496,16.5040626525879,
14.6046409606934,44.5438919067383,
15.3993291854858,20.0859909057617,
5.49194908142090,-26.5851688385010,
-9.18325614929199,-38.2601852416992,
-9.14883899688721,-2.77166986465454,
13.5510292053223,24.6636447906494,
35.7862014770508,8.37199401855469,
33.7790031433106,-17.7331752777100,
5.83372688293457,0.0920584201812744,
-26.4001922607422,54.3187675476074,
-44.3535232543945,73.5734329223633,
-47.1575698852539,21.1011409759522,
-41.4089202880859,-50.1062316894531,
-30.6726245880127,-60.6505661010742,
-11.0306930541992,-14.4354629516602,
18.3705387115479,11.4910936355591,
41.8038406372070,-20.8408050537109,
39.4888381958008,-62.1912956237793,
10.1031293869019,-46.6502037048340,
-19.4962234497070,13.6702213287354,
-22.6932525634766,42.3442306518555,
-3.95932865142822,4.14208936691284,
5.73354387283325,-45.0187225341797,
-9.89914894104004,-42.0244178771973,
-33.5840148925781,1.70639348030090,
-38.8214759826660,24.8856716156006,
-24.7603549957275,8.96490478515625,
-6.19228219985962,-4.02938985824585,
6.74727821350098,16.2014369964600,
17.0660190582275,41.9941596984863,
23.5643291473389,28.2240619659424,
19.0852966308594,-11.2078742980957,
6.30117416381836,-28.2337570190430,
-3.82095289230347,-8.33459854125977,
-5.37929487228394,7.21309232711792,
-2.57810473442078,-11.6474742889404,
5.36365222930908,-41.6533966064453,
17.0714759826660,-43.2751007080078,
25.3233547210693,-17.3547191619873,
21.6238098144531,9.77914333343506,
9.30267238616943,30.1482753753662,
2.09021973609924,48.2438926696777,
0.275179058313370,52.0447120666504,
-10.0751705169678,22.1915645599365,
-29.7540969848633,-22.9902172088623,
-28.5218753814697,-40.2955665588379,
6.93310737609863,-17.8538894653320,
45.1659545898438,-0.910316050052643,
42.4559288024902,-21.3487243652344,
8.80367469787598,-49.2830314636231,
-9.41749668121338,-32.5260963439941,
11.0372238159180,18.4339542388916,
37.8058128356934,38.9719963073731,
33.9393615722656,6.53942108154297,
5.52455949783325,-27.9657516479492,
-14.9031467437744,-11.5529985427856,
-17.2699470520020,39.5501556396484,
-16.3952751159668,59.9491767883301,
-15.5523900985718,21.4574699401855,
-0.632084965705872,-33.8876342773438,
24.6577796936035,-55.0647659301758,
36.2354354858398,-39.0618782043457,
26.6260967254639,-26.4252414703369,
17.1962146759033,-41.9649925231934,
33.1451110839844,-66.3841171264648,
58.3448410034180,-61.7972679138184,
61.5542984008789,-14.8860359191895,
40.3118705749512,42.9906997680664,
22.8717937469482,63.5722503662109,
21.3700809478760,36.2988624572754,
16.7955226898193,-0.00104880332946777,
-10.1671733856201,-5.95377635955811,
-40.8136825561523,18.9638729095459,
-42.6244773864746,40.5578269958496,
-23.2355327606201,33.4570236206055,
-16.5868301391602,11.2613506317139,
-30.9780941009522,1.37954545021057,
-31.1651592254639,7.27768278121948,
11.5470256805420,10.6459398269653,
67.8406066894531,6.28688812255859,
81.1359481811523,0.0831406116485596,
31.3188133239746,-3.59216928482056,
-29.0657329559326,-7.98247337341309,
-37.2725524902344,-9.22843360900879,
10.5815477371216,1.90420889854431,
57.6858787536621,25.0123805999756,
47.2541770935059,38.9737663269043,
-14.7190494537354,26.6603603363037,
-71.8562545776367,-3.47871875762939,
-73.3346328735352,-25.1248760223389,
-27.5573482513428,-31.9194297790527,
12.6736965179443,-32.7062492370606,
17.2723484039307,-26.7170333862305,
-2.43095612525940,2.60016202926636,
-20.9017429351807,46.8068199157715,
-33.2091674804688,64.4544219970703,
-47.3738822937012,30.6171264648438,
-57.7908782958984,-21.3030509948730,
-44.8944778442383,-34.7690696716309,
-10.5242624282837,-6.75185441970825,
9.93673229217529,11.2245702743530,
4.87193727493286,-13.5814275741577,
1.43909704685211,-45.7305259704590,
23.0811386108398,-32.3227462768555,
46.9699020385742,21.4495277404785,
28.3985157012939,59.2585525512695,
-23.6415901184082,49.5524520874023,
-47.9894752502441,17.4888248443604,
-15.0699062347412,-2.70463275909424,
34.1837081909180,-3.03159093856812,
39.8198966979981,0.666869163513184,
8.28770256042481,1.39321351051331,
-5.81742858886719,2.64413356781006,
15.9261856079102,10.1888494491577,
31.6487255096436,24.7928524017334,
7.78177547454834,38.4494438171387,
-30.8074131011963,40.9195899963379,
-38.1375579833984,24.1859474182129,
-15.5413751602173,-4.65076446533203,
5.46925115585327,-18.1021862030029,
15.0740442276001,-9.03417396545410,
26.8873195648193,-6.18160867691040,
40.4686126708984,-28.2676239013672,
29.4123077392578,-50.2948799133301,
-16.3675975799561,-42.1616020202637,
-57.8541755676270,-13.4120721817017,
-57.4448318481445,-7.40324592590332,
-30.9067420959473,-32.6273078918457,
-19.2186203002930,-49.7681274414063,
-33.6958618164063,-32.8295974731445,
-50.0427246093750,-8.72114944458008,
-47.1255455017090,-12.5739631652832,
-27.1814861297607,-23.1800498962402,
-1.51179254055023,1.96516954898834,
17.2075309753418,48.2780570983887,
12.7579517364502,61.8097381591797,
-20.6434593200684,24.7004585266113,
-57.8267478942871,-12.2129793167114,
-51.3101081848145,-4.29062128067017,
6.57434415817261,26.6227722167969,
61.5452423095703,33.8046646118164,
58.5058250427246,18.3865203857422,
8.32903099060059,10.0990762710571,
-36.9221572875977,15.0570087432861,
-53.0757522583008,2.62991714477539,
-54.3563919067383,-31.4729938507080,
-54.4060859680176,-43.9928703308106,
-44.5622291564941,-8.29430389404297,
-21.4221973419189,32.5529708862305,
-0.420538067817688,24.3060111999512,
1.76595497131348,-27.8737239837647,
3.06578779220581,-63.1549377441406,
16.4101543426514,-44.1844100952148,
24.6442604064941,6.31736755371094,
7.33249187469482,38.8757057189941,
-22.0350341796875,26.2101974487305,
-28.4487342834473,-14.4477443695068,
-7.38061618804932,-53.0140304565430,
9.60783767700195,-59.9759559631348,
10.9622964859009,-24.1003170013428,
15.3091764450073,23.9468898773193,
33.0232734680176,36.6044387817383,
39.8976287841797,2.05930638313293,
11.2260246276855,-38.5160522460938,
-27.2118473052979,-38.5733032226563,
-25.2771301269531,-6.30286121368408,
25.0147972106934,15.7353792190552,
70.1388778686523,13.5190343856812,
61.2391166687012,11.8335371017456,
9.34970474243164,24.2458362579346,
-32.3873252868652,20.9733085632324,
-29.0234794616699,-23.3369865417480,
7.35485553741455,-73.6932449340820,
40.5568351745606,-69.6832122802734,
40.4017066955566,-9.72196006774902,
7.82244968414307,43.1306610107422,
-24.5235900878906,33.4606323242188,
-26.3953742980957,-19.6222648620605,
5.41246986389160,-51.5675621032715,
38.5128822326660,-30.5654659271240,
41.0543022155762,21.1023464202881,
7.73441457748413,59.4359016418457,
-32.3810119628906,66.0442733764648,
-47.8062324523926,48.3281707763672,
-32.9094047546387,19.8494625091553,
-1.04310822486877,-6.47606706619263,
20.2887153625488,-20.2555313110352,
13.0538291931152,-21.7906246185303,
-10.8034114837646,-22.7994747161865,
-20.8684864044189,-32.8185043334961,
2.11818647384644,-37.9942741394043,
42.2748184204102,-20.4796123504639,
61.0547676086426,16.7672443389893,
48.7029800415039,46.2480468750000,
30.0520668029785,45.2661399841309,
32.6420173645020,29.2281208038330,
44.9175224304199,29.3454856872559,
30.0744800567627,49.3980827331543,
-23.0561218261719,56.2319831848145,
-75.8644638061523,26.6385517120361,
-77.8243560791016,-20.7754039764404,
-26.3035964965820,-42.6663780212402,
34.8812026977539,-27.1786403656006,
53.1480216979981,-2.14272403717041,
23.2711791992188,-2.55444502830505,
-16.6893653869629,-20.2716751098633,
-28.7678375244141,-19.2628459930420,
-7.43316078186035,11.4638538360596,
26.0063056945801,39.1493148803711,
49.8573341369629,30.7892055511475,
55.2347488403320,3.18221759796143,
42.3651084899902,2.17133712768555,
21.0642642974854,43.3615379333496,
-6.53107547760010,78.3253784179688,
-37.8967361450195,57.9304428100586,
-67.1301879882813,-3.07460355758667,
-76.8775711059570,-37.7320556640625,
-52.8290290832520,-25.1493167877197,
-10.4236297607422,-6.07859945297241,
18.3499126434326,-22.4751949310303,
12.8811635971069,-54.5248413085938,
-0.809471964836121,-54.7128410339356,
5.73056983947754,-23.8590812683105,
16.6230087280273,-5.57506608963013,
-4.54668998718262,-16.0420608520508,
-45.6715049743652,-17.2056694030762,
-51.8159904479981,12.8234043121338,
1.93995141983032,40.5837821960449,
59.1120910644531,29.3233337402344,
56.3279685974121,0.360221862792969,
3.07166385650635,8.07221603393555,
-31.5398712158203,55.3428001403809,
-22.5933380126953,84.1741714477539,
-18.0511741638184,62.8209609985352,
-45.3876838684082,17.7711906433105,
-70.1158828735352,-10.8276491165161,
-43.0364608764648,-18.1899318695068,
15.9091491699219,-22.2048301696777,
51.5638313293457,-21.3190174102783,
48.4142570495606,-1.50075578689575,
39.8088493347168,31.2395496368408,
42.9355392456055,44.0363082885742,
36.8022193908691,21.8356094360352,
13.8054847717285,-17.3495330810547,
6.91938018798828,-48.0629234313965,
33.4298782348633,-58.7665710449219,
56.3505630493164,-41.4579315185547,
27.4615955352783,-6.23037481307983,
-35.8783378601074,24.2015991210938,
-70.9154663085938,27.8095054626465,
-56.3484802246094,12.0334777832031,
-30.2400646209717,1.77386331558228,
-26.0244369506836,10.3674201965332,
-25.2659034729004,20.0766811370850,
-1.36682868003845,16.8406162261963,
34.5300292968750,10.4489898681641,
42.4132537841797,15.3741750717163,
15.8641767501831,17.8114776611328,
-5.57813549041748,-2.98653745651245,
3.86209726333618,-27.5784664154053,
27.5996742248535,-17.1894836425781,
29.6740779876709,29.7661094665527,
3.97067284584045,73.5778732299805,
-26.8377761840820,72.2723464965820,
-37.7709922790527,35.6329612731934,
-20.8076381683350,-0.586136460304260,
8.10284996032715,-17.2095222473145,
20.7109870910645,-16.2102031707764,
9.84745216369629,-0.148540973663330,
-14.2770671844482,25.7742214202881,
-26.2082862854004,36.8340644836426,
-18.5636386871338,7.15172052383423,
-5.48298406600952,-45.2442588806152,
-2.24567508697510,-59.1591377258301,
-7.43902778625488,-6.20020627975464,
-6.69906473159790,62.6368522644043,
-5.72108697891235,67.1212387084961,
-12.2270240783691,-1.58548641204834,
-17.5595588684082,-70.3746337890625,
-9.88997077941895,-71.7891921997070,
3.77389717102051,-18.2702465057373,
-2.23195791244507,21.8011817932129,
-35.2056045532227,10.7293739318848,
-67.1438903808594,-23.2028560638428,
-67.3063583374023,-36.5915679931641,
-41.1670265197754,-20.7472572326660,
-14.8507261276245,0.942233443260193,
4.07189369201660,11.9308271408081,
24.6544036865234,14.5399761199951,
39.6723747253418,18.0299968719482,
20.4376659393311,20.1266593933105,
-32.6075019836426,11.7380666732788,
-71.6940002441406,-7.55382490158081,
-50.1722908020020,-21.1711978912354,
13.4624118804932,-13.7399024963379,
58.2570648193359,4.49403572082520,
52.9638137817383,11.1731739044189,
29.7035160064697,-11.0780267715454,
26.6833686828613,-43.0537376403809,
41.0098457336426,-45.7873497009277,
37.7472686767578,-15.3996362686157,
5.35948467254639,8.62541580200195,
-25.1054821014404,-8.24866199493408,
-27.9232978820801,-50.5230178833008,
-11.6945438385010,-69.2455978393555,
-6.73307132720947,-42.7622489929199,
-18.6636199951172,-4.88419198989868,
-24.2190246582031,2.93889236450195,
-5.78741121292114,-12.7209568023682,
24.6516952514648,-19.9164009094238,
37.6582260131836,-16.2802734375000,
24.5921878814697,-26.3867378234863,
15.4120130538940,-57.0991096496582,
30.8581237792969,-71.6520996093750,
51.2925758361816,-41.1734848022461,
46.3392257690430,7.74292755126953,
18.2824382781982,21.3325138092041,
-0.696229696273804,-1.98330307006836,
4.32848119735718,-8.81229114532471,
6.42857170104981,26.9299201965332,
-16.7858657836914,54.9037780761719,
-41.0907173156738,20.2716178894043,
-29.6243171691895,-52.1673126220703,
3.59361410140991,-80.1376571655273,
12.6122293472290,-36.2092208862305,
-8.51965713500977,17.0869255065918,
-18.4742336273193,15.1793556213379,
5.51399612426758,-25.2195682525635,
25.6659259796143,-48.5766296386719,
2.42834901809692,-40.3627166748047,
-33.6733055114746,-33.6227569580078,
-22.5387096405029,-38.8696136474609,
32.5296058654785,-29.5326042175293,
59.5429687500000,5.32088232040405,
21.6504039764404,24.3874626159668,
-27.7663002014160,-4.02417469024658,
-16.2980957031250,-42.7074661254883,
46.0383453369141,-33.7096366882324,
78.4020462036133,23.0351123809814,
38.2617988586426,67.5591735839844,
-25.2414646148682,48.6568336486816,
-45.6067199707031,-9.13571453094482,
-17.6171607971191,-37.6231498718262,
9.59331798553467,-12.6469030380249,
4.59500122070313,27.6864051818848,
-9.86661052703857,36.0093955993652,
-3.24885559082031,10.1613254547119,
16.4734859466553,-11.4701499938965,
20.3415527343750,-0.129907488822937,
0.742403924465179,17.5345458984375,
-15.6889152526855,-0.0765299797058106,
-8.02688407897949,-52.6936073303223,
13.9022865295410,-82.0282516479492,
26.3616275787354,-45.5186767578125,
15.0162229537964,26.5765209197998,
-10.8312149047852,67.7087783813477,
-29.3211498260498,47.9138717651367,
-27.3538761138916,3.99317455291748,
0.768164932727814,-10.9127864837646,
39.5962753295898,5.73492431640625,
60.6423988342285,23.4960403442383,
50.5681152343750,26.6368064880371,
28.7815780639648,23.5465240478516,
27.0637912750244,25.0204887390137,
49.3361358642578,30.6946830749512,
62.3936576843262,32.8891334533691,
34.6456298828125,35.6471405029297,
-21.5214252471924,35.3764648437500,
-61.7226867675781,22.3880558013916,
-57.9131965637207,-8.75577068328857,
-24.7981452941895,-38.0638771057129,
9.25008964538574,-40.3107261657715,
25.7405242919922,-11.0891304016113,
29.3294048309326,25.4320964813232,
29.8078937530518,34.4797744750977,
28.7360382080078,10.4869213104248,
22.3597068786621,-18.5491275787354,
6.37671709060669,-20.7761516571045,
-19.8007564544678,2.55909490585327,
-42.8575363159180,20.4638061523438,
-45.8863868713379,4.14123249053955,
-20.9244537353516,-37.3299407958984,
10.7689857482910,-71.2321853637695,
22.7466983795166,-77.3699264526367,
14.6518096923828,-65.6424255371094,
14.4057197570801,-47.7478408813477,
35.9624023437500,-20.4723644256592,
56.5341186523438,16.6809806823730,
46.0147590637207,39.0526809692383,
13.0240802764893,24.3689403533936,
-4.70998477935791,-11.3536224365234,
6.11099243164063,-25.5175304412842,
20.7772026062012,-1.05312526226044,
14.4281673431396,32.7882156372070,
2.66215252876282,42.1797218322754,
7.53674793243408,29.8754920959473,
22.8201942443848,19.7763137817383,
20.1459293365479,17.3995075225830,
-1.79765212535858,9.05791187286377,
-10.4239149093628,-3.38933038711548,
9.91598510742188,-4.56916809082031,
34.5070533752441,10.3586044311523,
33.3681945800781,20.0233020782471,
8.07643795013428,14.1110744476318,
-11.2249050140381,8.68164348602295,
-9.16876697540283,20.2596168518066,
0.546654164791107,29.1788845062256,
6.51720619201660,9.97875022888184,
12.1028013229370,-26.0105686187744,
26.8129100799561,-34.0689620971680,
45.2652664184570,-1.80957841873169,
56.7018737792969,26.7473125457764,
50.7684936523438,8.81406211853027,
27.6499729156494,-30.6535320281982,
3.08440041542053,-30.2884674072266,
-8.17392158508301,24.2846889495850,
-8.62310981750488,73.5638046264648,
-14.2115173339844,59.3859329223633,
-32.7471008300781,-1.85658931732178,
-44.2245674133301,-43.0347404479981,
-23.5708484649658,-33.2258071899414,
19.4054355621338,-3.60945677757263,
46.9521026611328,9.91929244995117,
42.5672302246094,11.7267017364502,
32.7963104248047,24.8342819213867,
45.6134452819824,41.8345680236816,
60.2295036315918,36.4228286743164,
34.7813949584961,10.0952968597412,
-25.7346763610840,-10.4208841323853,
-68.4249343872070,-12.1926918029785,
-50.3525581359863,-13.9554462432861,
5.79883480072022,-31.3062725067139,
43.7397308349609,-49.5320320129395,
32.5554847717285,-46.0886154174805,
-4.48536062240601,-28.8031826019287,
-22.2854156494141,-20.2410697937012,
-0.830496430397034,-16.6061096191406,
39.2987098693848,0.799354851245880,
56.3949394226074,30.6348381042480,
26.9701805114746,45.7314224243164,
-25.3666362762451,28.3543014526367,
-48.9554939270020,-4.74929857254028,
-20.8464241027832,-21.8537750244141,
21.8517608642578,-16.7956447601318,
30.3942413330078,-9.16031360626221,
7.11917304992676,-8.57334709167481,
-10.8351430892944,-12.8622722625732,
-1.50806307792664,-16.9294967651367,
18.9071521759033,-16.4930305480957,
25.0678405761719,-4.57054519653320,
27.3763866424561,17.1854228973389,
40.5482063293457,34.3617362976074,
43.8953475952148,34.8435325622559,
12.5367536544800,23.8968887329102,
-34.6534347534180,13.9676570892334,
-47.8569602966309,2.59034252166748,
-18.9579868316650,-22.1166534423828,
4.19510459899902,-50.5465354919434,
-14.0665330886841,-49.0601844787598,
-37.6470260620117,-6.77640342712402,
-14.8102159500122,35.8270950317383,
38.5432968139648,38.0525550842285,
56.4181022644043,13.9210004806519,
10.2578258514404,8.74330997467041,
-47.3250045776367,35.5686836242676,
-56.5336265563965,61.4859008789063,
-26.7814121246338,59.1893272399902,
-11.9253129959106,38.0198478698731,
-29.4806041717529,17.6522102355957,
-49.8828086853027,-4.61777973175049,
-45.8842010498047,-32.3929748535156,
-26.6597824096680,-45.8997230529785,
-14.1579732894897,-22.7576103210449,
-11.7540092468262,15.8910856246948,
-8.02745246887207,29.3793144226074,
6.17331504821777,12.6429920196533,
27.8471145629883,1.42779433727264,
44.0668411254883,16.6433982849121,
44.8327484130859,33.7234725952148,
25.4198169708252,27.3269882202148,
0.939619898796082,11.6780252456665,
-3.68309903144836,16.3779449462891,
13.7584543228149,39.2156105041504,
22.5090122222900,45.6578483581543,
2.30193662643433,19.6053447723389,
-27.5657691955566,-13.4342489242554,
-34.0074348449707,-29.2667980194092,
-12.0735731124878,-33.7394447326660,
15.1830663681030,-39.3723335266113,
21.6894493103027,-38.1978302001953,
12.0533294677734,-19.7872982025147,
-7.12491989135742,-0.185624778270721,
-32.9409980773926,0.664848029613495,
-59.4582214355469,-16.4935779571533,
-65.9121017456055,-31.8841304779053,
-47.6096725463867,-35.5353393554688,
-30.2984085083008,-38.6928215026856,
-34.1646385192871,-44.9449462890625,
-34.3913459777832,-41.7825775146484,
2.91570639610291,-29.0159111022949,
57.2027626037598,-27.9300441741943,
68.4746398925781,-42.2507972717285,
18.7099037170410,-40.9999046325684,
-38.8916625976563,-11.3950662612915,
-41.0131492614746,14.7236776351929,
7.90808773040772,4.07404804229736,
51.4886131286621,-19.8712997436523,
61.9991569519043,-6.07397937774658,
58.4920806884766,40.6513786315918,
50.5070724487305,58.2681045532227,
29.3273468017578,14.5139884948730,
-0.976844131946564,-40.7669830322266,
-13.5059032440186,-46.2553215026856,
-1.76782011985779,-17.3750133514404,
2.97420406341553,-11.0447902679443,
-19.1198425292969,-33.7005844116211,
-30.7038822174072,-39.4492645263672,
3.78866338729858,-6.81259298324585,
52.7451591491699,32.2263526916504,
53.9318008422852,43.7535438537598,
2.93431663513184,36.7159461975098,
-27.6653099060059,32.9352569580078,
6.18758392333984,26.0215206146240,
49.9784507751465,5.10169458389282,
31.6384010314941,-12.6454992294312,
-35.3097877502441,-4.11422061920166,
-72.2547836303711,13.8606319427490,
-38.3490638732910,5.72395706176758,
19.8371582031250,-22.8376846313477,
35.0368728637695,-20.5491600036621,
-2.33828043937683,26.1661777496338,
-41.1921844482422,68.1462860107422,
-39.0343971252441,56.7849578857422,
-2.16883230209351,11.0396757125855,
29.5717582702637,-7.44817113876343,
29.5021476745605,23.8974552154541,
2.70607471466064,65.1117172241211,
-23.5852375030518,66.3846740722656,
-30.9058513641357,31.7885284423828,
-29.6785030364990,-6.13265991210938,
-35.9698104858398,-25.8722457885742,
-41.2719459533691,-29.6007461547852,
-19.0910968780518,-24.8326187133789,
24.8909015655518,-16.3796348571777,
53.0574493408203,-15.0822753906250,
37.1250877380371,-26.6785755157471,
-7.38044023513794,-41.2178153991699,
-35.5766143798828,-39.4573898315430,
-28.7761955261230,-19.1359653472900,
-10.5539684295654,7.55072402954102,
-8.42077541351318,28.0388145446777,
-22.1612720489502,46.3448486328125,
-34.6524429321289,63.1903533935547,
-35.0613365173340,61.8575973510742,
-19.5752677917480,31.1848564147949,
10.0673866271973,-2.69508481025696,
37.9291725158691,-7.99476337432861,
36.9239578247070,20.3638725280762,
2.71105575561523,49.7377853393555,
-35.2656173706055,51.3159751892090,
-38.2697639465332,32.9213676452637,
-12.4610166549683,18.5521736145020,
4.06753587722778,19.7130565643311,
-4.39532709121704,26.0457859039307,
-10.3280649185181,25.6730766296387,
13.9077720642090,14.5880584716797,
44.8081245422363,-4.41195487976074,
35.6720237731934,-22.0466766357422,
-13.9454154968262,-19.4576148986816,
-49.0511627197266,8.29126930236816,
-33.5489196777344,40.4606590270996,
5.48803758621216,49.5403137207031,
13.5293083190918,31.5838012695313,
-17.9138431549072,6.35939502716064,
-46.0768814086914,-9.92665386199951,
-34.9944915771484,-19.2866802215576,
1.99843442440033,-23.2747631072998,
24.7280864715576,-16.6851806640625,
18.5670433044434,4.06085109710693,
3.61134338378906,16.0737400054932,
0.991896152496338,1.77964806556702,
9.02260875701904,-22.4598140716553,
9.35942459106445,-21.1251716613770,
-8.32306098937988,4.08009624481201,
-33.5545616149902,16.5047569274902,
-37.9914894104004,-8.79395961761475,
-15.2215871810913,-50.8485221862793,
11.2741088867188,-69.9664916992188,
13.2967119216919,-53.1162796020508,
-12.2189655303955,-18.9108791351318,
-35.1979637145996,14.0750904083252,
-30.1371974945068,42.1510162353516,
-8.54365730285645,52.1034736633301,
-0.866763114929199,31.3009223937988,
-11.9483623504639,-5.02077865600586,
-21.7233715057373,-21.2775039672852,
-18.3639907836914,-7.91337490081787,
-11.1487388610840,-1.21525549888611,
-7.59609365463257,-26.7198753356934,
5.13247537612915,-52.6911926269531,
32.7102584838867,-33.3755226135254,
56.1267395019531,18.7923507690430,
46.0137443542481,39.7974510192871,
9.09669780731201,0.0418972969055176,
-16.8054847717285,-50.1683654785156,
-12.9869728088379,-44.4017105102539,
2.75465321540833,9.03388977050781,
7.68413448333740,49.3936271667481,
4.57709360122681,40.7043762207031,
6.14341688156128,10.6314125061035,
2.65238761901855,1.77670741081238,
-18.6748847961426,22.4301033020020,
-41.9406471252441,49.5272026062012,
-39.2471351623535,58.3210067749023,
-13.4222631454468,38.3779563903809,
-5.36505651473999,2.79814887046814,
-37.4006271362305,-25.4915809631348,
-72.2580871582031,-26.5051651000977,
-58.6023483276367,-5.71691036224365,
-1.69110250473022,11.7919931411743,
43.2742271423340,8.73954868316650,
41.1218070983887,-1.04767608642578,
9.38225841522217,-5.91227388381958,
-14.1306734085083,-14.3180351257324,
-16.0470199584961,-34.3876838684082,
-8.48296451568604,-52.5077667236328,
6.27847862243652,-54.0864677429199,
28.3402481079102,-45.3062210083008,
39.0345840454102,-45.5078086853027,
17.3605918884277,-47.2124404907227,
-21.7685031890869,-22.8717613220215,
-36.0861244201660,25.8463516235352,
-10.9125976562500,56.6586380004883,
11.8930778503418,38.6751556396484,
-0.364066243171692,-3.76553654670715,
-22.9863548278809,-17.7709655761719,
-8.78685188293457,9.61722755432129,
35.9361991882324,42.5050125122070,
52.8305892944336,49.8946609497070,
8.84556007385254,34.9042587280273,
-53.3153953552246,16.1325244903564,
-71.8221664428711,8.03342914581299,
-39.1626243591309,13.5698108673096,
1.67331957817078,20.6291160583496,
16.1464328765869,8.21133613586426,
10.6605138778687,-29.7325496673584,
5.89933872222900,-64.6811676025391,
12.7001171112061,-51.6703910827637,
32.8227195739746,7.61256122589111,
56.1189079284668,50.8631172180176,
59.8525238037109,28.6210346221924,
29.0307960510254,-27.7388381958008,
-20.4898872375488,-41.6191902160645,
-49.5965805053711,-3.49590778350830,
-36.7110939025879,23.5763587951660,
-2.34932231903076,0.867539882659912,
20.0011520385742,-29.4158859252930,
22.9082965850830,-7.79560422897339,
13.5746154785156,47.5980224609375,
-9.54693698883057,67.7261962890625,
-36.0795860290527,36.5307350158691,
-43.8540611267090,8.56277751922607,
-25.5983524322510,23.2832107543945,
-9.42564487457275,48.8281440734863,
-31.4723796844482,35.6552352905273,
-75.4841766357422,-9.55389785766602,
-86.6142654418945,-36.3194541931152,
-45.1284866333008,-31.7112178802490,
1.12131130695343,-24.3811798095703,
3.87031054496765,-28.8230228424072,
-20.7939929962158,-27.2252464294434,
-20.9704818725586,-3.09378790855408,
5.58717060089111,25.8821678161621,
11.8554706573486,27.7474689483643,
-17.8496761322022,-2.11920714378357,
-44.6550483703613,-34.9591903686523,
-26.5146179199219,-45.0716934204102,
21.6758460998535,-28.8420944213867,
53.6134834289551,4.48043060302734,
50.3643798828125,24.8412227630615,
27.3349456787109,8.37327861785889,
5.69345092773438,-30.9662532806397,
-3.57031297683716,-44.0706405639648,
9.20690822601318,-9.95088386535645,
43.7824630737305,31.0465354919434,
71.8906860351563,28.9401836395264,
50.0563354492188,-11.1489763259888,
-9.62475490570068,-33.0244636535645,
-45.0928306579590,-12.5805950164795,
-21.5347633361816,7.22873067855835,
25.2860450744629,-10.9318313598633,
43.8113937377930,-33.1703147888184,
27.4326381683350,-10.3963136672974,
8.20705604553223,35.3618011474609,
4.06543016433716,47.2117729187012,
1.96001732349396,18.4911041259766,
3.34112405776978,-3.50769472122192,
26.2459239959717,1.51995468139648,
53.4598121643066,-1.28810644149780,
42.6531639099121,-31.5711097717285,
-8.60419273376465,-45.2538337707520,
-39.4054718017578,-8.17016601562500,
-14.8702735900879,30.5135936737061,
22.4239444732666,6.49646759033203,
14.0087556838989,-53.7987594604492,
-18.2457485198975,-61.3715934753418,
-10.2647256851196,-1.65906858444214,
40.3132247924805,37.2434425354004,
61.0149612426758,-0.685706615447998,
12.9414825439453,-49.5634346008301,
-46.3614845275879,-26.1955280303955,
-48.9844512939453,41.4156417846680,
-8.88303470611572,53.4873619079590,
13.1006116867065,-14.0789985656738,
9.03213119506836,-70.2097015380859,
22.7306480407715,-36.2406158447266,
61.8879280090332,49.4134902954102,
74.9636917114258,89.5903091430664,
30.7749156951904,58.1061515808106,
-34.8269844055176,13.0748081207275,
-61.9999732971191,4.30583333969116,
-42.5324974060059,20.3621616363525,
-17.4192562103272,23.0552101135254,
-15.9714698791504,-1.49519538879395,
-25.5911140441895,-32.1879386901856,
-23.8718738555908,-38.1967353820801,
-11.0398855209351,-16.7834091186523,
4.81153535842896,5.73683500289917,
17.8905735015869,3.75841426849365,
15.5831508636475,-16.6801071166992,
-7.02224969863892,-22.9554557800293,
-31.4696063995361,7.61462688446045,
-30.9989948272705,48.7763900756836,
1.07152485847473,51.4662818908691,
37.5113029479981,19.0812549591064,
49.5086479187012,3.33012580871582,
30.4459877014160,28.0546264648438,
2.66817712783813,58.5932502746582,
-17.6070232391357,48.7711257934570,
-27.2903594970703,8.64380741119385,
-14.5276374816895,-13.2048568725586,
18.6678714752197,0.0681604146957398,
49.0308189392090,15.8250932693481,
46.3964233398438,7.73730134963989,
19.0740642547607,0.222470432519913,
8.61191558837891,12.9230175018311,
30.0108261108398,26.2077407836914,
48.9768524169922,6.90256452560425,
31.0309753417969,-29.9077396392822,
0.811981678009033,-39.6528205871582,
5.49879646301270,-14.2456541061401,
40.6200904846191,4.92140817642212,
46.9505920410156,-9.27344036102295,
-4.73678207397461,-32.9191436767578,
-60.4896469116211,-33.6543388366699,
-52.2092170715332,-18.3144340515137,
15.4464426040649,-11.5762596130371,
72.6691894531250,-10.9827527999878,
71.4691009521484,13.7550821304321,
27.8652019500732,60.3027648925781,
-12.9320354461670,86.6762161254883,
-33.7741050720215,71.5523300170898,
-41.5628890991211,43.6292610168457,
-46.3378601074219,34.7992858886719,
-42.9628906250000,39.7234268188477,
-25.9324645996094,27.4368953704834,
-2.44345521926880,-7.68712425231934,
15.7824077606201,-39.7757072448731,
16.3457450866699,-48.6123580932617,
-2.70207524299622,-38.4243316650391,
-20.8294811248779,-21.6925163269043,
-9.18377494812012,-1.74278163909912,
26.4276657104492,12.2041177749634,
45.1456184387207,3.10509943962097,
21.8306655883789,-18.2186279296875,
-23.9090728759766,-20.2066421508789,
-49.9488449096680,8.46302700042725,
-43.2191276550293,31.0400009155273,
-31.8528938293457,6.58423709869385,
-31.5204792022705,-47.1558799743652,
-23.8015804290772,-73.5353088378906,
2.18324804306030,-46.0785217285156,
21.3330898284912,2.02899074554443,
6.44933032989502,30.2609272003174,
-26.0807514190674,41.0886077880859,
-30.0835990905762,51.1279335021973,
1.65237545967102,48.1188430786133,
29.1352806091309,14.7929248809814,
16.1324291229248,-28.9451427459717,
-19.2650356292725,-32.1264114379883,
-36.9121475219727,12.0947933197021,
-23.1751537322998,52.5653305053711,
0.705223441123962,42.8274192810059,
9.93814277648926,-0.835722684860230,
8.94497680664063,-24.1991844177246,
11.3505544662476,-5.72504234313965,
18.9207820892334,25.3180446624756,
27.5085926055908,31.3125171661377,
26.2932929992676,15.3408632278442,
8.42953109741211,3.06923413276672,
-26.2955017089844,6.42184829711914,
-58.6488456726074,17.5125503540039,
-69.2848510742188,13.2698955535889,
-59.6511344909668,-14.6139411926270,
-48.0047874450684,-48.9946784973145,
-42.8757324218750,-57.9496726989746,
-27.9325714111328,-35.2334518432617,
12.0975971221924,-9.74133491516113,
53.0336723327637,-11.2302999496460,
50.3297080993652,-34.4497566223145,
8.43202209472656,-46.9069252014160,
-25.2057476043701,-33.4061393737793,
-13.7845640182495,-22.6947402954102,
20.7201194763184,-37.9717369079590,
35.4643402099609,-53.8894691467285,
25.5695209503174,-34.3918571472168,
21.7173652648926,9.19544410705566,
29.9247207641602,29.2884902954102,
24.3047485351563,10.0998716354370,
-1.35619068145752,-13.9300098419189,
-14.0576534271240,-6.31982374191284,
9.33964920043945,15.7670955657959,
27.9552612304688,17.6742362976074,
-3.81851100921631,-0.956286132335663,
-62.5490112304688,-16.2335300445557,
-74.7788467407227,-18.7577705383301,
-15.7477912902832,-24.8100471496582,
52.8861961364746,-38.3235206604004,
66.2252960205078,-34.9612045288086,
33.0831985473633,-5.69986057281494,
12.1292095184326,22.0656185150147,
27.2940635681152,23.1914062500000,
49.5123023986816,9.46248817443848,
50.3079414367676,10.2010002136230,
36.1959419250488,32.0900955200195,
16.4537334442139,56.0883102416992,
-6.34822702407837,65.3224945068359,
-22.9706859588623,55.3787040710449,
-13.8756275177002,29.1761131286621,
19.3721313476563,-2.03571510314941,
42.6629257202148,-13.4924077987671,
27.4470100402832,15.1268863677979,
-10.5032463073730,65.6908950805664,
-36.4900360107422,87.6004333496094,
-38.7821540832520,59.5538787841797,
-38.5638580322266,12.2375183105469,
-42.8482322692871,-12.9853496551514,
-33.7430496215820,-14.0239057540894,
-11.5557775497437,-16.3284854888916,
-4.01981639862061,-31.0022907257080,
-25.5897216796875,-43.9980468750000,
-49.1866378784180,-41.4559593200684,
-41.6383514404297,-27.3753242492676,
-8.45685386657715,-10.2861642837524,
10.5135707855225,8.41097831726074,
-1.30410981178284,20.4060974121094,
-24.7345790863037,10.0540056228638,
-32.6391677856445,-23.1995830535889,
-25.7840652465820,-49.7067413330078,
-17.3592681884766,-39.4317359924316,
-2.52601480484009,1.40769541263580,
23.2736358642578,33.7511024475098,
46.6727600097656,36.4262351989746,
50.0746154785156,15.4790964126587,
36.3924865722656,-4.62661647796631,
24.5741138458252,-9.99067020416260,
22.1786804199219,-3.27034282684326,
20.9493274688721,7.45191621780396,
11.2883138656616,12.4433279037476,
-3.75469064712524,2.60604333877563,
-21.2793846130371,-17.7518062591553,
-43.0212440490723,-31.0514926910400,
-58.7940864562988,-25.3397426605225,
-46.5260124206543,-8.58321571350098,
-5.19201898574829,4.53781366348267,
31.4037036895752,15.8290157318115,
39.0500793457031,29.0453128814697,
31.1482429504395,33.9771995544434,
37.8343811035156,24.1850337982178,
51.3870658874512,12.5067996978760,
38.8492584228516,23.0716285705566,
-0.556057929992676,55.1996116638184,
-25.9420337677002,66.8659591674805,
-8.45376586914063,29.7414264678955,
22.9968433380127,-25.3300952911377,
24.1638603210449,-49.9556083679199,
-3.06800913810730,-35.6151618957520,
-17.4765224456787,-19.3182086944580,
-4.69399404525757,-18.4318408966064,
6.91183567047119,-5.31126403808594,
-5.92069292068481,31.8825016021729,
-28.1997699737549,54.3771514892578,
-38.1633186340332,24.0749816894531,
-35.8450584411621,-30.1714096069336,
-30.0738086700439,-38.2927284240723,
-25.2507648468018,8.07924461364746,
-13.6524639129639,40.7394790649414,
2.67330455780029,5.46610116958618,
17.1580333709717,-53.5018959045410,
25.7341823577881,-56.5914840698242,
28.8805618286133,10.1560363769531,
19.6403598785400,76.8634948730469,
-3.01483607292175,84.5962982177734,
-15.9036569595337,39.5067710876465,
-1.25351142883301,-8.30157184600830,
21.2896575927734,-27.7002010345459,
17.8825340270996,-20.4578094482422,
-3.59122538566589,2.96111869812012,
-1.90292179584503,24.6384277343750,
36.3013534545898,31.1449470520020,
69.6180496215820,22.1952400207520,
51.2228012084961,21.6386184692383,
4.36760282516480,43.8826522827148,
-15.4630241394043,62.1145133972168,
5.27783489227295,46.2385673522949,
23.5555744171143,7.99970054626465,
11.2739753723145,-11.5896329879761,
-4.81524848937988,-1.73018872737885,
5.82666444778442,2.34723615646362,
28.7660980224609,-31.4312896728516,
30.5379066467285,-73.3945312500000,
16.3430557250977,-66.5070419311523,
16.2167816162109,-6.86110401153564,
33.3958969116211,55.2390136718750,
33.4983787536621,72.5734100341797,
-3.74970579147339,49.9739608764648,
-52.7165794372559,15.6340742111206,
-69.2653656005859,-13.5415325164795,
-46.6321487426758,-32.5082778930664,
-15.7905435562134,-37.3250732421875,
3.94533681869507,-27.4597301483154,
12.5201663970947,-11.3374958038330,
18.2113533020020,3.10853958129883,
29.1975116729736,15.9561977386475,
44.7946929931641,35.3626518249512,
51.3821983337402,51.4462471008301,
31.3717575073242,48.8206253051758,
-10.2041378021240,30.4347305297852,
-38.0179328918457,11.4057550430298,
-27.9467010498047,-9.18857383728027,
0.322894334793091,-42.7184562683106,
-0.790315508842468,-69.3770599365234,
-36.9388122558594,-58.4245872497559,
-54.4996376037598,-14.4882946014404,
-15.6810693740845,10.4239025115967,
37.8177871704102,-17.2378101348877,
44.1713905334473,-56.8664131164551,
-1.42303347587585,-41.7359848022461,
-42.2301788330078,24.9751510620117,
-39.6763267517090,66.0569305419922,
-9.90840816497803,43.0594253540039,
14.8113384246826,-2.05104446411133,
24.6320133209229,-17.0414161682129,
23.1578960418701,-11.5971927642822,
0.359871625900269,-20.7788085937500,
-35.6237335205078,-30.5323524475098,
-49.4982147216797,-6.14472866058350,
-16.8253402709961,36.1250305175781,
26.1989440917969,34.8737144470215,
22.7021980285645,-16.4223804473877,
-21.4868812561035,-45.7106170654297,
-44.1708984375000,-7.11444711685181,
-22.0099983215332,44.0496139526367,
3.72161340713501,29.5748329162598,
-5.85969781875610,-38.3078765869141,
-31.7174091339111,-77.3128585815430,
-26.0871925354004,-56.0727653503418,
12.4416208267212,-17.3721256256104,
39.8026275634766,6.84246397018433,
35.0859222412109,29.4243087768555,
15.8111171722412,61.8968811035156,
-4.43891382217407,72.0349578857422,
-32.2140922546387,32.5449295043945,
-54.5112800598145,-19.2793216705322,
-43.0045776367188,-30.7304916381836,
-3.30635595321655,-9.02902507781982,
12.4888420104980,-6.22277498245239,
-17.2824249267578,-32.1609497070313,
-48.1734695434570,-43.8059730529785,
-28.8931007385254,-24.3628044128418,
24.1999378204346,-3.91237401962280,
47.3982315063477,-0.142411485314369,
24.2769985198975,5.21814346313477,
1.79325187206268,24.7176876068115,
3.64831972122192,37.6553573608398,
-7.69736576080322,17.8716487884522,
-47.8158454895020,-12.9907827377319,
-67.0685272216797,-17.8600883483887,
-25.4989471435547,1.47765552997589,
37.7168083190918,12.0252285003662,
49.2950553894043,7.48923730850220,
11.3361730575562,11.6555938720703,
-1.39316308498383,24.2803783416748,
35.5321350097656,18.9855613708496,
60.4959831237793,-3.15454006195068,
26.2991027832031,-6.42681074142456,
-21.6357879638672,19.8250083923340,
-11.6791973114014,34.3365592956543,
37.2871971130371,8.58338546752930,
38.6673851013184,-27.3542137145996,
-24.1836738586426,-28.1848011016846,
-73.8931579589844,-5.94695186614990,
-44.5276985168457,-14.3697776794434,
28.7772521972656,-60.7141342163086,
66.4694747924805,-85.0657653808594,
48.9155654907227,-45.1949653625488,
23.8542995452881,20.8694381713867,
28.9396476745605,51.7675590515137,
43.3008308410645,33.5423507690430,
28.6576442718506,0.516157448291779,
-11.7671232223511,-16.1681976318359,
-44.4693222045898,-15.4928989410400,
-44.4475173950195,-1.10117685794830,
-16.6054420471191,21.2645397186279,
20.4234733581543,35.5466957092285,
41.9920463562012,21.3963088989258,
39.2038383483887,-15.9326848983765,
26.9822139739990,-40.5178985595703,
19.9137001037598,-29.8292427062988,
21.3896389007568,-9.49701309204102,
25.6376724243164,-16.3019313812256,
23.9000568389893,-47.3507232666016,
16.6269359588623,-61.2783241271973,
7.63537120819092,-41.2422180175781,
-3.72004127502441,-8.54964160919190,
-12.1910438537598,1.51913475990295,
-9.22441864013672,-16.7867889404297,
0.634971022605896,-36.8336219787598,
-2.51788806915283,-39.4490013122559,
-23.3972568511963,-30.3262405395508,
-35.1738166809082,-20.5807228088379,
-11.2585296630859,-15.6164417266846,
33.7118568420410,-12.6115741729736,
55.1286659240723,-9.04368877410889,
35.9331512451172,-2.47766184806824,
2.76663637161255,2.38054037094116,
-9.43537807464600,-6.43072223663330,
-5.73401927947998,-28.7453155517578,
-12.7204465866089,-45.3764915466309,
-33.4098968505859,-35.3338432312012,
-38.7334175109863,-6.60451459884644,
-13.1114959716797,11.8003616333008,
22.6215934753418,1.33899307250977,
39.5159988403320,-10.3884744644165,
34.4730072021484,6.27777910232544,
19.8754787445068,38.4311256408691,
3.25747585296631,43.6052093505859,
-16.4936408996582,15.2660417556763,
-27.1997547149658,-8.28085231781006,
-14.2643585205078,-0.124044120311737,
12.4189443588257,18.2486553192139,
28.1728878021240,12.8663082122803,
18.4793567657471,-5.62369966506958,
2.44014024734497,-3.66747236251831,
-2.16370940208435,15.7628030776978,
-0.456159472465515,11.2677078247070,
-5.01811695098877,-28.9307937622070,
-6.40867280960083,-62.8789291381836,
11.1674432754517,-47.4960937500000,
34.1083488464356,2.74787974357605,
30.2732257843018,36.6964416503906,
-10.2582378387451,34.9504470825195,
-55.9043579101563,19.3627948760986,
-66.2260360717773,6.79874134063721,
-42.1368026733398,-7.65442085266113,
-9.28605270385742,-30.4023017883301,
11.9000387191772,-47.5840415954590,
22.4304962158203,-41.3407249450684,
29.2682247161865,-18.5529670715332,
31.7207012176514,-4.81283664703369,
32.8924102783203,-9.74475002288818,
34.3507461547852,-17.1631832122803,
32.9307327270508,-9.13786983489990,
21.3351821899414,18.4692420959473,
5.66405963897705,50.4906730651856,
1.79279518127441,64.5799331665039,
15.8252439498901,49.0965538024902,
29.2535114288330,22.2589397430420,
18.9364013671875,13.4026985168457,
-15.7203588485718,32.3805999755859,
-48.1497497558594,55.0449142456055,
-54.0667762756348,50.6800384521484,
-37.3507614135742,21.7602310180664,
-9.32057476043701,1.19902658462524,
16.3493804931641,6.58670043945313,
30.5340366363525,17.4843826293945,
31.3047332763672,1.30093908309937,
25.7447204589844,-32.2454109191895,
25.3249111175537,-48.2249488830566,
32.7445678710938,-32.6371536254883,
35.9876670837402,-4.64224576950073,
23.3900966644287,8.02679061889648,
5.28172826766968,3.41065073013306,
3.17944407463074,-1.36633801460266,
14.9157476425171,2.43099784851074,
21.1350021362305,16.6674079895020,
17.6375255584717,32.8138389587402,
23.0295124053955,42.1453437805176,
43.4963645935059,32.8616409301758,
49.2554664611816,10.1426219940186,
17.0623645782471,1.91435611248016,
-29.3244895935059,26.9729309082031,
-40.7838478088379,61.6939506530762,
-14.0339231491089,61.3809127807617,
-0.246735721826553,16.5583953857422,
-31.9948425292969,-31.8541793823242,
-67.1951904296875,-46.7555732727051,
-49.4371719360352,-32.6698799133301,
13.7149991989136,-15.2099399566650,
50.9031143188477,1.46109580993652,
26.6000785827637,27.6666088104248,
-21.4040679931641,53.7626838684082,
-36.0427131652832,50.4244728088379,
-9.74816417694092,15.7125167846680,
19.9146022796631,-11.0928535461426,
23.6290016174316,2.28128528594971,
8.28409194946289,41.7888641357422,
-10.4960155487061,61.6686019897461,
-24.0801544189453,40.6143989562988,
-25.0375919342041,-1.41194915771484,
-9.14802837371826,-30.5747718811035,
13.9962444305420,-27.9601898193359,
28.0799064636230,0.0165574550628662,
33.5333557128906,24.2700843811035,
43.0161895751953,20.4067001342773,
51.3440742492676,-9.51669120788574,
36.7358093261719,-35.4872779846191,
-2.33122515678406,-32.8199272155762,
-30.6290016174316,-10.0526428222656,
-13.2882709503174,-2.97745943069458,
29.3653774261475,-28.1947822570801,
46.4849243164063,-59.3777809143066,
23.9184837341309,-66.3360214233398,
5.66613578796387,-41.7445907592773,
21.9791755676270,0.0279440879821777,
48.7308311462402,33.6762504577637,
41.8255310058594,39.3652458190918,
2.42206835746765,16.9881210327148,
-26.2664394378662,-13.2343502044678,
-16.0682506561279,-15.6787157058716,
17.0703201293945,16.9246253967285,
33.7304496765137,43.2342338562012,
23.1449890136719,18.6168193817139,
4.41633605957031,-41.1843719482422,
4.46759700775147,-67.4614257812500,
30.5429248809814,-24.8222198486328,
64.0597076416016,36.8048324584961,
68.0615005493164,50.6666336059570,
22.7389316558838,20.0786991119385,
-37.9393157958984,8.16289615631104,
-58.8485069274902,40.3715858459473,
-30.8091449737549,70.2431564331055,
-4.21954822540283,43.8244552612305,
-16.7593231201172,-16.7101078033447,
-38.8542480468750,-46.1068077087402,
-20.0244750976563,-25.9644603729248,
33.8854026794434,1.37205481529236,
57.9146270751953,4.43132686614990,
22.1242275238037,-3.54301238059998,
-22.9492874145508,0.512765049934387,
-20.7302227020264,4.99004411697388,
15.0013580322266,-5.63362836837769,
23.8708095550537,-16.8775577545166,
-12.4356460571289,-9.28264331817627,
-55.7426261901856,4.08258199691773,
-63.6783676147461,-10.1139354705811,
-38.1752853393555,-52.3620643615723,
-1.26337790489197,-80.2292556762695,
29.7482109069824,-68.5579071044922,
40.6177711486816,-38.9162902832031,
25.3969287872314,-16.8677387237549,
-7.62086486816406,4.52433443069458,
-30.3133983612061,34.8753509521484,
-25.4262962341309,57.6834411621094,
-7.59829425811768,49.2709579467773,
-2.47517156600952,19.8087310791016,
-2.86178350448608,4.58343696594238,
9.58233737945557,13.6786699295044,
29.6662979125977,20.7806015014648,
34.0988273620606,8.77344894409180,
15.6855163574219,-6.08182096481323,
-3.48091864585876,-6.75857162475586,
-1.57758581638336,-5.12277841567993,
20.5738906860352,-15.7574739456177,
41.4025611877441,-23.2308902740479,
51.2043685913086,-1.18520140647888,
48.2630653381348,35.2315254211426,
29.4014244079590,45.8895988464356,
1.10057020187378,12.1941766738892,
-15.8762359619141,-31.0255622863770,
-2.73237371444702,-40.6294937133789,
28.2426280975342,-19.3326034545898,
40.3509483337402,-0.692508041858673,
21.3451862335205,-3.21662807464600,
-6.66536426544189,-12.6875457763672,
-17.9586505889893,-7.99870920181274,
-16.5562953948975,6.95705890655518,
-21.1221370697022,14.5290670394897,
-35.2287139892578,5.27744007110596,
-35.7851333618164,-16.1901035308838,
-8.22934532165527,-30.8538894653320,
33.6287231445313,-20.9320831298828,
61.7371444702148,12.6907882690430,
63.4523849487305,45.5932083129883,
42.7071380615234,49.8562355041504,
18.0783538818359,17.0473575592041,
4.98462057113648,-28.5503101348877,
13.3993234634399,-51.5730400085449,
31.4469604492188,-41.1899337768555,
36.6704254150391,-8.65542125701904,
22.7532463073730,27.7567100524902,
5.75384235382080,44.1038703918457,
4.97567272186279,25.0735721588135,
20.8555374145508,-20.9156475067139,
30.2782020568848,-54.7061309814453,
23.6393547058105,-40.8526916503906,
13.9767713546753,5.93872451782227,
12.8534078598022,32.1108741760254,
16.1397933959961,13.6076917648315,
17.6385459899902,-12.8012752532959,
16.0958023071289,1.31129944324493,
8.55209732055664,44.3886718750000,
-11.4583015441895,56.5560607910156,
-40.9247894287109,13.0472183227539,
-49.9982681274414,-39.3910751342773,
-15.6967124938965,-42.0052757263184,
34.4146575927734,2.48218131065369,
41.2552490234375,44.9241523742676,
-10.6857900619507,46.2648162841797,
-67.5320892333984,16.4630432128906,
-60.9543075561523,-13.3683395385742,
7.39335441589356,-22.8674602508545,
62.9310035705566,-6.21691274642944,
49.7257575988770,29.7456016540527,
-10.5094203948975,59.8780059814453,
-53.7403831481934,50.9657821655273,
-45.0504684448242,0.975203037261963,
-6.31090879440308,-48.7782363891602,
19.7738342285156,-55.2613296508789,
23.5050182342529,-25.1164054870605,
25.3250656127930,5.79211807250977,
36.2131500244141,19.1722373962402,
38.4353675842285,26.6965942382813,
8.93878269195557,32.6720848083496,
-37.4709281921387,22.1772651672363,
-57.0228996276856,-10.4118337631226,
-23.7761783599854,-33.5280723571777,
29.4653472900391,-15.6503906250000,
36.5621299743652,23.4159278869629,
-12.4633598327637,39.0748596191406,
-57.8056449890137,13.8214397430420,
-46.0733375549316,-23.9352817535400,
7.11006450653076,-45.0236892700195,
39.2656173706055,-51.3546180725098,
21.8509216308594,-48.0132560729981,
-4.20744228363037,-27.1139259338379,
2.24089789390564,13.7171497344971,
21.7338619232178,56.3191108703613,
15.4319458007813,70.0961837768555,
-7.29431247711182,52.3000946044922,
-2.30119442939758,27.3335971832275,
33.6003417968750,12.8676862716675,
46.3152236938477,2.46711540222168,
6.68539619445801,-13.4984321594238,
-39.4596405029297,-31.6422920227051,
-30.4537315368652,-45.3899917602539,
15.6898708343506,-43.5817260742188,
26.2538490295410,-20.0740871429443,
-14.9384870529175,8.55992507934570,
-43.8707351684570,12.8044061660767,
-9.84886550903320,-12.8787040710449,
40.0086021423340,-37.3225021362305,
33.4334945678711,-18.5360431671143,
-20.5137500762939,28.8521080017090,
-46.7979698181152,47.3875541687012,
-10.0376672744751,13.2254600524902,
41.3573608398438,-20.4462795257568,
56.5260810852051,3.34471225738525,
44.8597984313965,54.9484863281250,
39.4939270019531,56.8175506591797,
36.6633644104004,-3.97421383857727,
13.8645048141480,-51.5113601684570,
-22.0598239898682,-29.1122989654541,
-33.1434211730957,22.6676559448242,
-16.0857505798340,22.1526355743408,
-12.7238893508911,-31.3835124969482,
-42.1716690063477,-67.0727844238281,
-66.9422454833984,-47.7097282409668,
-44.3645172119141,-12.1646728515625,
16.8461055755615,-8.50934123992920,
62.2866058349609,-21.8985671997070,
55.0541229248047,-4.34893560409546,
17.0490264892578,44.3827934265137,
-2.82641339302063,72.4359130859375,
7.85874843597412,56.3065605163574,
21.1898059844971,26.4495124816895,
6.48141765594482,17.5671043395996,
-31.5323429107666,21.0901966094971,
-52.6178131103516,0.652953386306763,
-30.7624664306641,-47.2100868225098,
14.3540735244751,-74.6327819824219,
33.9115715026856,-44.0140037536621,
10.7978401184082,19.0525894165039,
-22.9671058654785,55.0420875549316,
-25.8408432006836,37.4705200195313,
-3.41696929931641,-1.71116185188293,
8.35638427734375,-11.6703710556030,
-13.0232372283936,11.2096214294434,
-46.3785705566406,22.9084510803223,
-51.7922554016113,-6.41612148284912,
-23.6345672607422,-45.9920005798340,
12.5088729858398,-41.8346176147461,
28.7698116302490,10.7408094406128,
22.5955162048340,60.4361000061035,
7.40987110137939,56.0253715515137,
1.18527436256409,9.83159446716309,
5.84062290191650,-23.1501255035400,
12.4531097412109,-11.2703590393066,
6.47636556625366,17.1300544738770,
-18.8860569000244,24.9642925262451,
-45.2178153991699,13.0258836746216,
-43.0930824279785,4.74953031539917,
-5.76728343963623,11.0857095718384,
36.7735633850098,11.6105089187622,
43.6940040588379,-3.41487264633179,
18.2329120635986,-14.3830995559692,
5.81374311447144,-4.42472743988037,
32.8951416015625,16.3437461853027,
65.2312393188477,27.8028240203857,
51.3903770446777,26.8247909545898,
-10.2575044631958,24.1546821594238,
-66.3509826660156,20.3395195007324,
-74.4975051879883,0.914884805679321,
-47.3561363220215,-37.6061248779297,
-23.1503868103027,-65.3635864257813,
-11.2511730194092,-49.9778060913086,
0.526219606399536,4.07647466659546,
5.55231332778931,56.6049423217773,
-10.3671846389771,64.7749481201172,
-36.7503623962402,23.9855613708496,
-40.2231903076172,-26.7514953613281,
-7.51493167877197,-41.1451454162598,
30.6215305328369,-14.3961095809937,
40.7832221984863,17.5533466339111,
27.2086391448975,19.4450054168701,
15.3988428115845,-4.78795337677002,
11.4139242172241,-23.8737869262695,
10.1311826705933,-19.0192165374756,
15.2374305725098,-7.51292419433594,
37.0583076477051,-4.15531015396118,
57.7901229858398,-0.308684349060059,
38.0701293945313,14.3280754089355,
-20.3475379943848,26.6122531890869,
-59.2854995727539,13.2397327423096,
-28.5403385162354,-15.6583805084229,
40.9357299804688,-23.7227592468262,
72.4454498291016,4.41225194931030,
30.9111385345459,34.0830307006836,
-35.6132354736328,30.4511928558350,
-51.2423171997070,6.58624076843262,
-7.85366582870483,5.58154869079590,
35.6823959350586,38.0315170288086,
29.7177543640137,63.9287757873535,
-12.0249862670898,43.8722991943359,
-37.4977493286133,-2.53720784187317,
-20.7232456207275,-24.4871883392334,
9.94785022735596,-1.56891083717346,
6.94236087799072,36.3162956237793,
-27.7534065246582,49.5214118957520,
-43.1441535949707,33.4141120910645,
-1.31193065643311,9.95654869079590,
60.4797439575195,-3.23815345764160,
73.0116958618164,-4.61248254776001,
19.0592117309570,3.21937084197998,
-44.5561485290527,15.7263240814209,
-52.5304832458496,25.1388416290283,
-21.9715805053711,25.9812831878662,
-16.9691314697266,27.1303997039795,
-47.9403076171875,36.3771858215332,
-62.9522285461426,42.3425979614258,
-30.8330001831055,21.4454269409180,
7.30108356475830,-19.2280769348145,
-2.02371335029602,-44.5553855895996,
-41.9045829772949,-30.3046474456787,
-49.7781867980957,3.87353324890137,
-15.9885206222534,19.4894084930420,
3.43538570404053,10.7530183792114,
-24.1080875396729,9.75926399230957,
-49.9844284057617,30.8114223480225,
-20.6866989135742,50.3377952575684,
43.6626014709473,41.5991821289063,
66.7647247314453,8.75489425659180,
26.2504158020020,-14.9710140228271,
-22.3425388336182,-8.07779979705811,
-31.3639831542969,21.3117160797119,
-12.3068513870239,41.5944900512695,
-0.779422104358673,29.3379669189453,
0.629667699337006,-10.2093601226807,
11.4080238342285,-42.0010681152344,
34.4055862426758,-41.7537727355957,
48.8108558654785,-19.7131271362305,
43.1223754882813,-11.3076934814453,
33.1536712646484,-30.8433666229248,
29.4461002349854,-45.2124824523926,
26.1692314147949,-18.7392234802246,
22.9864368438721,31.6156139373779,
26.6803092956543,60.2235527038574,
29.5889339447022,50.7513465881348,
14.6822500228882,28.2158699035645,
-6.24711179733276,16.6622180938721,
-9.61869430541992,9.41178417205811,
8.61845397949219,-4.45033454895020,
23.7249736785889,-8.53114795684815,
16.5333023071289,17.8819904327393,
11.8365659713745,51.9423179626465,
31.6743984222412,51.7063179016113,
49.2255172729492,17.3717803955078,
23.7275810241699,-7.18591356277466,
-30.4666404724121,0.503503859043121,
-52.9653549194336,7.04983329772949,
-27.7407894134522,-17.6924629211426,
-3.80647897720337,-48.0049781799316,
-14.7471666336060,-33.3807678222656,
-27.1712551116943,15.3072328567505,
1.57638096809387,37.7941131591797,
44.9996757507324,9.91829204559326,
41.6851005554199,-16.7935657501221,
-17.0255851745605,2.01675868034363,
-69.2936553955078,37.0582656860352,
-66.6040954589844,30.5088043212891,
-27.9626026153564,-12.3340415954590,
0.779259085655212,-31.4228324890137,
10.6726245880127,-4.85865449905396,
17.0726852416992,16.7842864990234,
24.5523891448975,-2.23036217689514,
25.5548610687256,-30.6758136749268,
26.6212844848633,-15.0304183959961,
38.4949607849121,31.7143421173096,
52.2646675109863,52.4230270385742,
51.5976371765137,29.2600955963135,
38.7774963378906,7.33856582641602,
32.1813812255859,23.2656726837158,
36.4858322143555,48.1202850341797,
35.7178192138672,40.4054641723633,
19.2146263122559,8.89297866821289,
1.79702889919281,-8.89756488800049,
2.61298370361328,2.26104831695557,
15.2417182922363,19.3488464355469,
21.1209621429443,24.9393997192383,
9.89549636840820,30.0713481903076,
-10.1844329833984,50.1132240295410,
-28.6193580627441,66.8240890502930,
-39.6583709716797,52.5455818176270,
-41.4515838623047,10.2088479995728,
-39.7538833618164,-29.1029605865479,
-36.7113151550293,-38.6542015075684,
-31.3262271881104,-16.4844532012939,
-17.7168712615967,18.4509048461914,
-3.49578523635864,35.6766204833984,
0.509539008140564,20.8489780426025,
-7.73010349273682,-14.5601167678833,
-10.9667558670044,-42.3813781738281,
3.63286733627319,-42.9116744995117,
20.6179466247559,-30.6512355804443,
10.8009986877441,-34.5621566772461,
-24.0504951477051,-50.1055793762207,
-42.9977569580078,-45.3353500366211,
-22.2759590148926,-10.7123718261719,
18.8507423400879,21.3964424133301,
39.6062469482422,15.5068979263306,
26.7450466156006,-11.2601480484009,
3.27843976020813,-19.6047821044922,
-12.2102470397949,-5.93002080917358,
-20.2537708282471,-2.92738771438599,
-27.8412609100342,-24.7689228057861,
-22.6806240081787,-34.5183258056641,
-2.40847039222717,-2.45630645751953,
10.8297662734985,45.1895904541016,
-5.43666458129883,51.2351722717285,
-30.4840888977051,3.23714852333069,
-21.3428783416748,-49.1227111816406,
27.4110965728760,-58.0546417236328,
69.8359909057617,-22.6651535034180,
63.3918647766113,19.0154991149902,
23.0374031066895,33.6348876953125,
-3.63610100746155,9.66927433013916,
-1.01454949378967,-33.2110977172852,
6.27020931243897,-62.6293907165527,
6.28404235839844,-59.3407135009766,
18.6084880828857,-35.4067840576172,
45.1772804260254,-13.4977750778198,
54.8922729492188,-0.104821324348450,
31.8550567626953,21.1134014129639,
7.97190761566162,48.7474937438965,
19.1554851531982,54.9962081909180,
41.2654991149902,20.9389686584473,
19.9595565795898,-20.5253791809082,
-35.4151878356934,-25.9981632232666,
-56.5419960021973,-4.29880046844482,
-10.0578918457031,3.12438035011292,
46.0611953735352,-17.6337852478027,
40.4459762573242,-37.2624092102051,
-7.83591842651367,-31.7331523895264,
-27.4400157928467,-23.2263145446777,
-0.346914768218994,-36.4580993652344,
22.3141098022461,-58.8098487854004,
4.08342647552490,-56.9349746704102,
-21.0861244201660,-26.6156997680664,
-9.51358318328857,3.88681364059448,
21.0191192626953,22.3366889953613,
22.7330684661865,38.7845954895020,
-16.6518039703369,50.6093902587891,
-54.7478752136231,38.8736000061035,
-56.6166992187500,4.97342252731323,
-35.4127044677734,-12.7605590820313,
-16.7461624145508,9.44346046447754,
-5.96532344818115,45.1319313049316,
-0.115472622215748,52.4172592163086,
-2.32496500015259,35.9535980224609,
-14.9159669876099,33.6070327758789,
-35.6591224670410,57.3509292602539,
-50.1938285827637,68.6650085449219,
-42.8412971496582,44.3130798339844,
-13.4099836349487,13.9041252136230,
17.2672328948975,15.6240844726563,
22.1915874481201,32.3985137939453,
-5.95945262908936,27.1304168701172,
-37.5510711669922,-0.590830922126770,
-25.6940212249756,-14.4660081863403,
30.5504951477051,2.25662922859192,
74.5148468017578,18.6170749664307,
58.1082496643066,5.92427873611450,
11.1221847534180,-20.9206123352051,
-3.07898473739624,-35.4395751953125,
24.8230743408203,-36.9958648681641,
45.5808792114258,-38.6203193664551,
24.3374423980713,-31.5843887329102,
-7.55243062973023,-6.82740211486816,
-5.54288482666016,13.9918832778931,
21.8219623565674,1.41009998321533,
27.5147304534912,-25.6096038818359,
9.73026275634766,-26.5068759918213,
6.20711660385132,3.36362695693970,
30.3689823150635,15.9759950637817,
47.7619209289551,-11.9733428955078,
37.8833236694336,-39.1837806701660,
25.8628883361816,-14.6869039535522,
34.9799232482910,43.1667175292969,
37.2341880798340,70.2735748291016,
-4.91887998580933,44.1452484130859,
-61.9234924316406,6.72800636291504,
-72.0748596191406,-11.6243886947632,
-27.0147113800049,-15.5317287445068,
10.8048601150513,-20.6200027465820,
-6.33190441131592,-13.9538526535034,
-46.3829002380371,12.3942689895630,
-52.8785247802734,40.8140602111816,
-31.1070346832275,47.1290855407715,
-26.3685359954834,36.6262130737305,
-46.0653877258301,33.1666603088379,
-51.2107009887695,41.8960304260254,
-22.2340049743652,43.9138946533203,
8.91198730468750,33.2954750061035,
4.98386192321777,24.1070518493652,
-25.8221035003662,13.8301229476929,
-45.8878707885742,-16.0142841339111,
-37.6728401184082,-59.2179679870606,
-15.9953222274780,-82.3798980712891,
-0.922132730484009,-69.8976898193359,
2.31979107856751,-47.6742630004883,
-8.71413803100586,-43.7182769775391,
-27.0051536560059,-46.4343490600586,
-36.4930419921875,-28.0527954101563,
-27.3470916748047,2.24826622009277,
-16.1203689575195,7.54258298873901,
-15.6043062210083,-14.7740545272827,
-16.2878036499023,-20.1194744110107,
1.13069939613342,10.3535089492798,
32.3053283691406,35.5076332092285,
53.1039390563965,14.8064842224121,
49.8579216003418,-27.3258590698242,
41.4400062561035,-33.6968879699707,
42.7084426879883,6.05164146423340,
36.2451705932617,44.3038635253906,
7.62950325012207,47.3305664062500,
-21.4432048797607,34.5445671081543,
-23.3378753662109,32.0875358581543,
-11.5323781967163,32.4167785644531,
-21.0050582885742,17.0014572143555,
-49.3541030883789,-5.93029356002808,
-48.4090728759766,-11.1835527420044,
1.74474978446960,-4.98214769363403,
49.6921844482422,-15.0316381454468,
36.4151306152344,-36.5896034240723,
-24.4872169494629,-37.1704902648926,
-63.9727630615234,-3.51242589950562,
-45.0650177001953,36.6231384277344,
-5.84130525588989,46.6198272705078,
-2.27989172935486,26.2631072998047,
-27.4123191833496,5.22479915618897,
-42.9139099121094,4.96122074127197,
-31.1728687286377,16.8661003112793,
-15.9178714752197,25.9061145782471,
-19.8857116699219,21.6510410308838,
-34.6222724914551,-0.232975870370865,
-28.7236175537109,-24.8682594299316,
7.73361587524414,-20.8553657531738,
49.7766532897949,24.6755371093750,
59.8100318908691,72.2006683349609,
25.5421009063721,68.2166290283203,
-22.9778594970703,11.3035221099854,
-34.6250877380371,-44.5981445312500,
7.75957202911377,-50.7125587463379,
56.6353416442871,-14.8577022552490,
45.8490486145020,16.7675399780273,
-18.6251792907715,27.2067241668701,
-62.1825027465820,33.6866302490234,
-34.7092399597168,39.8130111694336,
19.5561313629150,33.5305404663086,
24.9390258789063,18.0693874359131,
-29.0711803436279,11.3563508987427,
-67.0286102294922,10.2817974090576,
-35.3392601013184,-9.55433750152588,
23.5930881500244,-44.3052787780762,
40.0908699035645,-43.6278533935547,
7.26980209350586,12.7900848388672,
-29.1679534912109,69.1082305908203,
-36.6251869201660,53.3145027160645,
-29.3392639160156,-22.5772171020508,
-24.4341526031494,-66.6778640747070,
-19.4576835632324,-29.0497188568115,
-16.2902622222900,32.3450508117676,
-22.3942985534668,43.3879165649414,
-24.4418277740479,8.58431625366211,
6.86546564102173,-13.3887968063355,
66.1020584106445,2.77460384368897,
93.8237762451172,25.2824554443359,
44.1602325439453,26.1742610931397,
-38.4291801452637,7.19974946975708,
-67.2449951171875,-16.4585132598877,
-24.0982856750488,-41.6657104492188,
24.6850891113281,-58.9915847778320,
33.7221870422363,-52.7464294433594,
20.9273548126221,-22.0041694641113,
18.2113056182861,0.897481441497803,
13.1447439193726,-8.62246990203857,
-21.6526470184326,-26.3850994110107,
-59.2919082641602,-21.0644550323486,
-49.2544860839844,1.93994164466858,
0.910145282745361,20.6878318786621,
28.0085353851318,28.5341968536377,
8.43311119079590,27.7777633666992,
-11.0602226257324,14.9540510177612,
6.17194032669067,-15.2131805419922,
29.6590881347656,-42.3240203857422,
20.1865653991699,-37.3078460693359,
1.15179824829102,-8.72862911224365,
12.9719572067261,-4.75412416458130,
41.7741050720215,-36.1108436584473,
34.3385581970215,-53.0158767700195,
-13.7249908447266,-17.8954200744629,
-40.6576919555664,30.9152755737305,
-14.3544111251831,36.2410812377930,
23.2946147918701,4.52864265441895,
23.2964191436768,-8.13025760650635,
5.17881584167481,10.5154247283936,
9.03395843505859,11.9999618530273,
22.1745376586914,-26.6162014007568,
12.4551134109497,-60.4239540100098,
-9.34773635864258,-40.9722061157227,
-1.34528040885925,3.29101872444153,
32.8350715637207,8.02630329132080,
38.9520683288574,-30.7720947265625,
-3.83956480026245,-51.6991195678711,
-46.0000801086426,-16.8331985473633,
-36.2128639221191,32.0170135498047,
2.23874592781067,39.8863677978516,
18.4730529785156,5.54116630554199,
13.9540843963623,-29.3613739013672,
30.1761684417725,-30.7257652282715,
62.6435356140137,-0.822134435176849,
61.1993141174316,36.7614135742188,
7.29504585266113,57.6106338500977,
-52.0199851989746,48.2773780822754,
-61.4750480651856,14.8415431976318,
-24.7633209228516,-17.5639953613281,
11.4174337387085,-24.2991199493408,
18.5365295410156,-9.62867355346680,
9.39602375030518,2.45083427429199,
-1.75166130065918,5.86920213699341,
-15.1909322738647,15.0780553817749,
-27.7710018157959,31.7961750030518,
-31.9202232360840,37.0432739257813,
-29.5669937133789,19.8687667846680,
-32.5796432495117,-7.81847429275513,
-35.2016792297363,-25.0283298492432,
-24.7536067962647,-28.0804443359375,
-0.735672473907471,-27.5626773834229,
11.6179904937744,-22.8214874267578,
1.24316966533661,-4.77959823608398,
-12.7498817443848,23.0808105468750,
-9.55154895782471,45.8649101257324,
-1.81008887290955,48.3225059509277,
-21.3537750244141,34.2403907775879,
-57.8197555541992,14.4683456420898,
-64.0593414306641,-6.40788888931274,
-15.0409011840820,-23.3980312347412,
48.1524353027344,-28.7329273223877,
67.1168441772461,-19.5500431060791,
35.2315254211426,-4.71056032180786,
6.28842878341675,3.73592782020569,
20.1365242004395,0.979282975196838,
57.3295173645020,-7.06674337387085,
64.8696899414063,-10.8855056762695,
24.5664939880371,-4.72392177581787,
-26.4436092376709,9.31646156311035,
-43.9119033813477,19.9699230194092,
-25.7017974853516,18.3686237335205,
-9.28135681152344,5.33380079269409,
-21.6061248779297,-9.84548950195313,
-49.2996406555176,-18.6850757598877,
-59.7603874206543,-27.1351680755615,
-37.6069602966309,-36.6497611999512,
2.23252773284912,-37.5675544738770,
33.1660919189453,-19.4245700836182,
43.9189186096191,9.89463996887207,
40.7556228637695,28.8741531372070,
32.7173500061035,28.7386302947998,
29.9002532958984,24.0430088043213,
32.9014396667481,23.2499160766602,
28.1314144134522,20.3589725494385,
8.31748676300049,6.31393718719482,
-20.4694271087647,-9.79324436187744,
-35.2364234924316,-8.33903694152832,
-17.4715671539307,9.40329742431641,
18.8809318542480,23.3299160003662,
44.6353187561035,19.9166984558105,
39.7239189147949,10.9441137313843,
18.0676441192627,14.2060642242432,
-0.304057240486145,26.4464473724365,
-11.3567667007446,34.2802085876465,
-26.8242530822754,24.6396007537842,
-45.9852981567383,-0.552167177200317,
-46.2038345336914,-36.9943084716797,
-8.59591293334961,-70.4256057739258,
49.0019226074219,-80.5921249389648,
73.6509933471680,-52.9307136535645,
41.9059600830078,-2.12486720085144,
-9.30238819122315,34.2033462524414,
-29.6819515228272,35.9648208618164,
-22.0644836425781,21.1756076812744,
-28.6768970489502,12.7207059860230,
-62.4889221191406,5.28387880325317,
-76.3644332885742,-17.5929718017578,
-29.9766502380371,-44.0984420776367,
35.8211479187012,-40.2097473144531,
53.2630653381348,1.03080534934998,
19.7390060424805,40.5288276672363,
-3.01016783714294,42.9209365844727,
12.4211530685425,24.3227157592773,
22.7585582733154,26.7589988708496,
-4.04494905471802,47.1605911254883,
-33.9062271118164,46.7463684082031,
-19.2969837188721,12.7902889251709,
13.5403270721436,-16.5174636840820,
4.37416028976440,-4.38079786300659,
-40.4546966552734,26.4836120605469,
-51.0387611389160,27.6563358306885,
4.71819496154785,-4.94552135467529,
63.9045524597168,-24.3900585174561,
59.4386825561523,-13.6004934310913,
6.91356182098389,-3.70097422599793,
-20.4937019348145,-19.1765327453613,
2.80095338821411,-32.4591674804688,
35.9477958679199,-8.91990756988525,
41.8891677856445,27.5863780975342,
28.9231948852539,20.4567546844482,
20.6738033294678,-33.7901077270508,
23.4025268554688,-68.6943664550781,
26.4122028350830,-41.6119232177734,
24.5014801025391,-3.46207356452942,
22.2633018493652,-17.4581203460693,
22.7311420440674,-62.1130523681641,
14.1883821487427,-55.9857139587402,
-8.58178138732910,21.5234222412109,
-30.3521823883057,87.0544128417969,
-34.5839309692383,74.3622741699219,
-12.3338508605957,24.6164760589600,
18.4408683776855,15.8399419784546,
23.5055999755859,45.1063880920410,
-5.59844207763672,39.2694549560547,
-28.4196186065674,-17.6714553833008,
-2.53191208839417,-53.2801399230957,
50.7717475891113,-14.8775329589844,
68.8916015625000,42.8051490783691,
28.5310897827148,34.1518898010254,
-12.6575145721436,-29.1690082550049,
3.32309770584106,-59.3438034057617,
55.0350914001465,-16.2505683898926,
63.4658470153809,50.8164520263672,
3.22366905212402,73.1611480712891,
-63.1596984863281,46.1585426330566,
-75.6806869506836,8.25782108306885,
-53.7363662719727,-10.8521223068237,
-45.3940620422363,-17.1066150665283,
-48.7135047912598,-17.9059581756592,
-26.3023090362549,-19.0159149169922,
23.2027206420898,-22.2687320709229,
49.1085395812988,-19.4815216064453,
22.2981796264648,9.06914329528809,
-19.8845634460449,54.3230705261231,
-35.7770919799805,73.6765747070313,
-35.5161972045898,42.9304351806641,
-46.8722381591797,-6.67807865142822,
-59.3861618041992,-23.4975280761719,
-31.7533035278320,1.64920830726624,
27.4238872528076,30.9539737701416,
54.2002716064453,32.2274360656738,
19.8813419342041,20.6632251739502,
-20.8848724365234,19.1072807312012,
-7.46371841430664,18.4472675323486,
46.1446418762207,6.40021991729736,
67.5378952026367,-1.20639932155609,
24.2571544647217,13.5488491058350,
-40.1318893432617,36.5895042419434,
-64.1482543945313,39.0194778442383,
-42.6877746582031,21.7744903564453,
-12.1532030105591,13.2003669738770,
0.328726559877396,21.4034805297852,
-7.94329357147217,23.8005352020264,
-26.4477787017822,12.3730783462524,
-35.9866790771484,7.92624330520630,
-20.2499923706055,26.5689105987549,
16.1984939575195,44.0202941894531,
41.6518402099609,26.6054573059082,
34.4532737731934,-14.9815654754639,
15.4229116439819,-30.8802585601807,
16.9624633789063,-3.84915971755981,
36.2129058837891,34.8844566345215,
32.0626258850098,45.8137130737305,
-12.6885499954224,29.0444259643555,
-59.8495674133301,9.99808502197266,
-64.5611038208008,3.40852594375610,
-29.1172294616699,2.37803411483765,
8.41363716125488,-4.68846893310547,
25.6921215057373,-11.3281068801880,
32.5225982666016,-9.16916275024414,
40.2880935668945,3.98006772994995,
35.9970474243164,16.6221351623535,
6.72680521011353,17.9377479553223,
-30.2017841339111,1.94296967983246,
-44.9654846191406,-26.5359039306641,
-27.9402904510498,-49.7150382995606,
-4.32110023498535,-53.1931991577148,
-7.49729871749878,-42.4652709960938,
-32.0306701660156,-31.5635509490967,
-44.7017898559570,-29.4273395538330,
-24.8055019378662,-28.2265052795410,
15.3367624282837,-14.1480865478516,
48.1273689270020,11.7419099807739,
57.1049270629883,37.4442901611328,
55.2057952880859,52.3090095520020,
47.4282798767090,52.5476493835449,
26.8483085632324,37.2129859924316,
-5.14385890960693,7.70115232467651,
-22.4401378631592,-17.4805984497070,
-1.55486738681793,-13.3019437789917,
32.7409400939941,22.7928066253662,
34.6551551818848,55.8378715515137,
-11.1044654846191,45.1308288574219,
-59.4412574768066,-8.61034774780273,
-54.4134941101074,-58.2434043884277,
-6.42319154739380,-62.7600975036621,
21.6393699645996,-29.7667961120605,
-3.97667264938355,2.84926486015320,
-50.7794799804688,11.7590608596802,
-66.5028228759766,5.30862760543823,
-46.0726089477539,-5.29611492156982,
-29.7753124237061,-19.4554767608643,
-32.3352890014648,-30.6928462982178,
-24.3765182495117,-31.0752182006836,
15.6582984924316,-14.2285861968994,
51.6444053649902,7.20237064361572,
32.5883369445801,23.7952041625977,
-26.7003421783447,33.6745719909668,
-56.3283500671387,36.3792114257813,
-22.3222389221191,24.7464580535889,
29.0762176513672,0.197886466979980,
32.2173194885254,-20.1470413208008,
-5.60200405120850,-18.7510375976563,
-23.6094379425049,-9.36075305938721,
2.89181017875671,-11.2953071594238,
32.0835342407227,-16.3694038391113,
25.0017013549805,0.925201952457428,
-6.58520984649658,36.2576980590820,
-24.2274360656738,59.8677101135254,
-25.5035209655762,55.6972236633301,
-33.9860267639160,44.0085296630859,
-52.8806800842285,46.0420646667481,
-56.2467117309570,49.7550430297852,
-36.5191116333008,31.8822898864746,
-17.6359214782715,5.52687644958496,
-18.4399833679199,-0.211220711469650,
-29.7869529724121,9.18217277526856,
-34.2831573486328,0.351160168647766,
-29.9472637176514,-31.3375988006592,
-34.2428359985352,-51.1447410583496,
-51.5418701171875,-40.4805107116699,
-64.2527618408203,-31.2247486114502,
-55.2053184509277,-51.2992172241211,
-23.8440780639648,-74.3763732910156,
11.8707132339478,-51.9256210327148,
27.6835079193115,7.71313381195068,
10.2936124801636,42.9309120178223,
-22.4017047882080,18.5750656127930,
-36.8775749206543,-26.0469608306885,
-24.4173069000244,-42.2830429077148,
-10.2329034805298,-30.4019145965576,
-12.4566907882690,-24.5774135589600,
-21.4253387451172,-25.5208168029785,
-9.78131866455078,-9.41575431823731,
20.9767436981201,24.0964355468750,
38.3380737304688,43.2965774536133,
25.3685626983643,32.7102279663086,
6.31878280639648,15.4046220779419,
2.48543167114258,17.0865650177002,
-3.79680061340332,30.0972385406494,
-33.1391792297363,28.6529769897461,
-57.2544212341309,7.03070974349976,
-29.1081981658936,-10.2927350997925,
40.4906997680664,-8.17265701293945,
75.4259338378906,6.69776916503906,
29.6481513977051,24.0798854827881,
-42.1193695068359,31.9828872680664,
-54.9417114257813,19.2279357910156,
-2.59903025627136,-6.40867900848389,
39.1713867187500,-26.7223072052002,
24.2314243316650,-27.5854034423828,
-9.08309459686279,-17.1264801025391,
-12.1412687301636,-10.5740146636963,
0.419955521821976,-9.07642173767090,
-10.2905864715576,-6.25334739685059,
-33.6230354309082,-6.41270112991333,
-24.7206516265869,-24.7277355194092,
16.4906501770020,-46.3987159729004,
37.6075096130371,-30.3750877380371,
8.55090522766113,23.6894817352295,
-33.8044509887695,58.1628532409668,
-43.5930023193359,24.4076652526855,
-22.9448661804199,-45.7881126403809,
-6.05626392364502,-75.9584274291992,
1.59174966812134,-39.4845848083496,
13.4485073089600,9.78517150878906,
19.0805416107178,21.0427913665772,
2.30987596511841,6.37218570709229,
-21.9092102050781,1.55635023117065,
-18.5726184844971,7.34786844253540,
15.6754283905029,-5.80708885192871,
43.2934379577637,-34.9925079345703,
37.1207847595215,-39.5080261230469,
19.6929168701172,-3.59651708602905,
27.6779441833496,37.6515083312988,
55.0814056396484,44.2542076110840,
64.2476730346680,21.2931766510010,
44.0923423767090,7.27080726623535,
16.8915729522705,17.2607765197754,
-1.68784236907959,34.5191078186035,
-11.2255382537842,33.1544189453125,
-18.3354701995850,7.35838317871094,
-17.7576694488525,-24.4807682037354,
-5.52688837051392,-45.2137680053711,
12.4022235870361,-47.2827682495117,
27.9647674560547,-32.3350257873535,
40.1382255554199,-16.0962638854980,
43.5294456481934,-13.1079502105713,
26.2767105102539,-25.9307250976563,
-10.1872463226318,-38.2803230285645,
-36.9925270080566,-33.3229942321777,
-26.8100624084473,-8.61480903625488,
2.72956323623657,26.0921688079834,
7.45473670959473,47.9450454711914,
-24.6934719085693,42.3058929443359,
-58.0877838134766,12.6050443649292,
-52.6301994323731,-14.2993249893188,
-19.8264122009277,-15.1013936996460,
-2.93692731857300,8.01330375671387,
-19.1255264282227,33.8319587707520,
-38.9140548706055,48.3925743103027,
-31.5863113403320,54.0459022521973,
-5.36163425445557,47.3295745849609,
7.89322280883789,22.4529819488525,
1.40405130386353,-17.1231594085693,
-7.52598142623901,-42.7527122497559,
-1.42897510528564,-31.7828216552734,
7.81764268875122,3.67946386337280,
5.78588342666626,30.5051574707031,
-3.86289811134338,39.2480506896973,
-7.32772302627564,40.4275169372559,
1.06534266471863,37.1625289916992,
12.2660083770752,18.5645637512207,
18.2393627166748,-10.8635377883911,
23.7957649230957,-31.3534107208252,
28.4370632171631,-30.8515758514404,
30.6001091003418,-26.8668251037598,
31.8414001464844,-34.7144546508789,
40.5148429870606,-43.8961906433106,
54.6667594909668,-33.8712997436523,
57.0277748107910,-15.5499095916748,
33.0460395812988,-12.2552766799927,
-6.33953237533569,-20.3685798645020,
-32.5076217651367,-13.3416872024536,
-28.5660591125488,14.4784612655640,
-6.14779090881348,29.8632450103760,
11.0245466232300,12.9821681976318,
14.3287296295166,-10.2562074661255,
6.85942506790161,1.61955881118774,
-6.07514667510986,45.9581680297852,
-19.7024154663086,74.7867813110352,
-30.3747406005859,62.6312942504883,
-30.3334217071533,33.1582107543945,
-15.5104932785034,20.3572196960449,
11.0943384170532,21.1267700195313,
30.5396385192871,6.10713577270508,
25.2330017089844,-26.1097602844238,
0.195037364959717,-37.8732795715332,
-14.1403627395630,-9.40059757232666,
-1.03750348091125,28.3574886322022,
21.8776016235352,29.7867870330811,
15.7665424346924,5.24658298492432,
-22.6310882568359,0.917834997177124,
-49.6691932678223,30.6269207000732,
-33.5713310241699,46.3570365905762,
6.00127458572388,4.48307132720947,
26.2060585021973,-57.6769905090332,
18.3200016021729,-64.1131286621094,
12.2189569473267,-3.96226358413696,
21.5851612091064,58.0137481689453,
22.4603099822998,62.3197631835938,
-2.59168958663940,31.2307605743408,
-27.8791065216064,11.6409606933594,
-19.7265014648438,5.88794994354248,
16.6619033813477,-19.3236274719238,
38.3591270446777,-58.5596580505371,
18.6317310333252,-61.2221527099609,
-18.0713958740234,-10.4204883575439,
-30.7494182586670,41.8364982604981,
-8.77192211151123,39.8757286071777,
19.2615451812744,-5.16060638427734,
20.9405994415283,-34.7438011169434,
-2.02927803993225,-22.6193180084229,
-20.5011405944824,5.10178422927856,
-6.28349876403809,18.2040596008301,
30.2759475708008,24.1090965270996,
45.6534996032715,41.2255477905273,
14.4563875198364,58.4716796875000,
-40.3839492797852,52.6832237243652,
-68.9174423217773,26.0500545501709,
-44.1882019042969,6.04472970962524,
9.39813423156738,7.01963233947754,
45.7031364440918,13.0392580032349,
44.8020133972168,0.577388286590576,
24.4952774047852,-22.2631816864014,
10.2529792785645,-25.1330299377441,
10.0899257659912,-4.42401981353760,
19.8972663879395,10.0712718963623,
29.4710731506348,-1.70880079269409,
31.6675415039063,-20.4044685363770,
17.7099819183350,-8.77482223510742,
-12.8843984603882,34.5491981506348,
-43.3265876770020,58.8729362487793,
-47.7866516113281,23.3929939270020,
-19.7869434356689,-44.8141632080078,
17.3694553375244,-73.8274154663086,
34.3453216552734,-32.4057617187500,
24.7804145812988,38.2024345397949,
6.34286499023438,71.1817474365234,
-10.0088853836060,49.6910667419434,
-27.6135311126709,13.1812286376953,
-46.3589096069336,-1.80815112590790,
-54.6457481384277,0.167425706982613,
-39.1620063781738,-3.22257208824158,
-9.64092063903809,-11.7019462585449,
15.8677568435669,-8.97957801818848,
28.0109291076660,8.61933231353760,
31.4334926605225,21.1653537750244,
24.1679077148438,10.5845384597778,
1.04591655731201,-11.9063167572021,
-27.8892040252686,-22.6422424316406,
-35.4891166687012,-14.0358772277832,
-11.4905233383179,-0.248958677053452,
20.5634574890137,1.29305553436279,
31.1503467559814,-11.8039360046387,
13.8737716674805,-23.7520503997803,
-5.02507114410400,-20.0831813812256,
0.149561583995819,-8.25514793395996,
25.0901317596436,3.27757263183594,
45.8987426757813,7.66976547241211,
38.9868736267090,10.9310798645020,
7.93502521514893,20.6142387390137,
-26.1673183441162,28.9718761444092,
-31.4085845947266,14.3762168884277,
-4.41051292419434,-24.4402236938477,
18.3069515228272,-54.8493118286133,
9.68506813049316,-39.0798530578613,
-13.3828525543213,14.4113502502441,
-5.44721460342407,54.2382469177246,
34.4839057922363,40.6245841979981,
56.0867118835449,3.27032804489136,
25.0868701934814,3.20813512802124,
-27.2590370178223,47.7883720397949,
-41.9375267028809,79.4139175415039,
-23.4706592559814,54.9963226318359,
-24.5972251892090,5.83724308013916,
-56.8683395385742,-9.89787864685059,
-67.6099395751953,9.52811717987061,
-24.0453872680664,10.8024349212646,
28.8551769256592,-27.7697772979736,
24.9565505981445,-60.2806854248047,
-27.7026748657227,-44.0691413879395,
-63.9059257507324,-6.28939151763916,
-51.9642791748047,-3.43992328643799,
-25.4422588348389,-37.8396453857422,
-14.2300577163696,-55.3274879455566,
-2.27801060676575,-24.8847827911377,
31.5068206787109,17.3367252349854,
67.6235733032227,29.1046371459961,
63.0223159790039,16.1773796081543,
20.3581085205078,13.5427198410034,
-17.1346244812012,28.9346656799316,
-23.9038448333740,35.8179359436035,
-13.1505184173584,13.3849449157715,
-8.38718891143799,-18.7082347869873,
-10.6569528579712,-30.4908733367920,
-15.3124341964722,-15.0199317932129,
-19.6937103271484,9.62090492248535,
-30.1219921112061,20.1678829193115,
-44.3444442749023,7.04923486709595,
-48.8531303405762,-22.6615180969238,
-36.6628189086914,-37.9748001098633,
-10.0198011398315,-14.4561357498169,
20.6899299621582,30.3246650695801,
39.7879562377930,48.2814979553223,
36.0780715942383,17.0103263854980,
17.2888927459717,-32.9297714233398,
6.21658134460449,-46.3359756469727,
8.68579006195068,-13.3480167388916,
7.25750637054443,23.2691783905029,
-13.8612298965454,28.2822666168213,
-37.6530685424805,15.6159620285034,
-29.3847522735596,13.9791736602783,
12.9076604843140,26.6039485931397,
50.9768753051758,36.7723617553711,
43.4765510559082,35.6012992858887,
-6.25198268890381,27.7040462493897,
-56.0212173461914,13.7683010101318,
-68.5438232421875,-12.6298398971558,
-49.6512451171875,-33.7683639526367,
-24.8092041015625,-19.7980880737305,
-17.5847797393799,23.7017993927002,
-25.8024139404297,50.6938781738281,
-26.4132556915283,26.9028625488281,
-4.40186691284180,-22.1342449188232,
25.6594810485840,-36.3854446411133,
30.8063583374023,-5.29417181015015,
-1.88059401512146,26.3636341094971,
-42.8380355834961,19.9991397857666,
-50.5413398742676,-7.73253726959229,
-21.8809471130371,-15.1639614105225,
3.51468324661255,1.26806950569153,
-4.56467294692993,7.17330932617188,
-22.4675598144531,-19.8792514801025,
-4.90689849853516,-54.3654708862305,
43.1918601989746,-55.0245742797852,
66.7268981933594,-17.3103466033936,
34.7785415649414,20.9851989746094,
-20.8642253875732,22.9879398345947,
-40.4541130065918,-5.83351230621338,
-18.7537460327148,-34.6272506713867,
1.34925079345703,-38.0990409851074,
-3.95243334770203,-27.6391811370850,
-7.99282789230347,-24.1359176635742,
11.4211311340332,-25.6673698425293,
32.6868476867676,-12.7958278656006,
24.5619831085205,11.6379289627075,
-1.83369302749634,22.5452556610107,
-1.18653726577759,7.73410129547119,
29.3358612060547,-9.39038848876953,
47.0276603698731,1.29248893260956,
25.9615287780762,32.2493743896484,
-5.11282014846802,44.4977455139160,
-3.47061729431152,24.0368938446045,
24.0649299621582,4.76125049591064,
40.8649330139160,16.6024017333984,
32.2930984497070,42.6453208923340,
23.5581512451172,48.8032913208008,
30.2526092529297,32.1384735107422,
33.8508605957031,25.8234386444092,
16.8714141845703,39.8042869567871,
-14.0866641998291,48.3434944152832,
-40.6005668640137,24.9514312744141,
-54.3213424682617,-8.93012619018555,
-48.3256568908691,-15.2564105987549,
-22.6341514587402,9.95386409759522,
12.5065860748291,37.7342147827148,
28.8691806793213,42.9503364562988,
7.52857542037964,32.8910751342773,
-31.7036724090576,22.8615016937256,
-48.5648994445801,8.91904163360596,
-35.6955299377441,-17.8300552368164,
-15.7526569366455,-43.3387031555176,
-5.05374765396118,-49.3993911743164,
4.00632286071777,-35.5400047302246,
14.3208646774292,-26.0411682128906,
14.2840204238892,-37.5218887329102,
5.05412149429321,-59.6533317565918,
12.6308832168579,-63.1529388427734,
49.8995552062988,-32.4952964782715,
81.0122451782227,17.1369323730469,
59.6989212036133,53.6084823608398,
-2.93022704124451,50.3749618530273,
-42.8359375000000,11.9036216735840,
-22.2538871765137,-27.2333393096924,
22.6446094512939,-31.3576908111572,
29.0565032958984,-9.16263580322266,
-9.50033187866211,3.90053272247314,
-44.6353492736816,-14.1297655105591,
-39.1722564697266,-41.6424484252930,
-5.55717134475708,-43.7638778686523,
15.6410074234009,-19.7330741882324,
7.98981952667236,-6.79842376708984,
-9.95071792602539,-23.9024105072022,
-12.5891895294189,-43.7657432556152,
6.70327091217041,-31.6771106719971,
32.0668601989746,-0.655266404151917,
44.3466529846191,18.3696784973145,
43.2668685913086,18.9189796447754,
36.0846290588379,25.9839420318604,
33.5859146118164,54.1033706665039,
32.9521064758301,68.3250885009766,
22.9302120208740,44.3737487792969,
3.58008623123169,10.6215696334839,
-15.6517505645752,8.23568534851074,
-22.4318904876709,26.4258861541748,
-14.5856409072876,12.7367038726807,
0.803987860679627,-39.8432579040527,
7.77643871307373,-74.8115234375000,
-6.99638891220093,-48.7800292968750,
-32.4216499328613,-5.69103527069092,
-40.9552230834961,-14.1830434799194,
-13.1663570404053,-60.9017105102539,
28.4788932800293,-67.7911148071289,
44.6114692687988,3.90612745285034,
24.5595626831055,87.2045059204102,
-6.95487117767334,98.9162597656250,
-20.6200046539307,42.8553009033203,
-25.4622173309326,-7.94087553024292,
-35.8656082153320,-8.73585033416748,
-38.6391868591309,14.2443714141846,
-10.2798452377319,24.8745098114014,
31.8401279449463,24.8195037841797,
39.0752220153809,35.1954269409180,
-6.82710599899292,51.1912193298340,
-64.3429489135742,49.0233650207520,
-78.6168441772461,16.1588439941406,
-53.7300720214844,-30.2834739685059,
-36.2951698303223,-60.7948684692383,
-43.4478569030762,-69.3810882568359,
-41.4948692321777,-61.2999191284180,
0.861152410507202,-43.5776062011719,
54.8423004150391,-27.1709957122803,
65.2100372314453,-18.5615863800049,
23.5239334106445,-17.4646682739258,
-18.1990032196045,-22.1378440856934,
-18.9000682830811,-23.1017436981201,
3.99538135528564,-10.4990329742432,
3.44359731674194,11.2071514129639,
-23.1305675506592,21.7448139190674,
-32.0476799011231,2.28164792060852,
-1.35927033424377,-37.9430580139160,
39.5329322814941,-56.2967224121094,
47.2643852233887,-25.4046325683594,
21.0584964752197,35.4321250915527,
-6.76828527450562,68.3376693725586,
-24.8601436614990,46.2955245971680,
-39.7711143493652,-1.88435578346252,
-52.3925285339356,-32.0249328613281,
-46.2770195007324,-31.5146713256836,
-25.5001239776611,-21.8566703796387,
-16.9610633850098,-23.0516624450684,
-28.8352203369141,-31.6169662475586,
-28.0041751861572,-34.6322708129883,
11.7476320266724,-24.3798370361328,
60.4418907165527,-3.65480279922485,
67.2620315551758,21.6548233032227,
30.0302581787109,36.0954971313477,
-4.23692274093628,23.7551250457764,
-7.04666519165039,-10.5466203689575,
4.51015949249268,-45.7026710510254,
5.33997821807861,-55.7662277221680,
4.95228910446167,-33.6124229431152,
25.7354850769043,2.05069088935852,
52.4132385253906,26.3041267395020,
47.9539260864258,29.2483825683594,
8.05027580261231,15.2210636138916,
-31.1110401153564,4.59989690780640,
-42.4419212341309,4.91634225845337,
-24.9305133819580,2.90009236335754,
0.495656788349152,-18.1987533569336,
15.8287525177002,-42.0649719238281,
6.59847211837769,-35.1371574401856,
-27.6253795623779,5.58591032028198,
-58.0606346130371,34.1609077453613,
-50.7324752807617,5.09207582473755,
-3.67119908332825,-57.9482994079590,
32.7740554809570,-85.9770965576172,
21.2893772125244,-45.9248428344727,
-11.0783920288086,14.0391330718994,
-9.13503265380859,26.0843639373779,
29.4878425598145,-9.45215606689453,
42.7337112426758,-37.8772964477539,
-3.14882016181946,-29.7739219665527,
-63.4898223876953,-10.1010284423828,
-76.3511734008789,-12.4677305221558,
-36.2743110656738,-26.3839530944824,
5.99676418304443,-14.9130477905273,
16.5212669372559,23.0579395294189,
13.0481033325195,48.5767059326172,
22.7163486480713,45.4631729125977,
40.0378074645996,34.3870544433594,
38.0795783996582,32.6045188903809,
7.80589485168457,29.1525535583496,
-27.0700740814209,6.74903249740601,
-35.0297317504883,-15.5280742645264,
-4.35773611068726,-7.89219427108765,
46.5729942321777,10.7367124557495,
74.1412734985352,-2.39764785766602,
52.6611785888672,-46.5108757019043,
2.72077894210815,-59.7025222778320,
-24.0101432800293,-6.97500753402710,
-7.30777406692505,55.3362579345703,
25.8670215606689,44.3066101074219,
33.5503921508789,-30.2007808685303,
15.2602024078369,-71.9629440307617,
0.682846665382385,-23.6373004913330,
8.85178470611572,60.0707511901856,
24.7085933685303,88.6633987426758,
23.6228961944580,43.2802085876465,
5.73876619338989,-14.2982625961304,
-15.8977985382080,-34.8104896545410,
-27.9463272094727,-22.7956714630127,
-28.6055679321289,-3.93346166610718,
-26.7672443389893,15.5999126434326,
-32.4704208374023,32.4878158569336,
-44.3153190612793,34.5028572082520,
-45.6920661926270,22.4875659942627,
-22.5873470306397,19.8137493133545,
5.64277267456055,33.6275329589844,
2.75514411926270,38.1912651062012,
-34.2320251464844,18.3875808715820,
-62.9025459289551,-8.44357204437256,
-40.3921051025391,-10.6844396591187,
16.5734558105469,11.2476644515991,
50.0041427612305,23.0608177185059,
36.7299957275391,13.0986986160278,
17.0256710052490,7.27103424072266,
25.1104202270508,12.6573534011841,
44.5455436706543,6.90665578842163,
39.2281494140625,-12.8534994125366,
8.79024696350098,-19.3958396911621,
-11.4446325302124,-3.83644151687622,
-4.08259105682373,-1.84984588623047,
11.3466739654541,-33.6898689270020,
17.2943668365479,-56.9733886718750,
25.7449760437012,-23.9783420562744,
37.1082534790039,38.0188598632813,
28.5548229217529,54.4098052978516,
-7.99640560150147,8.93298053741455,
-31.7177295684814,-28.4794673919678,
-2.32093334197998,-14.3625974655151,
52.3893394470215,5.40407514572144,
63.1653060913086,-16.7766799926758,
19.3984642028809,-42.1885719299316,
-18.0560436248779,-15.6713571548462,
-4.85787343978882,38.7371139526367,
21.4553680419922,50.7188529968262,
4.95913267135620,13.9797811508179,
-42.8063392639160,-7.36321163177490,
-51.9798889160156,16.2856063842773,
-4.45405149459839,33.8713645935059,
41.6025962829590,8.15391445159912,
39.3485527038574,-14.4473743438721,
9.98260974884033,12.9280538558960,
4.09739637374878,51.0368728637695,
29.9693164825439,34.3724822998047,
55.8177032470703,-13.9186296463013,
54.4710922241211,-13.8938655853271,
29.0387344360352,39.2218284606934,
-4.63923263549805,61.1885185241699,
-25.8446426391602,10.3884801864624,
-17.3095989227295,-44.3242874145508,
20.2795352935791,-27.9382476806641,
49.3585128784180,33.3355216979981,
31.3484115600586,50.4857406616211,
-18.3120861053467,5.27874183654785,
-36.8653297424316,-29.4068889617920,
1.03313410282135,-6.52856397628784,
48.8772697448731,32.3553504943848,
49.3464813232422,29.5609474182129,
10.4334201812744,-8.70611476898193,
-11.9554538726807,-36.3903770446777,
11.9622592926025,-30.2449493408203,
48.3329315185547,-3.16132760047913,
50.9256324768066,20.5999107360840,
21.3954010009766,24.9121227264404,
-6.01907062530518,6.96723079681397,
-7.86606550216675,-24.6872348785400,
6.98295879364014,-50.7255439758301,
19.5089416503906,-53.4161643981934,
20.9367866516113,-39.3611602783203,
10.7355861663818,-31.2389030456543,
-9.86880588531494,-26.5110454559326,
-31.6070842742920,-7.39004182815552,
-46.2414741516113,19.7232017517090,
-49.9299926757813,24.6582145690918,
-40.2735557556152,1.35145783424377,
-23.4080619812012,-20.3357830047607,
-7.80797719955444,-17.4889163970947,
-0.168619185686111,-6.42818641662598,
-3.84843850135803,-15.5982360839844,
-9.93540573120117,-37.4970054626465,
-2.76371407508850,-37.8814735412598,
12.1797838211060,-11.4817256927490,
15.6957139968872,5.10808467864990,
7.30356693267822,-14.3320188522339,
7.22183418273926,-48.4218711853027,
22.5899620056152,-59.1731719970703,
31.2023868560791,-45.1289710998535,
8.31549072265625,-22.3926448822022,
-25.4830284118652,-0.667835354804993,
-20.1954116821289,18.5413551330566,
29.8934764862061,23.2391223907471,
67.6171798706055,8.18772983551025,
43.3495407104492,-6.58276605606079,
-6.39559030532837,6.14529037475586,
-13.2102184295654,33.0815734863281,
23.5534820556641,33.1801338195801,
34.2039222717285,-2.91984558105469,
-12.5365085601807,-29.5830383300781,
-57.8838615417481,-14.3498563766480,
-33.3927536010742,9.66789054870606,
34.0894660949707,-1.86941063404083,
58.3054351806641,-34.8439941406250,
14.0911865234375,-39.4715499877930,
-31.8311500549316,-11.3816432952881,
-28.3661842346191,5.94436168670654,
0.199078798294067,-8.94341278076172,
9.13582706451416,-18.6922283172607,
5.22352552413940,10.6797838211060,
18.3572521209717,52.2741470336914,
31.7813873291016,58.8466224670410,
12.9446735382080,33.4859466552734,
-19.6647186279297,19.3345985412598,
-16.0293006896973,29.1814785003662,
29.2367248535156,34.0762443542481,
56.2779502868652,16.0174255371094,
29.2263355255127,-6.20097255706787,
-8.75872707366943,-13.2662839889526,
0.612944662570953,-7.76606273651123,
42.4363288879395,3.49907779693604,
57.4693527221680,16.6195411682129,
33.2144660949707,21.1465225219727,
6.06393337249756,0.294925451278687,
2.02467083930969,-43.9162063598633,
13.3779468536377,-68.3881530761719,
28.9411163330078,-41.1818542480469,
48.0991401672363,9.60593795776367,
60.7253761291504,25.4030437469482,
39.9817390441895,-1.25357711315155,
-15.6006774902344,-24.2660923004150,
-60.0146636962891,-18.5845680236816,
-55.1379508972168,-8.40609836578369,
-20.0040283203125,-14.1753015518188,
0.437233597040176,-12.0369863510132,
3.06725668907166,22.1706905364990,
10.1118555068970,60.2244262695313,
21.3539237976074,49.4526443481445,
15.0171623229980,-9.58834743499756,
-1.65470719337463,-55.3615875244141,
2.31205654144287,-50.1257896423340,
34.3393859863281,-20.8852996826172,
52.7417602539063,-6.73800182342529,
27.4898910522461,-4.64527988433838,
-6.96668529510498,12.4939765930176,
1.08594155311584,36.5348014831543,
42.1227340698242,42.1309585571289,
60.9142951965332,28.7217330932617,
32.6026992797852,20.1477451324463,
-0.741552531719208,23.7308769226074,
0.325816512107849,17.8650646209717,
18.4260272979736,-4.95530652999878,
22.0685806274414,-16.2393169403076,
11.9847183227539,5.99308919906616,
12.6335411071777,38.1396522521973,
27.3260211944580,37.6032714843750,
30.4133071899414,2.79655599594116,
4.67829418182373,-27.5006046295166,
-27.8998699188232,-32.6932182312012,
-37.7440567016602,-21.4343452453613,
-19.8230304718018,-8.88377666473389,
3.19253444671631,2.74332308769226,
12.0055046081543,14.7694196701050,
-2.77473688125610,16.6180953979492,
-29.0019550323486,1.74746680259705,
-35.5567436218262,-18.6624584197998,
-3.71848630905151,-23.7103385925293,
38.3950881958008,-11.7702751159668,
44.5937461853027,3.07930898666382,
3.15265178680420,11.3963031768799,
-35.7755393981934,6.21245384216309,
-21.5709552764893,-18.9055843353272,
29.3269882202148,-55.6692314147949,
55.0950889587402,-66.4654388427734,
35.7108306884766,-28.5844402313232,
14.7141847610474,33.9916610717773,
29.2017631530762,66.8301849365234,
51.2796325683594,44.2580566406250,
41.0803070068359,1.60313749313355,
10.5657110214233,-17.4698867797852,
2.72633767127991,-14.6701488494873,
23.6277942657471,-15.3059778213501,
28.6538925170898,-20.0078430175781,
-7.61938524246216,-4.17402505874634,
-48.0418739318848,31.7715663909912,
-50.4762763977051,52.0571022033691,
-23.4362373352051,40.2600250244141,
-7.99545764923096,27.2120189666748,
-17.3346405029297,41.2166900634766,
-32.5862541198731,63.2160530090332,
-41.8012886047363,50.6013450622559,
-52.6810722351074,1.67131733894348,
-52.6787300109863,-37.8697204589844,
-22.0451622009277,-29.0084476470947,
29.2873954772949,9.64615058898926,
54.5447387695313,30.0015888214111,
30.1606884002686,15.2911748886108,
-11.4415454864502,-13.3070697784424,
-18.6243190765381,-26.6458759307861,
10.4086437225342,-11.5792179107666,
32.5542106628418,15.6292915344238,
26.6666278839111,23.0692367553711,
17.2874336242676,-6.51933479309082,
23.8128223419189,-49.4756584167481,
37.1092300415039,-57.3612937927246,
47.9460067749023,-14.0564737319946,
55.3525543212891,34.3113670349121,
55.2988090515137,33.7137718200684,
37.2176399230957,-10.7394943237305,
3.74311852455139,-40.3179931640625,
-10.4646062850952,-25.4420299530029,
9.81594562530518,-2.21712088584900,
27.4067649841309,-9.85625457763672,
1.66826593875885,-32.5669822692871,
-47.7573852539063,-26.2252559661865,
-58.8335685729981,10.1639986038208,
-22.0092067718506,31.5337505340576,
1.36274421215057,10.9560432434082,
-25.1376438140869,-21.9483184814453,
-53.7812385559082,-25.4684448242188,
-22.6457653045654,-0.180564224720001,
47.7908706665039,19.4250030517578,
71.1714630126953,11.0077247619629,
15.5742282867432,-10.1260690689087,
-51.4255752563477,-19.2850532531738,
-53.4197387695313,-11.0179748535156,
4.35993099212647,1.04519486427307,
50.8081665039063,1.53102385997772,
44.6824073791504,-12.6470451354980,
8.90946006774902,-30.2962265014648,
-17.3934383392334,-39.6673049926758,
-24.9987583160400,-37.1756134033203,
-22.3536815643311,-30.6184291839600,
-12.7622470855713,-23.3443889617920,
2.56359624862671,-12.0800170898438,
16.1638259887695,0.317915022373199,
12.4862899780273,6.99357175827026,
-7.46615028381348,-3.55645036697388,
-26.1646423339844,-27.9652519226074,
-25.1570491790772,-48.9432716369629,
-8.71873283386231,-52.2721214294434,
8.03795528411865,-34.9770507812500,
14.8332996368408,-6.27431917190552,
8.15354251861572,18.9408473968506,
-0.805319130420685,22.1569938659668,
-1.93192923069000,-1.25800776481628,
6.48557901382446,-31.8188571929932,
16.7253894805908,-34.5493545532227,
14.9038982391357,3.21095705032349,
-2.80968308448792,50.1459083557129,
-23.2497901916504,62.8210258483887,
-29.7432518005371,27.9552383422852,
-14.2074193954468,-23.1280212402344,
10.6849575042725,-50.1817588806152,
26.4747371673584,-41.5261077880859,
22.7681274414063,-13.8230228424072,
3.57004928588867,10.8409614562988,
-20.0176105499268,25.6943225860596,
-34.5331153869629,33.1600875854492,
-38.6295776367188,36.4997978210449,
-36.9330444335938,37.8651695251465,
-32.2700233459473,37.5720710754395,
-18.8918781280518,32.9601364135742,
0.189649581909180,21.2699794769287,
11.1206436157227,6.29581737518311,
0.456010818481445,-2.35079288482666,
-23.2649040222168,1.26427125930786,
-32.6818733215332,8.97393321990967,
-13.1667966842651,10.1826057434082,
13.9395532608032,-1.37208127975464,
19.6864204406738,-15.0481090545654,
12.4891891479492,-24.3739147186279,
19.1050472259522,-29.1210861206055,
40.7752456665039,-30.5836372375488,
45.3972663879395,-26.2638912200928,
18.6483192443848,-14.9452896118164,
-2.93814897537231,-6.70267581939697,
15.9056549072266,-9.38339042663574,
55.5089416503906,-19.4841880798340,
56.9029617309570,-14.2709426879883,
12.6294765472412,14.2068271636963,
-23.6851863861084,48.1752586364746,
-10.8517227172852,62.0394096374512,
23.5932769775391,50.0520973205566,
25.8029041290283,25.8563556671143,
-0.642369747161865,2.05726504325867,
-8.76263904571533,-20.5488414764404,
17.0602951049805,-40.0322341918945,
44.5219230651856,-49.6120262145996,
42.2767601013184,-44.4720726013184,
19.3613204956055,-29.9999561309814,
1.58010601997375,-11.9556541442871,
-9.40013885498047,15.9627380371094,
-24.7114467620850,50.9433288574219,
-43.5105247497559,67.4552917480469,
-50.2562675476074,44.8445968627930,
-41.5416793823242,-0.773340702056885,
-21.8198032379150,-28.4033260345459,
15.3343286514282,-18.1146430969238,
60.3797302246094,5.75390577316284,
75.6765213012695,17.0032520294189,
38.4996948242188,15.6097650527954,
-22.3557586669922,16.8626632690430,
-52.2755546569824,15.6183395385742,
-35.9757843017578,-4.47375774383545,
-10.5572175979614,-28.3028087615967,
-6.44581985473633,-22.8677577972412,
-9.67785930633545,10.0469589233398,
2.09206724166870,23.8304233551025,
7.14199829101563,-7.45084142684937,
-18.9262809753418,-48.1880187988281,
-44.9813880920410,-45.8780517578125,
-24.7261714935303,-1.30402588844299,
25.4330577850342,41.3717346191406,
40.6266365051270,49.8882408142090,
-2.29505348205566,36.5974006652832,
-49.5596084594727,16.8243732452393,
-47.4504737854004,-18.7460575103760,
-15.1224756240845,-62.3246688842773,
0.0672370120882988,-74.4378890991211,
-8.17715263366699,-36.6902732849121,
-9.46615791320801,10.5370903015137,
-2.06680369377136,16.8515186309814,
-14.6054553985596,-14.0019607543945,
-40.2307014465332,-34.7609901428223,
-32.4010276794434,-28.6183319091797,
19.5741271972656,-20.1206779479980,
60.1085205078125,-19.4993438720703,
45.5509757995606,-0.210921525955200,
5.84539747238159,45.6624374389648,
-4.30129671096802,71.4614639282227,
16.1581668853760,33.9814605712891,
24.4159622192383,-31.8652553558350,
0.373412609100342,-53.4305191040039,
-22.5433292388916,-18.8491230010986,
-12.2361555099487,5.73975038528442,
13.4809265136719,-21.8602924346924,
28.2720375061035,-63.1176567077637,
29.7262516021729,-58.5154571533203,
25.4950981140137,-1.98783469200134,
11.4148292541504,50.1898536682129,
-6.24350547790527,53.2483749389648,
-6.29524183273315,22.9921798706055,
18.4195976257324,-0.834423601627350,
32.4765319824219,-3.33915948867798,
6.06592416763306,5.44102382659912,
-33.1091270446777,1.27378797531128,
-32.6847991943359,-24.7763957977295,
10.7753200531006,-49.6321334838867,
36.6736602783203,-32.8091888427734,
7.68184947967529,26.4175701141357,
-38.0809822082520,73.4351730346680,
-43.6563911437988,56.5768699645996,
-17.4076766967773,-8.04017925262451,
-7.20922660827637,-44.5985221862793,
-21.9870986938477,-20.1070766448975,
-24.2520828247070,14.4143495559692,
11.3219442367554,-6.02739810943604,
52.3182182312012,-56.2788009643555,
56.9215164184570,-54.6119194030762,
25.1042003631592,13.8673353195190,
-8.36163902282715,69.8292770385742,
-19.8121566772461,48.4903144836426,
-13.6779966354370,-13.4439086914063,
-6.78442239761353,-32.9249725341797,
-7.00690031051636,8.21039295196533,
-20.1093063354492,45.0997467041016,
-41.7549285888672,28.2575550079346,
-48.7054481506348,-22.0733928680420,
-25.1149635314941,-56.4259605407715,
15.6447219848633,-56.7289772033691,
44.3403968811035,-37.9555282592773,
48.5000877380371,-12.0428028106689,
34.8446807861328,8.74831104278565,
11.8858680725098,3.55340766906738,
-15.3909521102905,-27.2160720825195,
-37.3441352844238,-44.0015373229981,
-36.2648353576660,-13.1861820220947,
-12.3973197937012,35.6243286132813,
-0.175408929586411,42.3487243652344,
-22.0792942047119,-5.30955648422241,
-51.2865562438965,-54.9882354736328,
-47.6277999877930,-58.0093612670898,
-13.0917167663574,-30.9856376647949,
13.0881776809692,-22.8590526580811,
16.1782493591309,-32.0573501586914,
23.1765384674072,-24.1269741058350,
49.1882133483887,7.84782457351685,
61.2135047912598,31.6799907684326,
23.7519836425781,22.3603763580322,
-35.0152206420898,0.355983704328537,
-49.7919120788574,-5.88233947753906,
-7.68157863616943,6.31737709045410,
36.9081268310547,18.4799976348877,
36.4129714965820,17.7751083374023,
9.98218536376953,7.27457141876221,
6.02327871322632,-2.78159832954407,
23.8561859130859,-3.76808667182922,
26.5040321350098,12.0216293334961,
5.12357473373413,42.7097206115723,
-5.60433673858643,60.9701347351074,
16.9576740264893,47.7890319824219,
46.8568000793457,21.3489017486572,
38.0275726318359,9.96802425384522,
-11.3163881301880,7.58585453033447,
-54.1906051635742,-9.22821331024170,
-51.9267539978027,-35.7083625793457,
-15.1249008178711,-35.0523872375488,
17.5190391540527,6.95471572875977,
16.8894462585449,43.0615196228027,
-10.6405973434448,24.5359649658203,
-31.8858089447022,-27.8277893066406,
-23.7064971923828,-48.8519973754883,
-0.958257734775543,-27.5516204833984,
5.64908504486084,-13.3927297592163,
-12.2163953781128,-35.8124580383301,
-25.9021072387695,-57.1684799194336,
-10.4587068557739,-34.3975486755371,
19.5729427337647,5.71502542495728,
19.8029861450195,5.94915914535523,
-17.7256889343262,-27.5657348632813,
-50.2880668640137,-38.5553359985352,
-38.8561325073242,-3.57806968688965,
2.99314832687378,32.2606735229492,
32.5001678466797,27.0380306243897,
32.8075752258301,5.95970726013184,
20.7241973876953,17.1890697479248,
11.2738800048828,49.6383934020996,
-1.61366319656372,46.8872642517090,
-20.8455543518066,-2.17044043540955,
-29.4540596008301,-46.3887481689453,
-16.1184082031250,-37.2008552551270,
-0.132749736309052,14.1133050918579,
-7.89579868316650,51.1079978942871,
-38.4061088562012,37.3455352783203,
-61.7666816711426,-10.4957809448242,
-59.7671852111816,-48.8448410034180,
-39.3893623352051,-47.0871124267578,
-10.8519392013550,-9.59891986846924,
23.5972976684570,25.6071510314941,
53.8518104553223,24.3146324157715,
57.4088554382324,-1.00210893154144,
26.9203338623047,-4.08584260940552,
-10.3989562988281,26.4727935791016,
-17.7955570220947,47.4079513549805,
5.67450618743897,16.0658016204834,
23.3136310577393,-38.7900428771973,
10.3387413024902,-54.5477561950684,
-19.0465660095215,-17.8145637512207,
-37.1425094604492,13.7444181442261,
-40.9233398437500,-11.4363937377930,
-40.6576423645020,-62.8874206542969,
-37.0088005065918,-71.5541076660156,
-22.8595657348633,-26.6541824340820,
0.554220795631409,19.8000679016113,
23.7496471405029,27.2171173095703,
34.0557670593262,10.0003261566162,
30.8517360687256,2.53856849670410,
11.7673540115356,11.6662464141846,
-20.1609153747559,25.8041381835938,
-46.5994758605957,37.7013092041016,
-45.4873085021973,42.2674179077148,
-20.6854972839355,26.7548961639404,
-1.70601367950439,-12.3197135925293,
-5.24871397018433,-51.9292793273926,
-10.2252483367920,-61.5475730895996,
0.928757905960083,-41.5745658874512,
12.8396844863892,-24.8557319641113,
-0.871658623218536,-21.1216964721680,
-30.8023700714111,-13.3515071868896,
-31.2765827178955,5.17656087875366,
11.0453910827637,12.7534685134888,
53.3470420837402,-2.38429427146912,
46.0685997009277,-18.2983932495117,
-4.38585853576660,-8.75375556945801,
-48.1671676635742,11.3215913772583,
-48.7890968322754,7.49114799499512,
-16.5418701171875,-18.6507072448730,
20.0235157012939,-29.8091030120850,
46.5146446228027,-10.6212749481201,
56.5663261413574,9.48388671875000,
45.3575820922852,3.94283890724182,
16.3925075531006,-6.66262149810791,
-12.0268745422363,13.8685951232910,
-18.0650367736816,51.4122276306152,
1.84158539772034,58.8610496520996,
24.5539894104004,17.8784751892090,
22.4218597412109,-33.3532028198242,
-3.25778222084045,-45.9089050292969,
-26.2453784942627,-17.4297428131104,
-24.5300865173340,13.2555656433105,
1.56469225883484,14.9931583404541,
24.2390480041504,-5.70248222351074,
17.9415626525879,-27.0424156188965,
-2.40831685066223,-34.0043754577637,
-3.72066140174866,-27.2716293334961,
22.4616622924805,-19.5847873687744,
45.2286415100098,-23.8193321228027,
26.9457721710205,-29.5891723632813,
-20.2545490264893,-17.2984199523926,
-52.0267982482910,15.4755401611328,
-44.6049118041992,38.0720977783203,
-30.6632022857666,19.9783401489258,
-41.9483070373535,-22.8399658203125,
-58.7074050903320,-45.0008277893066,
-32.8888931274414,-25.5548419952393,
30.9340076446533,-1.14118337631226,
68.0296096801758,-11.0529155731201,
36.1326560974121,-39.5858154296875,
-23.9122257232666,-42.0285758972168,
-36.5990028381348,-9.75436878204346,
9.52750968933106,13.9690246582031,
50.5395660400391,-6.68075466156006,
40.7664985656738,-50.3847198486328,
9.90767860412598,-68.9570236206055,
13.1495275497437,-43.4696540832520,
49.5870132446289,3.00385999679565,
65.9124603271484,36.4692764282227,
33.4257240295410,42.8431663513184,
-18.9265747070313,29.7336044311523,
-50.1533699035645,8.94913578033447,
-44.9020690917969,-11.5639400482178,
-19.7817192077637,-24.0159130096436,
7.31308174133301,-24.9170303344727,
19.7958164215088,-14.7954397201538,
7.16536617279053,2.67011785507202,
-21.1206245422363,17.5552577972412,
-39.8533515930176,16.7118568420410,
-32.9618835449219,1.35586929321289,
-20.1535415649414,-3.94279980659485,
-22.7314910888672,15.1125926971436,
-29.8539638519287,43.2631607055664,
-17.4465885162354,46.4899902343750,
7.14329242706299,13.7059335708618,
11.0671596527100,-23.3149890899658,
-11.5730161666870,-31.1778373718262,
-28.8197803497314,-16.3916740417480,
-10.7577056884766,-8.64640235900879,
20.3494358062744,-20.0102729797363,
20.1775093078613,-31.1533107757568,
-9.85842514038086,-28.9277744293213,
-30.6784992218018,-24.3431072235107,
-20.9398536682129,-25.1651344299316,
-2.94042778015137,-19.6677093505859,
-2.41448569297791,8.38886165618897,
-16.2519912719727,44.1294136047363,
-31.4137878417969,57.9957580566406,
-41.2634162902832,44.1640472412109,
-42.2003402709961,25.8155632019043,
-26.2162132263184,19.7019901275635,
4.05607223510742,16.9819259643555,
27.4058094024658,7.57114553451538,
27.4238967895508,5.96027803421021,
19.0978355407715,27.8839359283447,
28.4494857788086,52.2436485290527,
44.7053375244141,48.4657630920410,
33.7755050659180,19.4854221343994,
1.08751726150513,-1.61485707759857,
-9.20337009429932,7.58168745040894,
13.8163890838623,31.7545032501221,
27.6806983947754,40.5386466979981,
4.50501251220703,29.9218196868897,
-23.0108261108398,12.4865913391113,
-9.69474029541016,-4.69450044631958,
27.9424018859863,-18.9300746917725,
31.5576992034912,-18.8609867095947,
-1.05163669586182,-10.9859476089478,
-13.1753492355347,-19.5504455566406,
19.3484306335449,-47.6562309265137,
45.7455520629883,-56.0384216308594,
20.2506237030029,-10.6706466674805,
-23.2142257690430,54.1399459838867,
-30.4034671783447,63.2707481384277,
-9.35314846038818,5.02643108367920,
-8.01920890808106,-43.6197166442871,
-26.9590663909912,-18.0670814514160,
-22.5632991790772,37.4391937255859,
15.2126808166504,38.4411773681641,
34.2568855285645,-16.0460891723633,
2.81603264808655,-42.0652465820313,
-39.2156219482422,-0.814798474311829,
-36.3031845092773,43.8222770690918,
0.835066318511963,21.1722278594971,
20.1518268585205,-39.5084304809570,
13.1676998138428,-57.9097938537598,
8.10093021392822,-18.4548053741455,
13.1123390197754,15.0408992767334,
8.19489860534668,-2.53806710243225,
-5.87488031387329,-38.1448402404785,
-1.89725625514984,-34.7521629333496,
26.1994304656982,2.40712237358093,
41.2526512145996,17.3236408233643,
13.2659320831299,-12.1978816986084,
-30.4242458343506,-46.4323120117188,
-43.2817649841309,-40.7295417785645,
-27.1031074523926,0.394315719604492,
-18.2977313995361,32.3346900939941,
-19.3438549041748,19.8661155700684,
-0.0240173339843750,-19.7355556488037,
38.2411651611328,-34.3865852355957,
53.6835899353027,-6.66635894775391,
25.7508869171143,33.4228668212891,
-11.0066747665405,43.6854667663574,
-15.0711765289307,18.3848628997803,
5.95723962783814,-10.3245105743408,
11.6110467910767,-18.4881572723389,
-5.40209150314331,-10.8334350585938,
-16.1978092193604,-0.821316182613373,
-12.7542018890381,12.8681249618530,
-17.8295555114746,28.8180522918701,
-36.9393577575684,25.1937484741211,
-36.2221031188965,-6.86212873458862,
-0.212490558624268,-38.3979187011719,
35.3908271789551,-29.4297695159912,
35.9654731750488,16.4349842071533,
14.1667585372925,54.2640342712402,
9.76287460327148,55.0904502868652,
19.0266914367676,38.2675323486328,
3.85001373291016,29.3111610412598,
-42.2478294372559,21.1723060607910,
-67.6734542846680,-4.40773963928223,
-36.8822212219238,-32.3195495605469,
17.7398262023926,-23.1379165649414,
36.5345382690430,21.7467842102051,
9.71284008026123,54.9659004211426,
-23.3817138671875,40.0479011535645,
-36.2073593139648,-3.94225454330444,
-36.6753921508789,-33.0263824462891,
-34.6827354431152,-34.3279571533203,
-17.4499359130859,-34.2274055480957,
19.3756999969482,-42.3699035644531,
50.0888099670410,-38.4095916748047,
43.3710021972656,-8.36569023132324,
4.98210525512695,19.8688411712647,
-20.4898624420166,9.95877647399902,
-3.16812920570374,-25.0044250488281,
36.7077407836914,-33.8035736083984,
55.4595146179199,9.38975620269775,
38.9863395690918,61.8073501586914,
5.54341936111450,68.6584091186523,
-15.1817731857300,29.7173347473145,
-17.0642528533936,-6.99989748001099,
-20.1286144256592,-13.3068075180054,
-32.0787620544434,-7.78817319869995,
-34.0318222045898,-17.6785888671875,
-12.4010696411133,-36.2807807922363,
13.4908943176270,-43.2221870422363,
10.7946996688843,-43.1956062316895,
-17.8090419769287,-45.1666908264160,
-30.7207527160645,-42.6033210754395,
-4.60938930511475,-18.3607101440430,
29.3924121856689,17.7442131042480,
17.5218448638916,37.0645065307617,
-33.4433250427246,34.3947410583496,
-56.9932632446289,31.7965679168701,
-18.9106140136719,41.0463256835938,
35.6709327697754,42.5253982543945,
40.6832733154297,20.0656318664551,
-0.765074253082275,-6.39805746078491,
-23.7830104827881,-16.5042572021484,
6.00401115417481,-26.3990478515625,
49.6506233215332,-51.1005096435547,
53.3136024475098,-65.5764465332031,
23.9057369232178,-37.3707160949707,
0.0583782196044922,19.1459903717041,
-7.81193399429321,47.2509613037109,
-22.3905887603760,21.2561912536621,
-45.8918914794922,-18.1711196899414,
-42.7065086364746,-25.5549106597900,
-1.94549465179443,-7.97858905792236,
33.1866416931152,1.46516978740692,
19.0492973327637,2.41421294212341,
-24.5785636901855,3.14262580871582,
-41.3696098327637,-12.4441337585449,
-13.2539691925049,-54.6944427490234,
20.4980030059814,-82.8534545898438,
14.0368165969849,-46.8281593322754,
-22.7967510223389,33.7093467712402,
-45.1554565429688,72.5234146118164,
-31.1471061706543,30.0916595458984,
1.20852410793304,-31.5643634796143,
23.8051376342773,-41.1367378234863,
14.9136161804199,-13.5198822021484,
-20.4708557128906,-13.7772951126099,
-52.4146156311035,-42.9355506896973,
-54.2877006530762,-38.6917648315430,
-26.1775932312012,15.4163761138916,
0.634383201599121,51.7387123107910,
7.59625530242920,17.1887245178223,
10.6773881912231,-44.9069595336914,
31.3567314147949,-56.2563247680664,
52.7872543334961,-6.75069046020508,
37.2986145019531,44.5961494445801,
-4.49060297012329,53.1924858093262,
-19.4586734771729,34.8614158630371,
13.4699115753174,26.7822589874268,
39.7188796997070,32.2127876281738,
8.97258663177490,29.8187389373779,
-49.6629943847656,17.3078937530518,
-59.1797828674316,12.2196474075317,
-0.0224423408508301,19.9152030944824,
57.5132217407227,33.2800559997559,
51.3741760253906,34.6958312988281,
6.14749050140381,12.6056470870972,
-14.5136175155640,-23.9572486877441,
2.89868783950806,-41.8731346130371,
16.2102489471436,-18.4339675903320,
-0.875689268112183,27.1993274688721,
-28.8969287872314,56.5174140930176,
-45.4759216308594,47.0053863525391,
-56.1654624938965,21.9055442810059,
-62.5673217773438,9.63171672821045,
-49.0599861145020,-1.79582750797272,
-12.5175504684448,-34.5430908203125,
14.5624399185181,-71.6178207397461,
3.05169343948364,-64.5218505859375,
-30.8648872375488,-12.2274961471558,
-41.1189041137695,28.8906974792480,
-16.1102256774902,18.9629802703857,
3.61158919334412,-12.2258119583130,
-6.49092483520508,-11.7430610656738,
-25.7601203918457,15.2793712615967,
-32.4990768432617,13.4662017822266,
-28.3170986175537,-30.8591117858887,
-21.8301506042480,-67.5934295654297,
-11.6339368820190,-53.7832946777344,
5.81912899017334,-14.8311920166016,
17.6028842926025,-1.67108047008514,
10.6535158157349,-6.17287158966064,
6.96106815338135,7.46514225006104,
25.0353240966797,34.2394714355469,
49.2528305053711,31.9069824218750,
43.8920669555664,-10.6576538085938,
17.4883441925049,-42.2931556701660,
16.4805335998535,-27.0004653930664,
49.8291320800781,11.4313135147095,
61.6619796752930,26.0151195526123,
16.2174510955811,10.3664512634277,
-41.8817596435547,-5.25763416290283,
-40.8360443115234,-10.4830589294434,
17.6054859161377,-20.2581176757813,
61.0264053344727,-24.3908729553223,
37.7534179687500,3.21435523033142,
-20.6261024475098,49.4463882446289,
-55.7391624450684,61.5591506958008,
-51.8224372863770,17.1773109436035,
-34.4440917968750,-42.7081985473633,
-21.0553264617920,-62.6536674499512,
-14.3832511901855,-40.7820968627930,
-20.4282112121582,-20.7724971771240,
-41.5811347961426,-28.0093784332275,
-56.0135536193848,-46.8699455261231,
-44.0343780517578,-54.8300132751465,
-14.2410039901733,-50.7124061584473,
6.22762537002564,-31.5989837646484,
10.0464010238647,7.97381019592285,
14.1927146911621,48.6582565307617,
29.1472606658936,59.5038223266602,
37.5177383422852,40.5553359985352,
25.5413780212402,28.2444477081299,
16.3830585479736,42.2049903869629,
25.0044994354248,54.4497985839844,
27.1756172180176,31.2104969024658,
2.66638064384460,-14.4345817565918,
-25.2675800323486,-37.8245849609375,
-17.0936012268066,-26.1489715576172,
15.0777559280396,-18.8937892913818,
20.7817249298096,-34.4864006042481,
-11.8636302947998,-49.5593681335449,
-30.2519416809082,-41.3167495727539,
-1.08356702327728,-31.3559150695801,
34.4709014892578,-36.4259605407715,
18.6091403961182,-40.7936744689941,
-28.0200424194336,-18.7464466094971,
-32.7183456420898,11.9312410354614,
12.2088203430176,11.5787296295166,
39.9351882934570,-15.3234796524048,
12.3614444732666,-26.8452644348145,
-24.7278556823730,-10.8260650634766,
-17.7731971740723,-6.75070762634277,
15.1809301376343,-37.4613609313965,
19.5890445709229,-64.1885757446289,
-8.06101608276367,-49.0004539489746,
-20.9738616943359,-24.1783447265625,
-1.35112237930298,-36.0288925170898,
17.3352966308594,-66.5541229248047,
11.0005826950073,-49.9241371154785,
-1.87408769130707,18.3918132781982,
-3.81019306182861,64.8342056274414,
-15.8105096817017,35.4251022338867,
-45.5864448547363,-24.9327430725098,
-57.5870018005371,-39.8361206054688,
-22.1825904846191,-2.14042615890503,
28.0011463165283,25.2949085235596,
34.7996139526367,9.39977073669434,
-4.92027950286865,-16.7143554687500,
-37.2294082641602,-19.9022750854492,
-22.0032978057861,-13.6408729553223,
15.7441101074219,-22.6214809417725,
29.6297473907471,-40.2542533874512,
14.8718147277832,-43.6270828247070,
-6.94511175155640,-25.3564853668213,
-23.8885593414307,-8.33934497833252,
-34.1028785705566,-10.0818166732788,
-26.4674663543701,-26.6395072937012,
3.63499331474304,-39.5714302062988,
38.3786048889160,-34.8566627502441,
48.1723442077637,-8.75119400024414,
28.4290218353272,26.0069541931152,
3.10950565338135,39.3970451354981,
-13.8812656402588,16.5194530487061,
-25.0573844909668,-13.0806312561035,
-34.7762641906738,-6.47935390472412,
-28.5842094421387,30.7555274963379,
4.54113006591797,49.5507926940918,
40.6120567321777,19.1476287841797,
47.3275222778320,-30.7507934570313,
27.8552589416504,-43.6979293823242,
13.6310520172119,-8.59222793579102,
23.3916511535645,29.8789024353027,
43.0919151306152,31.4571571350098,
48.0978431701660,4.92508172988892,
32.0971984863281,-18.8780708312988,
9.22645282745361,-23.5541324615479,
-0.693877577781677,-10.1650562286377,
10.0416727066040,11.6627464294434,
30.9985275268555,22.8361282348633,
44.4583129882813,5.48260307312012,
30.3433189392090,-35.4544525146484,
-2.00500798225403,-56.3018112182617,
-14.8674230575562,-26.6664295196533,
6.66561698913574,28.0125560760498,
30.3704662322998,55.6265602111816,
16.8517665863037,41.4371223449707,
-17.8490543365479,26.3211708068848,
-22.6447525024414,41.5866813659668,
15.9650688171387,59.2998352050781,
43.1224555969238,46.4174537658691,
14.6466064453125,22.7957687377930,
-42.3273735046387,24.2109603881836,
-63.4695434570313,43.4055938720703,
-43.0057907104492,35.2040214538574,
-32.7565765380859,-15.7704305648804,
-52.6107788085938,-65.0830383300781,
-60.1242332458496,-71.2739028930664,
-21.3466987609863,-44.2401123046875,
34.7966842651367,-18.0039405822754,
49.5833740234375,0.827106177806854,
21.5151882171631,17.3387126922607,
-4.55415964126587,18.8665847778320,
-3.41728782653809,-9.03997611999512,
12.0080976486206,-37.5080871582031,
23.9854984283447,-22.4488754272461,
37.5881271362305,29.2669029235840,
48.0060958862305,58.1876144409180,
31.2213783264160,29.9676513671875,
-21.7177200317383,-22.9529991149902,
-67.4452590942383,-46.8019371032715,
-59.6358604431152,-35.0454521179199,
-12.6806030273438,-20.0588665008545,
14.0743675231934,-12.9358177185059,
-10.1526069641113,5.22357845306397,
-54.2705764770508,37.2171401977539,
-70.2516479492188,49.2102317810059,
-43.2035865783691,27.1843795776367,
-4.66355037689209,-5.13011169433594,
16.6166267395020,-18.4298477172852,
24.8400192260742,-19.3487415313721,
35.1551170349121,-25.8262023925781,
50.5723457336426,-33.6366806030273,
58.2833900451660,-29.9180412292480,
46.6317787170410,-18.9321060180664,
26.4488067626953,-23.5321769714355,
20.2765388488770,-45.3385314941406,
36.2130470275879,-49.3683013916016,
46.5397300720215,-16.3657722473145,
16.1769065856934,28.6851310729980,
-36.0898704528809,53.0895233154297,
-57.0364608764648,49.4066619873047,
-18.3071804046631,33.2240371704102,
42.9895362854004,15.1224203109741,
60.1837692260742,4.16930770874023,
19.5226058959961,10.0109281539917,
-20.9116058349609,26.9769058227539,
-19.6879234313965,28.6095104217529,
4.39685821533203,-6.78852367401123,
8.64839363098145,-52.1257858276367,
-4.72252416610718,-55.9572029113770,
-4.27240800857544,-9.30754375457764,
12.6960582733154,34.6766128540039,
2.33383393287659,30.9219093322754,
-46.5127525329590,-2.13421440124512,
-80.3609619140625,-17.9643249511719,
-47.8204498291016,-11.7865476608276,
19.9116878509522,-7.66295719146729,
44.9194030761719,-8.51338386535645,
2.52168512344360,6.42271041870117,
-41.7239723205566,38.1864433288574,
-22.3080768585205,50.4426574707031,
40.2259979248047,20.1612930297852,
70.7200775146484,-23.4759502410889,
44.1005554199219,-36.0966949462891,
1.37391340732574,-20.3492031097412,
-4.60749912261963,-5.80488586425781,
25.5996341705322,-0.487256646156311,
48.7506217956543,10.5853939056396,
34.9907455444336,20.8233489990234,
-3.25019335746765,10.6149835586548,
-25.9817047119141,-11.0400810241699,
-9.05080795288086,-13.4078197479248,
35.1180419921875,14.2926559448242,
67.9859313964844,41.9708442687988,
56.1678924560547,44.6914634704590,
14.1690273284912,44.3999328613281,
-16.4275302886963,61.5356750488281,
-22.6427459716797,68.4193878173828,
-28.5450458526611,25.7784214019775,
-49.0740394592285,-39.8545684814453,
-66.2938766479492,-57.3497734069824,
-55.3493041992188,-14.1230707168579,
-20.3801670074463,24.7211036682129,
5.35826969146729,11.2255783081055,
12.7454357147217,-18.0102081298828,
25.8728809356689,-3.09610962867737,
45.5023422241211,43.3066787719727,
43.2456321716309,55.5346908569336,
7.61604785919189,10.2910327911377,
-26.0375881195068,-42.8725395202637,
-18.2177219390869,-55.3877220153809,
18.6855850219727,-34.9410667419434,
38.0363731384277,-15.4199285507202,
31.3676872253418,0.178202614188194,
29.3223991394043,21.3608283996582,
44.0372734069824,37.7054100036621,
38.9653778076172,26.3995475769043,
-7.20150756835938,-4.18474006652832,
-51.4970664978027,-22.2948131561279,
-36.7188110351563,-13.2464084625244,
28.7129917144775,6.70412302017212,
70.1410369873047,12.5881204605103,
45.0285301208496,4.11578798294067,
-6.52617073059082,-1.90136981010437,
-20.3535423278809,5.41059970855713,
4.22179174423218,20.7147026062012,
21.2301616668701,33.5615882873535,
2.34660530090332,31.5719127655029,
-28.1392192840576,10.2731819152832,
-36.6788635253906,-17.8863048553467,
-30.0870800018311,-31.8075828552246,
-38.6247520446777,-21.9293441772461,
-61.5538063049316,0.606162071228027,
-66.1830596923828,14.8743629455566,
-35.3218612670898,14.6073360443115,
5.40801811218262,5.97664976119995,
15.7226686477661,1.76848983764648,
-11.9374494552612,7.70835304260254,
-38.5153617858887,17.1973972320557,
-21.8893623352051,20.2106704711914,
25.8975677490234,11.5601263046265,
58.5007438659668,-5.19541883468628,
46.5466575622559,-10.6431646347046,
10.9396514892578,10.1365165710449,
-6.78396415710449,41.1661720275879,
1.35705876350403,49.1645812988281,
5.63903522491455,19.9653320312500,
-13.3616781234741,-21.9311485290527,
-26.8576946258545,-43.3423614501953,
1.83134806156158,-40.5104713439941,
55.2310256958008,-34.8032569885254,
71.6735992431641,-32.6521072387695,
27.2458381652832,-15.6344165802002,
-33.6075286865234,16.8448791503906,
-48.5992126464844,29.8976879119873,
-12.2656517028809,-3.90962171554565,
25.8110523223877,-55.7548713684082,
31.6430091857910,-63.8491134643555,
20.3505058288574,-16.2948398590088,
8.19974613189697,29.5144042968750,
-12.1945047378540,20.6286182403564,
-38.5102272033691,-20.8830261230469,
-34.8834533691406,-32.2796287536621,
14.1813497543335,8.11437225341797,
59.9803047180176,58.4053840637207,
47.9899063110352,66.3565521240234,
-1.39966559410095,35.0488739013672,
-18.8889770507813,11.4276399612427,
12.8102350234985,20.0496520996094,
26.9958209991455,42.8608970642090,
-13.2514400482178,43.7665061950684,
-51.9952163696289,9.80591201782227,
-21.5944252014160,-30.3707370758057,
42.2369308471680,-39.0956077575684,
48.5355453491211,-15.0471467971802,
-7.00843572616577,1.00639975070953,
-41.5907974243164,-17.2713718414307,
-14.9778556823730,-45.0168914794922,
16.4288978576660,-39.2667884826660,
-2.76521944999695,3.92809581756592,
-31.4292297363281,33.5448226928711,
-10.0921993255615,12.4064855575562,
37.7699890136719,-23.1523704528809,
35.0947341918945,-17.9768142700195,
-26.0670471191406,17.4857788085938,
-67.7738952636719,21.3708477020264,
-43.7362785339356,-30.3353424072266,
-3.02455306053162,-77.9743881225586,
0.865327656269074,-60.9596138000488,
-15.2421302795410,1.62123680114746,
-11.4667072296143,36.2248611450195,
3.02633333206177,20.2881145477295,
-4.90433979034424,1.47258996963501,
-33.2059669494629,23.0595436096191,
-50.4576950073242,56.5477828979492,
-45.5724372863770,47.9929771423340,
-44.0822715759277,-5.58071041107178,
-53.6276588439941,-55.5023689270020,
-52.6538238525391,-63.3262901306152,
-32.0317420959473,-36.8402404785156,
-18.0565261840820,-2.82540583610535,
-17.9478206634522,19.8245468139648,
-4.64935016632080,21.0943889617920,
32.4942398071289,2.62100458145142,
53.3543586730957,-19.4229106903076,
28.6110706329346,-22.3565483093262,
-13.9776096343994,-10.5813150405884,
-19.1351623535156,-14.4262208938599,
13.9232463836670,-50.9987068176270,
31.3231735229492,-80.5025711059570,
2.52687287330627,-57.2858619689941,
-38.2891540527344,6.33757019042969,
-45.1050109863281,49.3028526306152,
-27.7342262268066,44.2555503845215,
-28.2093601226807,17.6223793029785,
-56.1333694458008,5.25468444824219,
-75.3456420898438,3.83649301528931,
-58.3061294555664,-6.68679618835449,
-12.6606273651123,-12.8963613510132,
29.2711105346680,9.11341762542725,
47.5648002624512,43.5285720825195,
43.3096122741699,45.1672782897949,
30.8857707977295,11.6554517745972,
24.8971405029297,-7.17832136154175,
21.3087387084961,18.2381172180176,
12.1844196319580,54.4885139465332,
-4.44909954071045,58.0088691711426,
-15.8675508499146,37.3864097595215,
-3.32590866088867,31.2386398315430,
26.2113189697266,40.3561477661133,
39.7213211059570,38.6169242858887,
22.5494880676270,19.1939888000488,
-5.75986480712891,12.7610530853271,
-21.6725158691406,20.2111740112305,
-24.9130725860596,5.43984651565552,
-21.2071170806885,-41.0566368103027,
-7.04351425170898,-65.9467468261719,
24.8657760620117,-27.6585464477539,
49.4572944641113,33.7306175231934,
27.9707660675049,44.4772872924805,
-30.0178375244141,0.936945438385010,
-63.0276336669922,-34.6189689636231,
-27.6039276123047,-22.8842163085938,
37.1318588256836,4.89176702499390,
57.2426567077637,8.70741653442383,
20.3478584289551,2.51275658607483,
-12.3686256408691,20.6018447875977,
6.88278579711914,53.1994018554688,
47.5472526550293,59.8876152038574,
54.4182357788086,37.0987243652344,
16.9915218353272,19.2454090118408,
-21.9796886444092,26.0736122131348,
-30.5225067138672,33.5798072814941,
-25.6169033050537,22.1836051940918,
-28.1761970520020,0.598291158676148,
-36.8040733337402,-13.7055721282959,
-34.0297317504883,-15.4867868423462,
-15.6820535659790,-15.7960376739502,
1.19071137905121,-14.9442167282105,
8.08949375152588,-2.74428153038025,
8.54684448242188,17.4196968078613,
6.45823049545288,30.2993259429932,
6.97320175170898,30.2637310028076,
16.8858985900879,21.0394783020020,
36.2087020874023,7.28379964828491,
54.0627746582031,-3.25685024261475,
47.9573097229004,8.40152168273926,
4.33817243576050,47.6515960693359,
-57.0576782226563,83.7805328369141,
-93.7572402954102,69.7012557983398,
-76.2343444824219,1.00385725498199,
-18.6361236572266,-63.9816894531250,
28.1004943847656,-60.2055282592773,
27.6227111816406,5.85187673568726,
-9.98563194274902,64.1570281982422,
-36.6834983825684,60.9786148071289,
-27.9480094909668,15.9176893234253,
-3.88070964813232,-13.8547487258911,
3.32164192199707,-4.78243446350098,
-10.1600341796875,18.0604076385498,
-20.3110980987549,22.0377082824707,
-15.9298858642578,2.44546985626221,
-9.02842521667481,-18.9436416625977,
-10.8306875228882,-26.5410575866699,
-13.1127138137817,-24.9011058807373,
-1.21337842941284,-20.7714595794678,
15.8360424041748,-14.2308101654053,
8.97704029083252,2.60435056686401,
-24.2870368957520,23.9017524719238,
-58.8694496154785,32.5336685180664,
-66.0408401489258,16.8306064605713,
-45.1814880371094,-18.1667671203613,
-23.4340305328369,-39.5620002746582,
-17.0390682220459,-24.3748741149902,
-18.4745330810547,7.41694641113281,
-18.4054584503174,20.1047954559326,
-19.3208274841309,-1.11971652507782,
-25.3415145874023,-25.4454669952393,
-28.6421642303467,-16.3124637603760,
-17.1359996795654,20.1345100402832,
-2.23228335380554,42.4919090270996,
-5.70224761962891,30.4718189239502,
-29.3271846771240,2.83336544036865,
-40.4912414550781,-11.6377305984497,
-11.1645202636719,-15.3614387512207,
37.4886398315430,-30.3021316528320,
60.7689552307129,-56.3961715698242,
43.2133331298828,-67.3431930541992,
10.7478399276733,-51.0341949462891,
-0.251823902130127,-27.9810771942139,
5.73310232162476,-25.9497680664063,
6.31596517562866,-45.7680969238281,
-6.11777830123901,-58.0395317077637,
-18.9108028411865,-40.1842002868652,
-27.0871696472168,-5.51231622695923,
-35.6702270507813,14.1082353591919,
-48.1365013122559,1.34490609169006,
-49.8370552062988,-27.2783546447754,
-26.2384414672852,-35.2579421997070,
15.3114032745361,-2.86524009704590,
48.7329788208008,37.1395530700684,
46.3078155517578,29.9752044677734,
7.24609851837158,-27.5662384033203,
-42.0634689331055,-74.0855026245117,
-63.4431953430176,-50.4411849975586,
-37.9990692138672,17.2931671142578,
8.34236812591553,48.5118408203125,
35.2279968261719,5.24798774719238,
27.4410076141357,-44.8630714416504,
12.3157339096069,-29.5262565612793,
17.8318939208984,30.4051837921143,
38.1392517089844,48.1267204284668,
43.0193977355957,6.50122451782227,
18.1703300476074,-26.0357475280762,
-16.3803005218506,-2.92348289489746,
-35.9064941406250,28.1732196807861,
-35.5925598144531,2.95884943008423,
-28.8997020721436,-52.8706893920898,
-24.4902896881104,-60.7675094604492,
-20.9146804809570,-12.1199474334717,
-8.32938766479492,14.1280574798584,
14.4763088226318,-25.0267124176025,
34.9525680541992,-76.6837387084961,
38.7360191345215,-66.8692855834961,
17.9779567718506,-4.59246158599854,
-12.5002880096436,43.2851638793945,
-28.2807273864746,50.9409141540527,
-22.6610412597656,43.3367156982422,
-7.73434686660767,36.6668624877930,
3.19653129577637,18.7615737915039,
11.0926685333252,-5.90938282012939,
17.9299030303955,-9.35217571258545,
22.9224109649658,16.8568592071533,
19.7795848846436,29.5133895874023,
12.7221612930298,-5.94382762908936,
9.51856899261475,-61.3835258483887,
7.92109918594360,-74.6711730957031,
-3.16095352172852,-33.4164733886719,
-16.7073993682861,14.2365989685059,
-15.7266931533813,28.7604732513428,
-0.422637104988098,20.9446716308594,
9.01948833465576,15.8559198379517,
-3.87461137771606,19.7993335723877,
-22.2176456451416,15.2510976791382,
-19.6379470825195,-6.41716670989990,
-0.268243432044983,-27.0893383026123,
2.11147856712341,-31.5525360107422,
-26.0805892944336,-27.4086990356445,
-50.8131027221680,-32.2645874023438,
-34.0968971252441,-48.4430122375488,
5.64121770858765,-57.0795745849609,
15.7707872390747,-34.2314491271973,
-19.4858093261719,17.7089080810547,
-50.6078681945801,60.8644371032715,
-29.6633453369141,46.0628890991211,
22.1329593658447,-14.8805122375488,
41.1134567260742,-55.3807449340820,
14.8441696166992,-28.3608512878418,
-3.18688511848450,35.7757873535156,
21.8707866668701,66.4864578247070,
54.3717727661133,43.3482704162598,
42.7579269409180,17.0850830078125,
0.0253698825836182,32.5651016235352,
-23.1042041778564,60.8337326049805,
-13.8315792083740,52.1249465942383,
-9.59399700164795,11.7046613693237,
-27.1380577087402,-14.2004537582397,
-37.1106491088867,-19.1331157684326,
-20.8606548309326,-37.9692649841309,
-7.48784685134888,-71.1277618408203,
-22.3480758666992,-70.9077148437500,
-41.0088272094727,-17.5714721679688,
-24.1072139739990,30.8751945495605,
14.5110082626343,13.6336917877197,
32.4894447326660,-41.2483711242676,
29.5373172760010,-52.4221725463867,
36.1007194519043,0.402995824813843,
51.4048881530762,50.2174720764160,
34.8929138183594,41.7920265197754,
-20.6435890197754,1.26282024383545,
-66.1125335693359,-26.4264755249023,
-54.9433097839356,-39.6191825866699,
-15.1677360534668,-57.2394828796387,
-6.29250621795654,-61.6337547302246,
-32.7130851745606,-32.4417419433594,
-48.6495399475098,5.07870149612427,
-32.4816360473633,0.686846494674683,
-11.6142139434814,-42.2702217102051,
-5.91641759872437,-63.0910453796387,
-1.58400869369507,-24.5066261291504,
10.7486867904663,28.9567394256592,
18.7671604156494,33.2729225158691,
12.2291908264160,-6.53368568420410,
5.65583419799805,-30.7711277008057,
18.7526111602783,-12.7125511169434,
33.0158920288086,23.9486999511719,
21.6942844390869,44.5687522888184,
-8.70879268646240,37.2657737731934,
-23.0924663543701,12.1047840118408,
-10.1036005020142,-12.9030542373657,
0.0134416595101357,-25.5041770935059,
-4.69907140731812,-18.8737812042236,
-3.49533867835999,-6.60949707031250,
10.7944087982178,-6.48837757110596,
13.3020381927490,-14.4784173965454,
-11.5976133346558,-8.25820350646973,
-38.3727760314941,14.2675113677979,
-26.7687339782715,16.4679050445557,
16.2481250762939,-17.8002223968506,
48.3973999023438,-50.9598121643066};
