shortreal out[16384] =
'{0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
-4.36648497270653e-06,
-0.000747180718462914,
5.23935086675920e-05,
-0.00178522011265159,
0.000276090431725606,
-0.00315736024640501,
0.00100479775574058,
-0.000899338629096746,
0.00277266860939562,
0.00704684760421515,
0.00541969249024987,
0.0237905196845531,
0.00902761239558458,
0.0529022961854935,
0.0128122316673398,
0.0992690101265907,
0.0211915671825409,
0.0915164351463318,
0.00204224651679397,
0.119120717048645,
-0.0186217594891787,
0.140451192855835,
-0.125730335712433,
0.150780171155930,
0.0127733349800110,
0.219489634037018,
-0.0655424594879150,
0.0131699889898300,
0.0569725930690765,
-0.477253139019012,
0.202010393142700,
-1.14943146705627,
0.250376790761948,
-0.994743764400482,
0.133997678756714,
-1.49767589569092,
-0.196828484535217,
-2.11689448356628,
-0.911162853240967,
-4.30467176437378,
-1.23879337310791,
31.2400722503662,
-3.54356336593628,
-26.1557102203369,
-7.79165840148926,
1.22459912300110,
17.6930999755859,
15.2593269348145,
52.8402404785156,
37.2271842956543,
-11.4445581436157,
3.96658182144165,
3.53592967987061,
-9.58977127075195,
-9.77703952789307,
-50.0300865173340,
5.11400699615479,
64.0068511962891,
-40.0134963989258,
-11.7667703628540,
10.0384483337402,
6.50500869750977,
9.17521381378174,
-10.0754299163818,
36.2389678955078,
-23.0716400146484,
28.3180694580078,
17.0692539215088,
-48.0458641052246,
-11.1223602294922,
-6.67004108428955,
-10.8243083953857,
-48.2845764160156,
45.9763488769531,
35.5136833190918,
-28.4864177703857,
44.4487190246582,
35.4106903076172,
-18.5612297058105,
-50.5984878540039,
-2.74568557739258,
-13.6671037673950,
-10.5406513214111,
40.8392105102539,
-39.6200866699219,
-26.2053470611572,
9.42117500305176,
-31.4042892456055,
-0.386880874633789,
22.9769401550293,
-20.1259460449219,
4.42750549316406,
54.0993003845215,
25.1013031005859,
45.4781112670898,
53.6026306152344,
59.4080123901367,
37.6259956359863,
-23.0044612884522,
-12.4784173965454,
10.0456151962280,
19.3202037811279,
19.5989513397217,
69.2128067016602,
-8.82177734375000,
9.25082111358643,
58.4806022644043,
-55.6166229248047,
14.2877712249756,
32.2141075134277,
33.5107154846191,
16.1133422851563,
-15.5691289901733,
52.6962547302246,
-13.2556877136230,
-45.3768844604492,
-7.76243305206299,
6.89634561538696,
57.0280380249023,
10.8147926330566,
-40.7040863037109,
34.2829322814941,
17.5894107818604,
-27.7612648010254,
2.10851764678955,
36.5171928405762,
29.6674766540527,
-18.1586894989014,
35.3764495849609,
-7.35634422302246,
-19.1063499450684,
50.9577941894531,
-24.7376060485840,
34.5031089782715,
28.7340888977051,
-35.3985290527344,
9.96474456787109,
-33.6677436828613,
-3.46980094909668,
69.7668533325195,
2.74073576927185,
8.62287330627441,
26.5207366943359,
-37.0269508361816,
20.6266345977783,
32.6397781372070,
30.7916488647461,
31.8266468048096,
-9.50194835662842,
11.6434497833252,
-6.33880186080933,
25.9981956481934,
40.0197143554688,
-42.7410774230957,
40.8537979125977,
34.9554748535156,
-16.6180400848389,
52.6161804199219,
-28.3701972961426,
-9.96270370483398,
14.4374628067017,
-43.0025787353516,
-11.2655963897705,
77.9197921752930,
2.69919967651367,
-27.5453758239746,
69.5471725463867,
2.34175729751587,
33.3479499816895,
7.92644023895264,
-10.0538854598999,
54.1327438354492,
49.3649253845215,
-9.10667419433594,
0.553097963333130,
23.9000625610352,
-49.7763290405273,
-23.8864059448242,
11.2395191192627,
34.5446701049805,
14.1101760864258,
21.9295082092285,
-5.70205354690552,
8.75474929809570,
14.8303689956665,
-33.3999404907227,
20.8965435028076,
-19.1962184906006,
-5.70614385604858,
-5.16263341903687,
26.9686584472656,
49.9360961914063,
-6.80894184112549,
61.5069885253906,
-5.33454322814941,
-18.1610908508301,
95.3027267456055,
-0.988546848297119,
-33.0551147460938,
-7.17101430892944,
3.06470108032227,
55.5128593444824,
22.0493774414063,
32.0901489257813,
42.3924789428711,
-5.57402610778809,
-53.9039611816406,
29.2379837036133,
12.7760038375855,
-33.4739913940430,
70.1904373168945,
7.53231000900269,
-15.9694938659668,
10.2047090530396,
1.91303420066834,
14.2189054489136,
12.4335460662842,
36.5745239257813,
51.8352050781250,
-2.83018374443054,
22.3332843780518,
38.5922012329102,
-50.8824577331543,
33.8174362182617,
58.9347229003906,
13.9308738708496,
-7.56905746459961,
-32.6379089355469,
50.9085693359375,
-5.31897544860840,
-60.5835304260254,
28.1854553222656,
52.2372627258301,
3.06904053688049,
23.1700210571289,
-28.2376556396484,
-25.5243053436279,
64.0157470703125,
-52.8022804260254,
43.8390426635742,
38.8378219604492,
-7.95340061187744,
36.9797134399414,
-46.9399795532227,
24.3409137725830,
1.88263821601868,
44.1051216125488,
5.93641471862793,
-7.97888851165772,
52.6567344665527,
-23.2779216766357,
-15.7320356369019,
-20.9294223785400,
36.2117156982422,
39.7686271667481,
1.23998689651489,
-7.96164512634277,
-5.87530899047852,
27.3634166717529,
29.0579605102539,
9.88562583923340,
-40.6915512084961,
8.63047409057617,
13.8013057708740,
-51.9633712768555,
-7.19797515869141,
33.3328819274902,
21.9221305847168,
11.4901924133301,
51.9305114746094,
-0.905254364013672,
-27.8309516906738,
53.1786422729492,
14.5083036422730,
12.1202497482300,
31.8629341125488,
-40.8554878234863,
20.8463134765625,
45.8774833679199,
-47.7182960510254,
15.0313739776611,
35.9676361083984,
2.72911834716797,
-14.8326120376587,
-38.2085647583008,
-9.28870582580566,
-25.0940780639648,
-25.5199356079102,
22.9000320434570,
5.81539916992188,
-47.5068969726563,
29.4747314453125,
-15.5700340270996,
-56.5953216552734,
78.2079620361328,
20.4092063903809,
13.8852043151855,
-11.2901077270508,
2.02415752410889,
42.2248153686523,
-48.0538330078125,
63.2717323303223,
35.9720726013184,
-39.6885452270508,
9.59564018249512,
8.63940906524658,
-32.3345565795898,
-13.8495254516602,
21.7789707183838,
34.9500274658203,
33.9155158996582,
9.52370834350586,
38.0561180114746,
-22.3283176422119,
28.1079082489014,
10.7839803695679,
-22.5873756408691,
41.8044738769531,
26.9525108337402,
54.6135864257813,
-4.97745513916016,
2.84913420677185,
67.5051879882813,
24.0971622467041,
-21.8976058959961,
26.2237663269043,
-12.7868785858154,
-29.8806495666504,
60.7927970886231,
-23.5096950531006,
-25.3418560028076,
-16.7422084808350,
-3.56266188621521,
45.1649475097656,
-11.2102479934692,
9.63737010955811,
-31.5471973419189,
16.4455680847168,
20.3996295928955,
13.6805706024170,
65.3045654296875,
-51.9049758911133,
47.0212135314941,
40.4404220581055,
1.40559375286102,
27.9350261688232,
-44.3829650878906,
39.0394973754883,
-16.9465179443359,
19.4083728790283,
38.6163330078125,
-63.1704750061035,
-15.8239498138428,
27.2696723937988,
34.4184646606445,
-59.1428604125977,
-29.0026245117188,
-7.65918684005737,
-32.1021156311035,
22.3302459716797,
12.7433300018311,
-5.69897890090942,
3.83952236175537,
69.8979415893555,
-4.27690362930298,
-29.4062194824219,
41.6185913085938,
-0.892475128173828,
-8.75788402557373,
-13.9065332412720,
23.8167648315430,
45.4065856933594,
20.8610076904297,
-18.0559158325195,
14.9132843017578,
12.9760112762451,
-44.7619438171387,
70.5763092041016,
33.9339065551758,
-17.4320869445801,
24.5437297821045,
-17.0280914306641,
26.9696025848389,
15.3426570892334,
-61.3990097045898,
10.2591419219971,
2.48091030120850,
-44.1910667419434,
54.5015068054199,
2.54540443420410,
3.62370133399963,
-5.76203346252441,
-50.7644920349121,
37.8727226257324,
-27.1260528564453,
29.3218574523926,
9.27345085144043,
-35.9841423034668,
39.0630531311035,
-29.0526199340820,
45.7288208007813,
40.3839645385742,
-7.02909994125366,
5.54653167724609,
24.9895572662354,
46.2275390625000,
7.02409696578980,
38.6816787719727,
14.0787773132324,
-34.2175788879395,
14.9143142700195,
33.6453056335449,
-51.8049125671387,
-3.77425956726074,
-8.06125068664551,
-66.0393905639648,
10.7830572128296,
11.5929841995239,
-22.8739280700684,
21.0065193176270,
36.5568275451660,
-54.6902809143066,
-12.1895675659180,
49.2876892089844,
10.4903736114502,
29.6695671081543,
61.9583282470703,
12.8135433197021,
-14.6482410430908,
94.0389480590820,
14.7629432678223,
-25.8689785003662,
51.4437332153320,
-38.1559753417969,
-10.6137123107910,
8.97843647003174,
-3.52537488937378,
15.5552701950073,
-8.58090877532959,
6.06710004806519,
54.9063262939453,
0.840554237365723,
-18.3951263427734,
68.5332336425781,
-52.4331436157227,
-19.7965621948242,
79.6773529052734,
18.2178726196289,
-11.9622697830200,
-30.8367214202881,
-23.8521575927734,
-9.63116359710693,
73.3603286743164,
6.80529880523682,
-46.1434288024902,
47.2094039916992,
36.4206771850586,
-6.11949443817139,
-5.60782909393311,
49.4771804809570,
-14.1874809265137,
-11.1069297790527,
52.3636245727539,
-42.1893882751465,
31.8191699981689,
41.4301033020020,
-46.4650955200195,
-26.5954246520996,
-15.3128118515015,
39.0356788635254,
16.8183078765869,
38.0760917663574,
30.3154850006104,
-5.81820201873779,
50.8968353271484,
-24.7120933532715,
-4.66591739654541,
4.14768981933594,
-48.5884857177734,
12.0973625183105,
-26.0858230590820,
-37.1806144714356,
22.0940742492676,
34.3928756713867,
2.75750517845154,
14.4601755142212,
2.02506256103516,
-39.5502014160156,
-11.5595312118530,
40.8590965270996,
23.1320075988770,
-56.3849182128906,
25.9168834686279,
7.43653821945190,
9.83763408660889,
51.7549858093262,
-23.5472240447998,
30.9356155395508,
-2.66043186187744,
20.7977294921875,
45.9745941162109,
-7.05313491821289,
-21.3472328186035,
6.20927000045776,
17.8253593444824,
-28.2619838714600,
26.1166801452637,
-43.3319854736328,
-29.1065845489502,
54.3107185363770,
-10.5349302291870,
45.6708488464356,
13.6142501831055,
-40.1735458374023,
20.9125480651855,
-35.7438468933106,
-9.64843654632568,
5.44032716751099,
9.17816162109375,
49.8381690979004,
35.7371368408203,
53.4957046508789,
-15.8221435546875,
-13.1292715072632,
-24.9170780181885,
19.9780273437500,
35.0059127807617,
11.1314668655396,
53.9194145202637,
-14.9473352432251,
13.2138519287109,
5.52731800079346,
-30.0658302307129,
13.2152862548828,
-0.0473270416259766,
-62.0838165283203,
40.0271072387695,
11.4410190582275,
-30.3330135345459,
27.3408565521240,
-46.3378562927246,
8.26622962951660,
-18.8620910644531,
8.62357139587402,
48.3174514770508,
32.1018714904785,
29.0353584289551,
11.6745729446411,
54.6754798889160,
25.1094989776611,
34.9193191528320,
43.6295852661133,
-0.918533325195313,
-33.7426223754883,
-7.08774328231812,
-6.33222484588623,
-33.1882438659668,
-31.0943374633789,
-21.8723545074463,
-0.357658147811890,
-9.49373912811279,
-43.1649856567383,
1.77206230163574,
9.33415603637695,
6.63983345031738,
52.9506874084473,
-7.40110874176025,
37.2197113037109,
23.5681114196777,
23.3157196044922,
53.9344558715820,
1.83393001556396,
32.6468391418457,
47.5221138000488,
-7.18850708007813,
-25.1178627014160,
69.3527526855469,
10.5827579498291,
1.89696168899536,
16.6282558441162,
14.7796230316162,
22.3919639587402,
-21.0985546112061,
-1.82866644859314,
-33.0518760681152,
18.1375541687012,
-26.3558425903320,
-47.4236679077148,
4.38449192047119,
-11.3306188583374,
38.6986389160156,
-3.80652451515198,
-25.5520305633545,
68.8427505493164,
-3.01611804962158,
-35.1626892089844,
55.2419662475586,
-36.8586997985840,
-3.67088699340820,
58.2903213500977,
-8.45603084564209,
35.9408950805664,
13.8370332717896,
-21.3978939056397,
18.7901401519775,
26.1826038360596,
-11.4369621276855,
-29.2973346710205,
49.9040451049805,
18.8396778106689,
-30.7874145507813,
21.0890350341797,
18.5381679534912,
1.90547978878021,
-13.0257167816162,
48.3281211853027,
41.5191421508789,
37.9492454528809,
19.7507324218750,
-34.0772361755371,
32.0829315185547,
-15.6859312057495,
17.8156051635742,
38.8906326293945,
30.0056304931641,
13.1620903015137,
-12.4063644409180,
18.8432254791260,
-14.8403778076172,
39.9925956726074,
-14.1493911743164,
-32.7611885070801,
36.2247734069824,
19.4686737060547,
-35.3564605712891,
3.06590557098389,
43.2786445617676,
-6.32194137573242,
-0.740796566009522,
41.5374488830566,
21.3616237640381,
-41.2843475341797,
40.7318229675293,
10.0115280151367,
-16.4469261169434,
-9.19379615783691,
-17.2648086547852,
40.3293113708496,
16.4341697692871,
18.4207420349121,
-33.4156455993652,
34.5408668518066,
20.0081863403320,
-46.8864212036133,
30.1330490112305,
-31.2721710205078,
22.5358791351318,
23.9910030364990,
-41.3722190856934,
4.85309505462647,
27.9961605072022,
-3.89628791809082,
-39.9112167358398,
-24.7949867248535,
3.18325138092041,
11.3265743255615,
-57.2811203002930,
55.6156082153320,
6.34612464904785,
-24.3764114379883,
52.5581588745117,
-58.5079536437988,
12.3803329467773,
45.7016906738281,
-10.7651643753052,
-42.6195449829102,
52.7515716552734,
16.4283905029297,
-26.0732688903809,
10.6052513122559,
10.9420166015625,
33.1974449157715,
-26.2626838684082,
47.6246871948242,
-9.42806816101074,
-28.6917171478272,
22.4917602539063,
20.4540405273438,
42.1882247924805,
21.9935874938965,
22.7304325103760,
-45.1766242980957,
-13.3742437362671,
-4.40610122680664,
-7.87785434722900,
57.8058013916016,
30.8305664062500,
39.7186012268066,
12.0077266693115,
-0.742441773414612,
23.8506584167480,
-21.2610702514648,
-21.5673904418945,
-6.71121311187744,
5.04406118392944,
-7.88709306716919,
4.57534599304199,
51.9559745788574,
-0.335676193237305,
8.94919872283936,
60.2667541503906,
16.4574432373047,
-14.1145925521851,
-40.1948432922363,
8.66853713989258,
38.1824150085449,
-43.7177238464356,
39.0014190673828,
65.1630401611328,
-41.1346817016602,
41.6620063781738,
71.5950851440430,
-13.2053079605103,
-11.3554458618164,
8.95094394683838,
47.1553573608398,
43.6420593261719,
-44.8471183776856,
-17.6247901916504,
37.0303306579590,
-31.6028881072998,
-42.3185729980469,
-6.86293220520020,
-25.8726348876953,
-47.2460632324219,
-23.3542156219482,
-9.43541717529297,
-6.00687789916992,
16.3075790405273,
-15.1655244827271,
11.2505683898926,
-27.2157917022705,
-47.5473480224609,
67.8562698364258,
-4.10039234161377,
17.4565238952637,
16.4301700592041,
-11.9960632324219,
43.3217887878418,
-36.0435752868652,
7.12529754638672,
24.2705192565918,
1.38529324531555,
-26.6757373809814,
18.2695503234863,
32.7756042480469,
-20.9415531158447,
32.8861465454102,
18.0996990203857,
51.8171615600586,
29.9613227844238,
-3.14899539947510,
28.7186126708984,
46.5835342407227,
59.7047271728516,
7.94584369659424,
10.6566848754883,
26.9040985107422,
-7.68598747253418,
-3.13343334197998,
34.7156410217285,
-7.59805107116699,
-52.0607872009277,
-1.31379795074463,
-13.8403997421265,
-30.6142616271973,
5.80897045135498,
28.6812858581543,
44.3685798645020,
28.2476387023926,
15.5535850524902,
-23.3934097290039,
13.0561876296997,
-5.44197177886963,
-40.3500900268555,
34.5400238037109,
25.1255912780762,
42.9628562927246,
36.4072265625000,
41.3400611877441,
15.8037862777710,
27.3582458496094,
21.3088722229004,
-35.9282684326172,
45.2480278015137,
6.14863109588623,
3.87193202972412,
48.4440879821777,
52.0700912475586,
-23.7888450622559,
-10.8061876296997,
17.8070430755615,
-31.2572593688965,
63.5139579772949,
6.00113677978516,
8.19279575347900,
-17.0633926391602,
-30.6680450439453,
8.90075302124023,
-21.9092121124268,
72.3594055175781,
-31.6794509887695,
-11.9666023254395,
54.6225852966309,
-35.6992683410645,
68.0995025634766,
38.6914215087891,
-17.3773231506348,
20.9377307891846,
13.0766935348511,
42.4122238159180,
37.2946128845215,
7.10736656188965,
28.3834381103516,
46.3808441162109,
31.7327613830566,
33.1244316101074,
0.470155715942383,
33.3285446166992,
35.6963996887207,
-43.5586166381836,
-19.9510803222656,
34.7965278625488,
19.9488983154297,
6.20257139205933,
16.9955406188965,
-54.5780982971191,
-22.3693771362305,
62.1028480529785,
42.5089340209961,
41.6775817871094,
-16.7117309570313,
-43.8416786193848,
26.5547008514404,
57.5726127624512,
26.2590465545654,
-28.8200378417969,
-9.05296707153320,
44.7137870788574,
29.5549621582031,
-10.7688016891480,
64.6035919189453,
57.5217475891113,
-55.6335945129395,
42.9253082275391,
61.0864524841309,
-36.5865974426270,
-14.6722545623779,
-11.2911672592163,
27.1883354187012,
34.7706527709961,
-31.9438552856445,
-19.8672103881836,
13.1172943115234,
-31.4697685241699,
-25.2696266174316,
59.7656898498535,
-12.5694332122803,
-8.44999217987061,
66.1859207153320,
31.5259475708008,
23.8486728668213,
31.5441474914551,
22.7880210876465,
-23.3305587768555,
27.2971572875977,
1.19695091247559,
13.9097127914429,
36.9720458984375,
-28.9945621490479,
74.0922927856445,
23.5631027221680,
-47.5035934448242,
30.8609123229980,
52.8498153686523,
-4.34788227081299,
16.2034473419189,
65.7301101684570,
-5.01202297210693,
64.6790618896484,
22.3827533721924,
-9.45502662658691,
34.3106193542481,
-31.6029357910156,
50.1644554138184,
10.9813194274902,
-42.1497268676758,
17.3017883300781,
39.6518020629883,
-14.1285228729248,
29.1294708251953,
39.2219810485840,
-20.2560081481934,
51.0275650024414,
23.8325767517090,
43.3142547607422,
0.945938110351563,
0.334158897399902,
36.4101638793945,
-25.9261169433594,
7.37350082397461,
15.3280334472656,
26.8394031524658,
2.06720089912415,
-4.93438911437988,
53.2321281433106,
36.7992820739746,
-4.94238185882568,
-10.5109291076660,
-3.86231994628906,
28.6058044433594,
22.5595893859863,
15.0062084197998,
73.8214721679688,
23.7991600036621,
-37.8987236022949,
-1.80961513519287,
50.8403091430664,
54.6796722412109,
18.8200321197510,
5.73053550720215,
-28.3573379516602,
22.3867626190186,
10.9663143157959,
-21.3053207397461,
53.1498832702637,
48.8269195556641,
17.1416187286377,
-30.3069648742676,
9.79938697814941,
32.1501998901367,
-19.0693340301514,
35.9025764465332,
31.9630107879639,
11.5577249526978,
55.0954856872559,
15.6216802597046,
-37.5937881469727,
66.3242874145508,
40.8510589599609,
-55.0621261596680,
41.6453857421875,
8.36541366577148,
7.21025848388672,
13.1894941329956,
-13.8038539886475,
20.9457931518555,
-29.8119773864746,
0.965394973754883,
60.0906791687012,
41.6968193054199,
-45.5813827514648,
-39.2937393188477,
39.2932052612305,
40.5671310424805,
-27.2766723632813,
-7.87427902221680,
42.7057571411133,
-33.1020736694336,
19.7888889312744,
61.6133575439453,
-3.09898328781128,
23.1202640533447,
31.4587535858154,
29.3579120635986,
52.4384918212891,
12.7444410324097,
19.7824649810791,
70.5420913696289,
10.8150892257690,
-18.1472854614258,
80.9976043701172,
11.5455818176270,
-41.0251312255859,
73.1584091186523,
-17.9204502105713,
-32.5499877929688,
53.9478302001953,
56.1257553100586,
16.1006011962891,
-42.4887275695801,
-19.0340652465820,
-3.81310749053955,
44.8443222045898,
-17.5660171508789,
-46.9310455322266,
56.6755065917969,
7.21273994445801,
-33.6664237976074,
32.8121070861816,
1.31271219253540,
-23.6716346740723,
32.3359756469727,
24.6208839416504,
24.4314537048340,
-28.5077266693115,
-14.5863704681396,
39.2744369506836,
6.03423023223877,
30.5161838531494,
46.1644859313965,
18.4849090576172,
-10.2193794250488,
15.4570579528809,
10.5383090972900,
47.6055221557617,
65.2716217041016,
-0.501721143722534,
56.0329589843750,
31.0468215942383,
11.0051536560059,
-18.2828311920166,
-8.49192428588867,
56.6008224487305,
-9.21953010559082,
38.1721916198731,
-17.8919792175293,
-1.02942276000977,
57.3262863159180,
-23.3355140686035,
18.4799098968506,
41.7432823181152,
65.9743728637695,
-15.7642002105713,
-26.6313591003418,
18.2836380004883,
-20.0623378753662,
22.7709922790527,
-24.0385570526123,
-26.1953582763672,
29.1610164642334,
18.0138626098633,
-30.4347705841064,
-42.6262359619141,
-6.68032503128052,
26.0496196746826,
10.1800584793091,
-1.87908554077148,
65.8922653198242,
11.8514795303345,
-5.24831867218018,
-15.1884145736694,
20.5966129302979,
86.1697616577148,
-13.1502408981323,
-1.90467286109924,
26.1957473754883,
3.90901422500610,
30.5399246215820,
14.4003238677979,
-21.6562843322754,
45.8087692260742,
23.0804634094238,
-33.2539863586426,
0.188369274139404,
-49.2545890808106,
-13.6275682449341,
-20.3946113586426,
-19.8077354431152,
50.9559631347656,
-4.52710151672363,
2.34230422973633,
6.94026565551758,
21.4815101623535,
-6.70179414749146,
-45.4445037841797,
15.2696743011475,
24.1212596893311,
30.1881675720215,
-39.8489418029785,
17.4604148864746,
50.4113960266113,
-46.5879135131836,
23.1166057586670,
16.6640052795410,
32.5281105041504,
7.24121761322022,
-30.1323833465576,
55.5096282958984,
-52.2305908203125,
-19.2895774841309,
39.6221160888672,
-48.6506118774414,
-6.21966743469238,
-5.45612287521362,
18.5524215698242,
46.9239158630371,
47.2287330627441,
-16.7975769042969,
-19.5426483154297,
13.2828178405762,
-34.2447471618652,
32.8526229858398,
-32.1204185485840,
-52.4587631225586,
50.5438423156738,
38.2669143676758,
1.88702571392059,
9.18726825714111,
46.4113998413086,
45.5508842468262,
7.20235729217529,
-24.0532112121582,
-7.45231056213379,
30.4932365417480,
-0.655717849731445,
-42.8994674682617,
50.3731842041016,
26.1057777404785,
-16.5647125244141,
2.44792032241821,
-16.4860305786133,
-6.69712257385254,
-38.9765357971191,
2.96779966354370,
-30.5643997192383,
-15.3869590759277,
51.7222366333008,
-8.99725627899170,
20.7779579162598,
30.6648883819580,
-11.5363035202026,
-4.74769496917725,
1.38638186454773,
-16.4214744567871,
-15.1776065826416,
7.36452674865723,
-33.3624534606934,
-18.6082324981689,
46.2602920532227,
32.0671882629395,
3.74187898635864,
-51.1060752868652,
27.1112251281738,
26.1696147918701,
-48.3768386840820,
70.8401870727539,
12.7572250366211,
-56.1009216308594,
13.2632236480713,
16.0480594635010,
-24.4798927307129,
-21.5860710144043,
-0.147172972559929,
-20.0039787292480,
35.1945495605469,
18.9594058990479,
-31.2531185150147,
-5.95339488983154,
-18.6229095458984,
-15.8752355575562,
-15.3313627243042,
-33.6773757934570,
-23.7026233673096,
-0.725506901741028,
-12.6805047988892,
-3.83871746063232,
3.18414688110352,
-17.8677864074707,
-6.96294498443604,
-26.1745052337647,
-1.97877073287964,
7.48171520233154,
-24.6407852172852,
-29.6041622161865,
-28.6630287170410,
42.7756614685059,
-11.7230510711670,
-50.2756729125977,
54.3753166198731,
23.0538902282715,
0.546292603015900,
20.6840648651123,
-23.1433639526367,
-16.8540325164795,
4.43116617202759,
-55.5456542968750,
-18.7303409576416,
45.2177734375000,
23.8936462402344,
22.1762542724609,
-13.1381988525391,
10.9704284667969,
-4.24812507629395,
-28.4117507934570,
-1.64738011360168,
9.28935241699219,
-15.3270969390869,
-53.0679779052734,
-8.46103858947754,
21.0989875793457,
34.8205032348633,
29.3411064147949,
53.7045974731445,
-0.601284027099609,
-26.1759567260742,
7.34361362457275,
-27.2729377746582,
12.5459461212158,
50.6215972900391,
11.0469188690186,
3.17668151855469,
67.7710876464844,
-28.2801189422607,
-18.6351013183594,
57.3653106689453,
4.16944456100464,
19.7679061889648,
-3.17526531219482,
-25.2240371704102,
-9.96599864959717,
-4.61682653427124,
-25.3996562957764,
12.9120893478394,
52.7655830383301,
-35.7552413940430,
-23.4017829895020,
74.9176864624023,
-3.66041159629822,
-36.3776092529297,
64.6930389404297,
-25.7891464233398,
-32.9870376586914,
58.5977325439453,
9.31540679931641,
33.3580932617188,
-10.3509435653687,
-26.1798248291016,
27.9516201019287,
33.3335609436035,
25.9460601806641,
-4.44456386566162,
37.4257011413574,
15.3919963836670,
12.9572362899780,
24.4429073333740,
45.2648162841797,
54.2434997558594,
-33.6831588745117,
31.9579849243164,
15.8310098648071,
-48.7032966613770,
-18.5900554656982,
-14.0757694244385,
-18.4043979644775,
5.69306755065918,
28.1530036926270,
10.6950035095215,
41.3404235839844,
-14.8288974761963,
27.8658542633057,
15.6721658706665,
1.11386537551880,
30.5543460845947,
-41.7824020385742,
49.8755950927734,
15.2897338867188,
22.7489395141602,
67.1681671142578,
-3.18734550476074,
-26.0937500000000,
-28.4267616271973,
18.7695007324219,
30.5592994689941,
25.9389877319336,
-2.62192773818970,
-23.9705371856689,
28.8538303375244,
36.2681236267090,
45.3070907592773,
41.1078033447266,
-18.2958106994629,
-17.3001365661621,
1.34690999984741,
73.0919647216797,
0.700548171997070,
-11.8935642242432,
62.0394897460938,
-48.4350242614746,
-22.5004577636719,
-13.8800334930420,
-17.5464534759522,
8.60585117340088,
-40.2530441284180,
-39.1971778869629,
-2.25032401084900,
-28.2204589843750,
-31.3406028747559,
18.3309936523438,
-12.2267503738403,
14.4292745590210,
7.83662033081055,
14.2722759246826,
35.8429527282715,
23.9721641540527,
27.1046543121338,
-34.7373542785645,
6.33200931549072,
-0.846389770507813,
-31.1290893554688,
11.9134063720703,
-43.9829177856445,
33.9466781616211,
59.0805816650391,
-42.5710830688477,
56.7882614135742,
6.99605894088745,
-52.6499328613281,
-6.42529916763306,
-33.2865600585938,
22.5884246826172,
-26.1008415222168,
31.3288135528564,
67.5431900024414,
-32.9579772949219,
20.9146423339844,
-19.0837249755859,
-13.1874876022339,
36.0604667663574,
3.89232015609741,
16.5418338775635,
10.1575965881348,
-18.7240772247314,
-2.56517791748047,
41.7700080871582,
19.1533432006836,
33.3564834594727,
10.6850624084473,
29.5654563903809,
56.0363616943359,
-34.0882606506348,
-11.8102025985718,
54.2170486450195,
25.3838748931885,
2.60648155212402,
55.6782531738281,
2.20367240905762,
5.00955963134766,
57.1772766113281,
21.6674289703369,
14.0980701446533,
17.1497344970703,
-2.18119907379150,
-20.8548374176025,
7.72727394104004,
19.5491428375244,
40.9993171691895,
30.6033096313477,
54.5774841308594,
4.05429267883301,
-47.4841270446777,
70.8455963134766,
-0.395256996154785,
-31.9828987121582,
75.1746749877930,
28.9414787292480,
-37.3396301269531,
-8.59612464904785,
16.2561588287354,
-7.40290689468384,
0.330922603607178,
-5.94658899307251,
49.3432006835938,
26.5889511108398,
14.0818138122559,
24.6641139984131,
-33.3654022216797,
52.8707351684570,
-32.2836875915527,
-2.62553787231445,
68.0977325439453,
-37.0496978759766,
4.08697605133057,
25.3297386169434,
33.5510635375977,
-23.2238559722900,
31.7904396057129,
37.0366783142090,
-54.1800231933594,
19.6985530853272,
-18.6349182128906,
18.1512107849121,
37.6811981201172,
25.7944030761719,
79.2059020996094,
10.2888078689575,
-35.1920013427734,
9.55484580993652,
22.3627071380615,
-49.2335777282715,
11.2424716949463,
35.4597587585449,
-39.2989921569824,
-39.9218215942383,
0.276444435119629,
-6.36681175231934,
1.11293554306030,
28.4259910583496,
4.36021375656128,
11.3034706115723,
4.25990676879883,
56.3382225036621,
33.3688163757324,
30.2258892059326,
67.5444412231445,
21.3497638702393,
66.4284057617188,
30.0841636657715,
14.8519554138184,
54.2428588867188,
-19.7489891052246,
41.7007675170898,
64.7037963867188,
-43.7968406677246,
-13.6975927352905,
20.2667331695557,
1.89842820167542,
10.8582363128662,
55.7421493530273,
30.0005397796631,
-4.30161142349243,
16.5992202758789,
21.2838420867920,
9.73086261749268,
-35.1211433410645,
26.4294242858887,
12.1077966690063,
-45.9546356201172,
62.5536880493164,
21.9944629669189,
-37.7038078308106,
53.1483535766602,
54.0821075439453,
27.6364974975586,
31.7636680603027,
-4.90464067459106,
48.7117805480957,
75.0743560791016,
-8.92318344116211,
-23.6848602294922,
-16.4531650543213,
-4.09195613861084,
4.58173751831055,
-18.5046653747559,
-29.1808242797852,
-7.96646976470947,
-39.5808715820313,
-50.7249374389648,
55.6254348754883,
7.71734619140625,
-45.5355682373047,
21.7131881713867,
-26.6586093902588,
-12.6229152679443,
32.8874969482422,
9.01266574859619,
16.2936859130859,
31.8458557128906,
-2.30802822113037,
0.411577224731445,
50.4035339355469,
-4.79551410675049,
14.2802696228027,
-8.75318050384522,
-24.3100357055664,
23.1866569519043,
-19.3623828887939,
5.30543470382690,
-21.2280769348145,
14.1183052062988,
30.6622009277344,
-32.0308570861816,
-17.1967029571533,
16.6652107238770,
3.30759453773499,
5.04598522186279,
46.3922691345215,
41.6232910156250,
-5.94453811645508,
-14.9437942504883,
70.8914108276367,
-2.01689815521240,
19.0873146057129,
44.6432189941406,
1.85746026039124,
44.8346557617188,
-7.74031591415405,
8.00251007080078,
-17.0011749267578,
45.7470016479492,
18.1699943542480,
-49.8506927490234,
48.1676101684570,
-4.32596063613892,
-9.99264717102051,
25.3679618835449,
45.8425521850586,
38.1036376953125,
-26.9417705535889,
21.7685127258301,
42.2427177429199,
7.61120605468750,
-12.0280265808105,
-23.5258846282959,
51.7395553588867,
7.80849933624268,
-63.7626190185547,
10.3294181823730,
58.3918457031250,
25.1054611206055,
25.4344062805176,
9.02758407592773,
-28.2348251342773,
36.1854476928711,
-11.2411327362061,
-11.0873517990112,
3.79045414924622,
-58.7148590087891,
-9.74457359313965,
41.0963439941406,
31.0087089538574,
22.2482261657715,
38.7229347229004,
-41.6526870727539,
13.9349040985107,
87.5686264038086,
-13.0035743713379,
-37.9259262084961,
-4.51761150360107,
28.7606315612793,
-1.03780937194824,
4.39062356948853,
27.9642925262451,
-7.42965793609619,
-42.4561691284180,
-37.5470123291016,
14.8328456878662,
27.1574230194092,
58.4166297912598,
6.81324958801270,
-35.7194938659668,
-4.94510746002197,
8.37878227233887,
10.5689020156860,
1.77981567382813,
56.8362998962402,
31.1736488342285,
1.69834995269775,
-9.65771198272705,
45.1486892700195,
18.0619087219238,
-9.14599514007568,
38.8277397155762,
-33.3987541198731,
46.2666587829590,
10.3468055725098,
-24.4842758178711,
-7.03304052352905,
-27.6405639648438,
59.2075538635254,
9.66270828247070,
8.41573429107666,
32.9329681396484,
-20.2796230316162,
-8.59207630157471,
16.7150249481201,
-17.7643394470215,
14.5834541320801,
15.5557289123535,
-50.1222877502441,
33.7571945190430,
-14.7503356933594,
-20.5584812164307,
48.0376205444336,
-69.4186477661133,
-12.5933303833008,
36.9961891174316,
-40.8620185852051,
-17.2890319824219,
5.69771718978882,
7.64312458038330,
20.8052959442139,
-16.1873321533203,
-46.7680130004883,
-2.85185194015503,
-0.287467002868652,
-49.5932693481445,
37.8511657714844,
50.0761413574219,
-42.9755630493164,
37.2279205322266,
40.5360450744629,
31.6060543060303,
0.690052151679993,
-31.6560306549072,
40.2885322570801,
-5.89106845855713,
61.9901275634766,
27.2354316711426,
-52.5833969116211,
25.3413276672363,
33.0794448852539,
-3.33574867248535,
-60.2980003356934,
45.6904716491699,
-8.18734169006348,
-45.3692703247070,
24.6035861968994,
-4.11535835266113,
26.9633426666260,
-6.94771718978882,
29.7327251434326,
-20.3607826232910,
-34.0204048156738,
-24.7895545959473,
24.7954635620117,
25.3107166290283,
-15.0416927337646,
49.9768333435059,
-24.8520431518555,
45.3653450012207,
31.4080142974854,
-11.0930671691895,
-12.9896821975708,
-33.0046463012695,
-25.8098106384277,
-12.5423269271851,
26.8992843627930,
-5.28325748443604,
24.3127803802490,
-40.7610359191895,
30.6033058166504,
67.8188323974609,
-18.5189609527588,
24.2703533172607,
24.7042160034180,
69.7315979003906,
-1.54086220264435,
0.618056297302246,
69.6073989868164,
-13.9974040985107,
-46.7248115539551,
-20.8334693908691,
31.0025215148926,
5.44929742813110,
18.7653656005859,
-3.13350915908813,
-0.493840456008911,
21.5780429840088,
-80.5932540893555,
30.9709777832031,
46.4099426269531,
-55.2379608154297,
-18.4400386810303,
9.07194995880127,
18.4047031402588,
-29.9318904876709,
41.2634582519531,
56.4320526123047,
9.63980007171631,
47.2216873168945,
-41.0865135192871,
38.3216934204102,
42.8494796752930,
-46.6066741943359,
21.1683216094971,
-14.4143295288086,
3.98850679397583,
-30.9220619201660,
-8.90182685852051,
13.2465381622314,
-40.1495437622070,
-36.3274574279785,
-27.4342365264893,
21.6757411956787,
-37.4373245239258,
-21.6174259185791,
40.5154838562012,
47.2633895874023,
-24.9780521392822,
4.29905080795288,
78.1188659667969,
5.70079612731934,
-0.958901166915894,
-20.3408699035645,
-2.48872375488281,
61.9094848632813,
33.6872825622559,
-41.2444610595703,
13.9849815368652,
27.7686920166016,
-43.7292098999023,
-17.9847431182861,
35.2062072753906,
34.1907272338867,
0.221837997436523,
-37.9098625183106,
-2.29625320434570,
66.4623489379883,
-3.47371578216553,
15.5777359008789,
8.36769294738770,
-25.3158454895020,
-14.5031232833862,
-30.7545471191406,
61.9339942932129,
19.4716014862061,
-15.1773977279663,
18.7316036224365,
25.6319065093994,
54.7086105346680,
7.22586774826050,
41.5717849731445,
-0.304626464843750,
-36.3575935363770,
48.6325263977051,
-15.6988029479980,
-3.90502023696899,
-1.37946987152100,
-44.3522186279297,
-0.781435012817383,
14.2412824630737,
49.1281738281250,
9.76078128814697,
27.8695621490479,
60.7381401062012,
27.7434234619141,
57.5561828613281,
51.3081054687500,
-27.0602321624756,
5.44427490234375,
56.6080627441406,
-17.1700763702393,
17.3630943298340,
-20.1678791046143,
3.43199443817139,
58.7232666015625,
-0.422620773315430,
-8.11802577972412,
-15.9734268188477,
35.7057609558106,
-2.98367714881897,
45.7764511108398,
58.0419845581055,
-2.88008093833923,
42.0850906372070,
0.355934143066406,
41.4098014831543,
17.7628688812256,
1.21930193901062,
56.3015098571777,
-24.7256622314453,
-33.3846511840820,
-1.95895767211914,
35.2094612121582,
-28.7553901672363,
-58.8458480834961,
37.9885559082031,
-36.9105987548828,
-11.7490310668945,
64.4479675292969,
-6.44939613342285,
29.7832508087158,
17.8039989471436,
-13.8872299194336,
-9.86024188995361,
-6.61847686767578,
60.2302703857422,
-29.5553398132324,
16.3149719238281,
29.2250976562500,
-41.7377204895020,
11.1220722198486,
-32.3993148803711,
3.83432960510254,
37.8171653747559,
23.6717262268066,
-3.25968313217163,
-1.09217095375061,
-14.8662242889404,
37.0436477661133,
16.2839164733887,
-52.3217926025391,
3.67032861709595,
-34.4770812988281,
26.8614158630371,
-19.4771003723145,
-17.4228515625000,
62.7128334045410,
-36.8764762878418,
4.81894207000732,
33.4944648742676,
22.4240818023682,
33.3035354614258,
-23.1148853302002,
16.0271625518799,
63.3911819458008,
-12.1901187896729,
4.30377435684204,
-3.99570655822754,
-24.4766693115234,
71.4342803955078,
-10.2141523361206,
-17.6080303192139,
45.5040054321289,
-16.8371124267578,
2.65961003303528,
-2.40878868103027,
-23.1071853637695,
-24.2242469787598,
-26.4033298492432,
-37.0796852111816,
-24.4415321350098,
-30.3564224243164,
-10.9388275146484,
22.4109745025635,
-17.4205017089844,
-30.5747795104980,
-14.6049728393555,
41.8439140319824,
28.7075920104980,
15.6586685180664,
17.7692222595215,
-5.84992170333862,
19.8527011871338,
70.3461990356445,
11.4481048583984,
7.35960006713867,
59.6343498229981,
-32.9231758117676,
1.96264314651489,
-10.5539951324463,
19.2147960662842,
52.6712341308594,
-31.1561698913574,
30.7315101623535,
28.9917984008789,
-27.7222137451172,
-15.3543720245361,
-2.59024763107300,
15.5117444992065,
36.6561164855957,
-23.0408020019531,
-15.3042030334473,
18.4654884338379,
-11.8202037811279,
-18.6175613403320,
11.9164390563965,
36.7703552246094,
-39.2562789916992,
-16.1156997680664,
18.0891952514648,
-6.37044286727905,
34.2895545959473,
-25.9956722259522,
-38.3318862915039,
10.4354028701782,
-16.7227344512939,
21.6828460693359,
4.72433519363403,
-19.5941829681397,
17.2572555541992,
15.3442726135254,
39.3425827026367,
23.6688060760498,
-1.57534456253052,
20.0668506622314,
29.2030735015869,
-23.6982727050781,
8.03443908691406,
76.8154144287109,
-14.8183917999268,
-15.0137882232666,
34.1151466369629,
-20.3625240325928,
0.727823257446289,
41.7454223632813,
6.85002231597900,
7.19063091278076,
64.1547393798828,
-8.46708774566650,
-30.7005805969238,
51.6186485290527,
25.9331398010254,
-8.86004447937012,
10.6717977523804,
49.7279090881348,
38.9490470886231,
50.3447570800781,
40.6351928710938,
54.2870025634766,
31.2979011535645,
-21.8994865417480,
2.99286961555481,
4.02708625793457,
59.9816741943359,
20.2181282043457,
11.3234128952026,
16.1997947692871,
-27.2997779846191,
20.3146896362305,
-13.7719440460205,
31.1599693298340,
12.7558593750000,
-18.8929443359375,
72.6979446411133,
45.1897506713867,
-4.55756092071533,
-25.7431926727295,
35.5328788757324,
28.3443946838379,
31.4970016479492,
58.3020248413086,
23.1401996612549,
55.5818176269531,
31.2763462066650,
-17.2270812988281,
-13.5546712875366,
49.1476364135742,
0.692180633544922,
-44.2394409179688,
33.9599914550781,
39.8068466186523,
-2.38597488403320,
-6.22223615646362,
7.76016998291016,
-34.2525100708008,
2.79831123352051,
40.0559425354004,
-36.2713928222656,
-38.0996818542481,
53.7876205444336,
15.9202384948730,
-55.0909500122070,
19.7736282348633,
-11.2428150177002,
18.2387886047363,
18.1292457580566,
-14.9536285400391,
3.19338417053223,
-29.5601406097412,
61.4797210693359,
20.8217105865479,
26.1851310729980,
33.3527069091797,
22.5582427978516,
7.04780626296997,
-27.0471725463867,
6.66812658309937,
-27.1397323608398,
45.7833213806152,
35.2485733032227,
-7.26186895370483,
-26.7099571228027,
0.841989040374756,
-28.8180084228516,
2.78751277923584,
45.1221427917481,
-39.2883987426758,
68.4976577758789,
13.7305059432983,
19.7522563934326,
66.7203521728516,
11.2675104141235,
61.2636566162109,
10.4262981414795,
46.8433723449707,
72.7856140136719,
32.5776367187500,
45.8539733886719,
27.9451160430908,
-12.3722991943359,
-14.8922414779663,
-1.76400375366211,
-38.9745597839356,
25.5799179077148,
-10.7901830673218,
-66.7759017944336,
11.7229251861572,
-7.85123777389526,
-6.31813621520996,
-13.5871477127075,
53.7774810791016,
37.9375801086426,
-55.8284606933594,
36.5530815124512,
25.1457309722900,
16.8916587829590,
33.8755989074707,
45.9927825927734,
43.6567115783691,
14.9177551269531,
36.6127777099609,
22.8944816589355,
63.3382339477539,
28.9677143096924,
-13.8157501220703,
22.2588119506836,
23.1464500427246,
-31.8826789855957,
-4.71266889572144,
68.3008270263672,
-21.7160415649414,
-27.4331665039063,
14.4456996917725,
-18.2478542327881,
29.1728477478027,
30.4563808441162,
-40.0121154785156,
-2.97217559814453,
30.3354034423828,
-2.84114813804626,
16.3014450073242,
-14.1724319458008,
-22.4790210723877,
40.8332748413086,
38.1168441772461,
38.3483505249023,
-12.7562246322632,
-42.1885986328125,
20.2439842224121,
50.9906196594238,
25.3993530273438,
1.91967082023621,
28.7111263275147,
23.4803199768066,
23.3179264068604,
44.6000366210938,
59.3462448120117,
17.2899703979492,
26.7773475646973,
58.4159431457520,
-17.4411449432373,
15.0270442962646,
56.1450080871582,
21.0994014739990,
-69.0478591918945,
5.09762191772461,
49.7148818969727,
-45.5886192321777,
52.9135780334473,
0.689210891723633,
18.5724525451660,
49.3952255249023,
16.1863670349121,
69.1786193847656,
19.0524139404297,
-32.0758972167969,
11.8023500442505,
46.4488945007324,
-43.0999832153320,
45.3818168640137,
53.5440559387207,
-12.6852951049805,
24.5012454986572,
68.6518478393555,
0.644798278808594,
-25.0244140625000,
22.4110221862793,
-26.9663047790527,
56.0622253417969,
-41.1066246032715,
-23.9470233917236,
47.3654594421387,
-49.7178878784180,
-1.00500345230103,
13.2826862335205,
19.1692123413086,
10.9308719635010,
-25.3946495056152,
20.2099933624268,
6.20047903060913,
-6.55436134338379,
44.6374893188477,
41.6889419555664,
53.4432525634766,
21.9106044769287,
21.5735778808594,
-40.0394020080566,
18.3276710510254,
53.8893318176270,
-45.7857284545898,
27.6492729187012,
8.48558425903320,
39.7182159423828,
-12.6577987670898,
-10.3083076477051,
22.7048244476318,
-35.9195175170898,
-3.27864050865173,
-30.2665672302246,
83.0504837036133,
21.7724895477295,
-39.9030761718750,
42.8919563293457,
-10.8230066299438,
-8.78018188476563,
-31.7466354370117,
-6.99928045272827,
-0.885927975177765,
-6.03365993499756,
55.7798538208008,
-2.34716129302979,
55.1088829040527,
46.9629821777344,
-31.1108551025391,
59.2943267822266,
28.4881763458252,
-3.02081847190857,
-26.0490798950195,
2.12201642990112,
52.2857971191406,
36.3789215087891,
33.3697433471680,
-44.2136230468750,
-6.05707740783691,
34.2023963928223,
-7.06046581268311,
-20.9901542663574,
-28.3446979522705,
-27.0320968627930,
-14.1907615661621,
54.6773490905762,
2.02973747253418,
-34.5364837646484,
46.6716117858887,
-9.33547019958496,
20.4435863494873,
61.4626083374023,
-33.4396400451660,
18.3552131652832,
71.9138641357422,
12.6671762466431,
-10.2213068008423,
19.2592582702637,
61.5161514282227,
8.82384872436523,
27.3938426971436,
71.7567520141602,
-9.19920158386231,
-12.6296634674072,
-22.1214065551758,
4.47017383575439,
-4.26424884796143,
-13.4012422561646,
11.7948246002197,
29.7340183258057,
19.6815605163574,
-37.7666778564453,
25.9716949462891,
13.8955497741699,
43.7578544616699,
-12.0044956207275,
-22.8140144348145,
48.6261444091797,
-44.0215263366699,
34.6378326416016,
50.1198539733887,
18.4802589416504,
19.3201770782471,
0.846575736999512,
55.6900482177734,
54.4950752258301,
22.8816528320313,
-28.1156120300293,
-9.59991455078125,
-10.1330461502075,
-30.8498363494873,
-5.41248035430908,
50.6132202148438,
35.7113037109375,
-40.4300880432129,
53.5596389770508,
7.05552673339844,
-32.1788558959961,
66.7733764648438,
17.9806594848633,
-43.4667320251465,
48.5349769592285,
42.9493103027344,
6.20294475555420,
46.5019302368164,
-0.829537868499756,
38.2542228698731,
-7.98878574371338,
18.2786102294922,
71.7698211669922,
44.5506515502930,
-4.58509397506714,
-8.83385753631592,
66.8678665161133,
-49.5752182006836,
-9.23431205749512,
36.6374511718750,
1.15344250202179,
24.6801853179932,
-12.7608985900879,
2.28001785278320,
28.6821079254150,
-9.05294418334961,
-34.0633201599121,
10.3175277709961,
-32.6496810913086,
9.25427436828613,
55.3108520507813,
9.35226058959961,
47.3418083190918,
-15.4344911575317,
-24.8237247467041,
23.9195384979248,
-7.15045499801636,
-34.4795303344727,
-12.7085247039795,
56.3139038085938,
-44.2798461914063,
-42.3729553222656,
76.9597244262695,
-9.82863330841065,
-22.3456954956055,
5.47433710098267,
29.0903663635254,
12.7211675643921,
-50.0141944885254,
79.1575851440430,
35.5149154663086,
-50.8646888732910,
-3.30526208877563,
-34.4558715820313,
22.5854110717773,
13.4499893188477,
-23.6846065521240,
-17.7831268310547,
8.73077487945557,
-17.2969474792480,
-9.25282478332520,
47.8911895751953,
-12.3159656524658,
26.8992938995361,
-35.7556381225586,
19.0310401916504,
105.896560668945,
-40.1868286132813,
0.945231676101685,
37.0206527709961,
-46.0569686889648,
-24.3391265869141,
-1.35437965393066,
-45.8345489501953,
0.368103027343750,
7.02522945404053,
-10.6959314346313,
42.5059852600098,
29.9226646423340,
-5.14660549163818,
10.0487642288208,
-2.75015068054199,
-14.3655624389648,
-14.2676973342896,
-32.7381744384766,
0.150342941284180,
-21.8170585632324,
1.79507160186768,
41.0706214904785,
-7.87374973297119,
32.3147277832031,
48.8723258972168,
-22.4768371582031,
1.27923190593719,
-12.7565336227417,
-7.28539562225342,
21.5433235168457,
-42.1318359375000,
24.0743274688721,
-0.460560798645020,
-0.278153121471405,
13.0703086853027,
-50.8268165588379,
-28.5561141967773,
-2.97192955017090,
55.4211959838867,
-0.594694137573242,
-29.8394985198975,
0.496955394744873,
-17.5999488830566,
-6.57389974594116,
42.7944068908691,
10.4623441696167,
-4.77598190307617,
40.7691726684570,
17.0451965332031,
-12.7659645080566,
-11.2323875427246,
-1.03576660156250,
-20.2248649597168,
25.4409236907959,
-7.12281799316406,
-28.9704303741455,
-33.1237831115723,
-28.1496257781982,
-19.4153022766113,
-18.4993553161621,
22.9674568176270,
-23.5145034790039,
12.5213327407837,
-17.5708160400391,
12.2254533767700,
64.8755111694336,
14.3150405883789,
-28.4845142364502,
-5.37509346008301,
24.9301643371582,
-49.5097236633301,
-19.9378395080566,
16.7554397583008,
40.7440681457520,
30.7014255523682,
-1.40002989768982,
-24.9906139373779,
35.2058486938477,
32.3171768188477,
19.2514858245850,
24.2777214050293,
-16.8772506713867,
58.2688446044922,
-39.7098617553711,
-36.9349975585938,
26.0281925201416,
14.3613891601563,
26.5664005279541,
6.85600423812866,
75.1172103881836,
18.6628837585449,
-29.0750465393066,
52.2532119750977,
4.78822898864746,
-41.0526885986328,
62.7949028015137,
6.95290374755859,
-55.8194198608398,
63.6542053222656,
20.6185703277588,
-40.7382202148438,
17.9261608123779,
37.3762359619141,
-31.0098915100098,
-7.80078697204590,
60.8299064636231,
-50.7339401245117,
-19.7598190307617,
60.1945304870606,
5.40464115142822,
-23.6865329742432,
-46.5360794067383,
21.6099147796631,
34.5188522338867,
-80.2071075439453,
-12.6697120666504,
23.3256835937500,
-16.2929782867432,
37.8974266052246,
-13.9593486785889,
11.7151527404785,
18.4897537231445,
14.9327697753906,
39.7380981445313,
39.4562072753906,
47.8620758056641,
-30.3134918212891,
52.5174293518066,
68.6185760498047,
5.93795108795166,
6.72099494934082,
-9.77739524841309,
5.81586742401123,
1.25982928276062,
47.3278617858887,
20.5475311279297,
8.39594650268555,
41.2594261169434,
-28.7256469726563,
-0.484106063842773,
67.9315795898438,
46.9772644042969,
13.3700141906738,
-11.0997610092163,
45.0328483581543,
45.3236236572266,
-19.6615409851074,
19.2624435424805,
-21.5308361053467,
-27.0647640228272,
44.2427749633789,
29.9945106506348,
-6.71984720230103,
-13.0113029479980,
50.6760482788086,
-14.4201393127441,
-21.3179988861084,
94.0110778808594,
25.7299995422363,
-34.6054763793945,
10.9143562316895,
48.3695793151856,
11.4631729125977,
19.5237445831299,
66.2199096679688,
42.7203216552734,
18.9000358581543,
9.88801574707031,
-16.7594108581543,
-30.8884353637695,
-4.82127237319946,
21.5803356170654,
34.5570602416992,
-16.4844093322754,
25.1186752319336,
28.7982444763184,
-46.2933654785156,
-11.0273828506470,
16.8672389984131,
69.2411041259766,
16.8705863952637,
-28.3001518249512,
39.9064636230469,
-14.5651187896729,
32.7878189086914,
78.5433731079102,
-7.01758337020874,
32.0186500549316,
14.2662696838379,
19.4002113342285,
24.6864490509033,
-10.1221160888672,
37.4634017944336,
-28.3587341308594,
-17.8923835754395,
47.9288597106934,
50.5939750671387,
-10.2917938232422,
-50.3397827148438,
23.0299339294434,
-11.0341606140137,
-6.42543601989746,
-14.7803716659546,
-30.8292312622070,
-18.5580348968506,
-11.9209899902344,
54.0662918090820,
-17.9045925140381,
31.3498668670654,
29.4579524993897,
-34.2540740966797,
30.8525180816650,
38.3627586364746,
26.1262340545654,
-46.8425559997559,
7.27324676513672,
-7.87022781372070,
-46.4817428588867,
21.7510108947754,
5.05584621429443,
22.7526359558105,
-15.9897356033325,
-27.4451637268066,
-7.08769273757935,
-8.13629817962647,
28.4665298461914,
6.34650754928589,
-13.5552291870117,
-1.86115074157715,
32.0075378417969,
25.4893951416016,
38.6110992431641,
54.0615539550781,
-2.62074899673462,
34.5171012878418,
64.4903182983398,
14.5729169845581,
-30.7266578674316,
45.2270393371582,
49.4423751831055,
-52.1583442687988,
46.3755645751953,
32.7635459899902,
-29.3623523712158,
38.3968620300293,
15.7256803512573,
41.2883300781250,
45.0670700073242,
40.0583305358887,
-6.74204063415527,
-37.6845588684082,
68.9996566772461,
45.8479270935059,
39.4246215820313,
-9.30648994445801,
-9.78648281097412,
55.7946891784668,
50.0391731262207,
44.0077667236328,
16.2087211608887,
33.9754295349121,
-31.9273338317871,
28.0991859436035,
48.1192092895508,
10.2487173080444,
44.0909347534180,
-50.2277221679688,
2.48292064666748,
32.0647163391113,
-44.3728332519531,
44.2273750305176,
21.8937683105469,
-61.8193740844727,
52.3279228210449,
32.3003120422363,
17.6693592071533,
41.1740913391113,
-32.9253921508789,
21.0964660644531,
46.1145858764648,
20.9937992095947,
-8.76617431640625,
-15.5579900741577,
32.7715721130371,
54.9272232055664,
-13.7782535552979,
14.1527748107910,
61.4876861572266,
-29.2220840454102,
20.3376235961914,
73.2441101074219,
45.1143722534180,
29.2654705047607,
-21.0053062438965,
-3.28730773925781,
56.7718734741211,
24.5293998718262,
27.6347198486328,
65.8504180908203,
33.1746826171875,
-8.06091117858887,
-15.8508882522583,
72.7110443115234,
47.1760559082031,
-41.6551551818848,
59.3257369995117,
17.9152183532715,
-42.5359153747559,
57.2181358337402,
21.8675880432129,
2.74190211296082,
11.9237728118896,
7.65637397766113,
11.7708826065063,
-34.9825744628906,
5.28929996490479,
25.2644882202148,
-32.8611297607422,
-26.1347122192383,
-1.28715825080872,
-17.5706996917725,
-23.3918571472168,
31.5490646362305,
32.8340530395508,
14.0730266571045,
33.9126548767090,
-32.2886466979981,
-26.4556198120117,
18.0079574584961,
35.0637130737305,
48.0826263427734,
-29.8800621032715,
3.02445411682129,
48.3135108947754,
26.9076976776123,
51.0194168090820,
-15.6145000457764,
-8.76966190338135,
29.4238166809082,
-20.3957462310791,
18.2899856567383,
5.12388992309570,
-38.1639289855957,
-25.8721275329590,
-17.5419960021973,
-23.8491878509522,
-36.3819961547852,
-23.4447174072266,
-20.1872997283936,
-36.8836288452148,
17.0025253295898,
59.6352539062500,
-32.3902893066406,
7.29472923278809,
55.1413192749023,
18.4795799255371,
16.7593860626221,
35.0133323669434,
59.7378349304199,
18.6896877288818,
37.6160850524902,
10.6088981628418,
-10.3063659667969,
-6.91622543334961,
40.9050788879395,
18.1104335784912,
-61.7187385559082,
-6.51832485198975,
-15.4386739730835,
40.6570243835449,
21.5727825164795,
-3.25037860870361,
48.9753150939941,
-2.44684982299805,
2.53355240821838,
51.8402519226074,
26.6810550689697,
-39.0172080993652,
0.141798019409180,
71.6700592041016,
31.5108642578125,
-25.0025863647461,
24.9715538024902,
8.49619388580322,
-3.48845100402832,
28.3754501342773,
23.5426998138428,
56.4216346740723,
10.3287267684937,
5.13723230361939,
42.1328964233398,
26.0386276245117,
30.7331542968750,
-3.76210308074951,
-20.4648780822754,
7.82893276214600,
32.4918937683106,
25.4602203369141,
10.0043907165527,
57.9816284179688,
14.1611938476563,
-45.2823333740234,
49.3143348693848,
60.9888992309570,
-38.9298515319824,
42.8019828796387,
24.1539554595947,
-50.2818031311035,
77.2063064575195,
-1.16053962707520,
-20.3677310943604,
84.1825561523438,
28.7848205566406,
-42.6825180053711,
29.3012886047363,
78.4426956176758,
-49.8238983154297,
26.9994812011719,
60.4473495483398,
-32.2403144836426,
-48.1820030212402,
8.63057518005371,
51.7020187377930,
-39.8904647827148,
26.7689399719238,
39.2513122558594,
-6.63908052444458,
15.0337772369385,
41.5158958435059,
33.6276435852051,
-47.6322517395020,
2.00016307830811,
40.8188018798828,
12.3728122711182,
8.64328193664551,
26.4216194152832,
-3.83852481842041,
14.9708318710327,
21.1217288970947,
-1.44483470916748,
68.7785644531250,
-23.0277976989746,
-10.0786933898926,
72.3174209594727,
15.4189119338989,
7.61523723602295,
17.5768375396729,
60.3317260742188,
-11.6199579238892,
-15.1872224807739,
61.2580261230469,
-17.3785171508789,
-65.0447311401367,
17.2135486602783,
37.0745544433594,
-6.41529130935669,
33.4023208618164,
-11.8439025878906,
-9.31479072570801,
31.6794586181641,
33.2043800354004,
54.9507904052734,
38.7577705383301,
53.6991386413574,
49.5100097656250,
23.8800926208496,
46.9535064697266,
40.7361221313477,
-37.8429908752441,
23.8434467315674,
67.1729049682617,
-30.3034133911133,
9.17603015899658,
20.9930896759033,
-37.8769721984863,
-15.3055610656738,
-2.89224267005920,
-17.8194465637207,
-12.4648628234863,
14.4735584259033,
39.8635482788086,
-9.37529468536377,
-42.9972114562988,
39.3112335205078,
-4.95822334289551,
-19.3212299346924,
19.3667201995850,
-29.6071987152100,
13.9575309753418,
65.0019378662109,
25.8061180114746,
-36.6975631713867,
14.7824888229370,
-6.08479547500610,
-23.2334232330322,
1.77902531623840,
-58.1380271911621,
2.15533924102783,
15.3631706237793,
-16.9805412292480,
20.3671016693115,
17.5564823150635,
24.1621761322022,
0.170104026794434,
-22.3644981384277,
3.59510350227356,
-42.0409851074219,
6.58788108825684,
70.8509902954102,
13.9111680984497,
-15.4408950805664,
19.1576576232910,
14.6972579956055,
-35.4395751953125,
5.11794185638428,
49.5444412231445,
51.3456268310547,
-14.2538862228394,
-33.1614036560059,
16.9994144439697,
40.4960861206055,
-17.0445613861084,
-21.5320472717285,
33.8034286499023,
4.48071002960205,
26.8492393493652,
-27.7567901611328,
-5.89787578582764,
24.4921875000000,
13.2831382751465,
13.0737562179565,
-6.18291282653809,
65.7141876220703,
-0.152230262756348,
19.3717193603516,
29.0989704132080,
1.38684511184692,
-1.55935311317444,
-20.4429798126221,
78.9515380859375,
-5.57095670700073,
8.74248218536377,
47.5300407409668,
-27.6762008666992,
28.8817462921143,
53.4923782348633,
52.3045043945313,
-10.5252552032471,
15.7555923461914,
20.8863296508789,
-57.4077033996582,
33.8726196289063,
77.3630828857422,
25.5315818786621,
-7.27851867675781,
-13.7040758132935,
-15.0887966156006,
11.7699928283691,
39.7993049621582,
24.3077125549316,
12.2301788330078,
12.6354875564575,
13.1522274017334,
-25.2345485687256,
7.05638599395752,
40.9994125366211,
-8.02537918090820,
16.7209701538086,
59.4380264282227,
-6.57443428039551,
-20.6190872192383,
50.4820518493652,
-4.38051652908325,
-42.3616676330566,
32.8771934509277,
65.4839630126953,
14.3479957580566,
-47.9348640441895,
-2.14776420593262,
9.69304180145264,
20.6416683197022,
55.6135978698731,
7.35804653167725,
34.1065444946289,
-14.1147937774658,
-26.1641635894775,
8.46293449401856,
-2.00508975982666,
66.3650817871094,
-19.3494148254395,
-29.3480148315430,
25.0172672271729,
-14.3212060928345,
45.7885742187500,
-0.423778295516968,
-51.1330261230469,
45.0714569091797,
26.6029891967773,
-49.5553894042969,
-13.9840545654297,
61.1558837890625,
4.95441246032715,
-61.4596061706543,
28.2769508361816,
19.2136116027832,
-20.6130008697510,
40.4581794738770,
-4.79346561431885,
-44.4240303039551,
13.5438432693481,
-43.2840080261231,
-30.2341899871826,
34.6547012329102,
-22.1940364837647,
27.4854946136475,
21.6517276763916,
34.2438163757324,
23.4457111358643,
-52.4544982910156,
55.6914024353027,
8.35461997985840,
-21.9833946228027,
68.6715316772461,
18.5308952331543,
-29.6981391906738,
-31.3459300994873,
16.9051170349121,
48.4705467224121,
7.20845937728882,
-33.1732559204102,
37.7505798339844,
24.8458900451660,
-36.7452735900879,
39.9944305419922,
53.2634773254395,
14.4067192077637,
-38.0562324523926,
11.4047908782959,
77.4181976318359,
29.6557903289795,
40.0741233825684,
23.9106025695801,
-45.4018783569336,
-11.2285804748535,
74.7284851074219,
0.221050262451172,
-16.4997920989990,
45.1744232177734,
-26.6651744842529,
-31.6537456512451,
27.5796642303467,
64.5336074829102,
24.9305267333984,
-1.15677618980408,
30.0219993591309,
49.2495651245117,
50.3987121582031,
33.2379455566406,
7.81756210327148,
3.83164262771606,
31.2497367858887,
-29.1282596588135,
35.7141990661621,
10.6351976394653,
-14.0426025390625,
34.0269165039063,
-42.1755409240723,
41.1573028564453,
-17.0575771331787,
26.5609951019287,
82.8825149536133,
0.652007102966309,
48.6309127807617,
4.80419874191284,
-8.91874122619629,
11.7633228302002,
60.5438461303711,
-16.8874111175537,
-44.6315460205078,
11.0830421447754,
-35.1148529052734,
31.9214763641357,
24.3610877990723,
19.0943698883057,
22.4307994842529,
-29.2303562164307,
-22.3531894683838,
47.2688636779785,
43.9452285766602,
-54.5573959350586,
-8.81878280639648,
41.9035110473633,
59.9008522033691,
4.95431661605835,
-11.6536979675293,
3.09588789939880,
-14.0663566589355,
37.7102661132813,
1.35333383083344,
58.2876510620117,
18.3083477020264,
-45.0411415100098,
29.7648773193359,
-18.8330688476563,
15.8916282653809,
71.1717147827148,
7.37884330749512,
-20.4628906250000,
-9.66208267211914,
12.0584163665771,
25.6461334228516,
-38.6237945556641,
-24.4010524749756,
21.1523189544678,
22.6813449859619,
52.4139175415039,
-5.74378824234009,
3.26478719711304,
-4.75128936767578,
-27.6056060791016,
52.4767379760742,
-28.2415256500244,
-22.8881092071533,
51.8085746765137,
-13.4263353347778,
8.53488826751709,
33.0520782470703,
3.06646203994751,
-24.3007335662842,
-16.4593486785889,
1.26418590545654,
19.4582214355469,
45.3047409057617,
13.0818309783936,
37.6688385009766,
36.6550445556641,
-30.5267829895020,
-12.0838499069214,
38.6985893249512,
49.0695114135742,
12.7395563125610,
-14.4417009353638,
10.1138687133789,
35.6706466674805,
25.6415214538574,
7.42472648620606,
19.0084228515625,
1.69448757171631,
-42.3084297180176,
-2.08109140396118,
59.9233665466309,
8.42197990417481,
-45.0475311279297,
55.6408386230469,
17.8229293823242,
-46.5655441284180,
53.8714256286621,
-0.976986885070801,
8.34908390045166,
30.3759574890137,
-16.0037040710449,
22.0786075592041,
-12.2300148010254,
-26.3434276580811,
-1.48890972137451,
-29.9833602905273,
-45.0599937438965,
-33.9010200500488,
-43.5348510742188,
-16.6432018280029,
-4.45583391189575,
26.2208938598633,
-7.71140146255493,
-22.3306598663330,
67.1233673095703,
6.09433126449585,
20.1948814392090,
61.8855514526367,
-11.0618438720703,
33.3856735229492,
86.2333374023438,
-0.635427713394165,
26.4902324676514,
63.8542022705078,
-21.0483379364014,
-19.1381378173828,
23.7398757934570,
12.2857112884521,
-44.8813056945801,
10.3848514556885,
12.9424667358398,
-19.8168544769287,
22.0523014068604,
-30.0398674011230,
6.46334648132324,
14.7378749847412,
-28.1031894683838,
27.9331817626953,
13.1757907867432,
10.8825397491455,
54.0735130310059,
51.0799751281738,
37.3968505859375,
0.152779102325439,
-49.8903160095215,
23.9890537261963,
41.3220481872559,
-50.5641326904297,
-25.8819961547852,
12.7216205596924,
3.19867897033691,
40.7847099304199,
23.0983467102051,
-42.9635238647461,
39.2601776123047,
43.7008590698242,
37.1797943115234,
3.54935836791992,
-15.6241455078125,
32.2249145507813,
-31.8810081481934,
32.3878021240234,
18.3848114013672,
-42.9137840270996,
-34.2431068420410,
25.4051456451416,
1.46456146240234,
-27.8098621368408,
34.8164978027344,
4.98534345626831,
-2.44018363952637,
-34.7501831054688,
-5.29145908355713,
-17.7208538055420,
15.2479705810547,
16.5918693542480,
-34.5199508666992,
10.9622697830200,
-31.0741195678711,
28.5338821411133,
47.9233665466309,
17.4692440032959,
16.2559967041016,
39.5132369995117,
54.3297920227051,
-20.5548133850098,
-10.1875286102295,
-5.15945291519165,
9.03198432922363,
-31.2919483184814,
0.346690177917480,
31.1204624176025,
-54.5244140625000,
-9.90725898742676,
-6.07193422317505,
-46.9388542175293,
-23.6682701110840,
52.3636703491211,
15.9467735290527,
46.8059654235840,
9.95975494384766,
-10.9917907714844,
23.7634906768799,
-32.0516357421875,
44.2318420410156,
-14.8293657302856,
27.6660594940186,
-14.9078693389893,
-5.67111492156982,
36.9890899658203,
-26.8123016357422,
58.5300979614258,
20.2908096313477,
-4.41240596771240,
-39.7122421264648,
9.14689445495606,
34.6738853454590,
6.77376222610474,
43.6387100219727,
45.8168067932129,
-21.5880565643311,
-2.22818565368652,
93.9407196044922,
-0.709787368774414,
0.956016540527344,
70.4733505249023,
48.9202232360840,
23.9490013122559,
3.75194549560547,
-17.3317775726318,
15.2338428497314,
27.7078037261963,
-7.94839334487915,
37.1385078430176,
39.3405685424805,
9.73926258087158,
-34.5735282897949,
4.41127777099609,
39.5509643554688,
-35.9021644592285,
27.4377231597900,
21.8468456268311,
-40.6108970642090,
-8.70353126525879,
33.2252502441406,
18.4164047241211,
-41.5274429321289,
28.6821346282959,
61.1395339965820,
19.4964981079102,
-13.8933057785034,
23.5805892944336,
44.1442909240723,
15.3705291748047,
68.7961578369141,
25.7268066406250,
-18.8504180908203,
45.4177131652832,
48.3532066345215,
-32.0891876220703,
-14.6244678497314,
58.9675254821777,
37.7311515808106,
15.3205814361572,
38.4094200134277,
18.5229492187500,
-6.71328210830689,
-1.21452939510345,
11.8048696517944,
22.9283638000488,
-27.4299259185791,
-21.9716644287109,
44.4578857421875,
6.14978742599487,
2.74151110649109,
3.81903266906738,
-9.27207183837891,
84.6298522949219,
-5.69881629943848,
-26.8342514038086,
55.8588752746582,
-46.8678054809570,
-39.6492385864258,
-17.8225765228272,
15.9555187225342,
39.1381568908691,
-41.2452812194824,
-28.3360862731934,
15.2993803024292,
3.05924987792969,
-25.5242576599121,
-29.6490058898926,
11.7049856185913,
24.7338542938232,
-35.4459915161133,
-21.8608131408691,
10.3976449966431,
29.6312160491943,
15.3327102661133,
-37.4912986755371,
46.1559753417969,
47.9421882629395,
34.3084449768066,
23.1190414428711,
8.12560176849365,
51.0820808410645,
-31.7451019287109,
31.1526241302490,
27.9533653259277,
-45.5569267272949,
-9.13327598571777,
-51.0215339660645,
-27.3229293823242,
36.5033454895020,
41.2920112609863,
14.3973312377930,
33.7247047424316,
28.8956871032715,
22.0689201354980,
35.7885169982910,
38.3776512145996,
-15.1288738250732,
-17.0898208618164,
85.7707214355469,
47.7168540954590,
29.4926948547363,
13.6308898925781,
-29.9534473419189,
50.0002593994141,
40.9499244689941,
-41.1266784667969,
37.4908065795898,
44.7881965637207,
-16.4360122680664,
11.6473751068115,
-15.0983161926270,
-1.42448806762695,
-24.4291725158691,
11.5210561752319,
20.3871231079102,
-53.4327659606934,
39.7141113281250,
-4.02239322662354,
-29.1198654174805,
48.6100120544434,
-29.1095867156982,
-39.1831436157227,
-36.5738105773926,
-36.8601150512695,
34.4678573608398,
42.6962432861328,
16.5909500122070,
-28.6667098999023,
-23.1398563385010,
11.8165988922119,
20.6366558074951,
8.22701263427734,
58.8040008544922,
5.01934242248535,
-37.1947174072266,
62.6574478149414,
-13.4445133209229,
28.8071556091309,
56.6772994995117,
31.7276592254639,
25.2645206451416,
-12.4663257598877,
46.3011016845703,
11.3803062438965,
-45.9211502075195,
-24.6502723693848,
54.3706398010254,
-40.1521263122559,
-7.56929922103882,
32.7928466796875,
-26.2083683013916,
71.7828063964844,
-32.8285064697266,
26.5625953674316,
32.1456108093262,
-36.8623886108398,
31.0166683197022,
-40.9984016418457,
39.3710975646973,
37.8122138977051,
18.9208183288574,
2.54549551010132,
-15.2141761779785,
35.4402236938477,
-25.3180141448975,
21.5452957153320,
11.6490631103516,
-11.2516269683838,
-25.6952667236328,
-17.2046833038330,
-9.36640548706055,
-37.1172332763672,
33.8791007995606,
-31.9247474670410,
-36.1186599731445,
-25.9352607727051,
-33.1910591125488,
-12.1580495834351,
2.65626144409180,
30.5509471893311,
-37.2237663269043,
39.6437873840332,
10.1086435317993,
17.0889263153076,
17.2420082092285,
-29.3627624511719,
40.9135742187500,
-33.0356407165527,
52.3839111328125,
58.2092781066895,
-8.50445747375488,
-5.04272031784058,
24.2261943817139,
20.1537189483643,
-63.4561614990234,
43.2890396118164,
44.2747993469238,
-51.2774276733398,
-12.6861848831177,
-30.9408054351807,
-12.0197563171387,
45.4163780212402,
-29.8415298461914,
-6.93763160705566,
-16.6187362670898,
2.05381870269775,
23.0139541625977,
-14.3159017562866,
51.8498382568359,
-17.2549285888672,
6.20203876495361,
33.4127311706543,
-29.3207321166992,
-3.32919836044312,
-15.0149984359741,
-16.8336067199707,
38.3176193237305,
2.85703372955322,
-43.9647445678711,
26.3930549621582,
6.39735031127930,
-21.7868881225586,
36.7589912414551,
5.43085289001465,
3.86771893501282,
55.4835319519043,
2.56191444396973,
16.4938602447510,
10.5036563873291,
-23.5556011199951,
22.8221015930176,
-26.0642185211182,
2.30916023254395,
21.7548484802246,
-16.4500255584717,
37.1874580383301,
53.2056961059570,
23.1157951354980,
3.43852949142456,
41.2998809814453,
11.7453117370605,
-22.4960231781006,
1.78368186950684,
-25.9192619323730,
-7.15712165832520,
-31.5378208160400,
-29.0125656127930,
59.4438591003418,
-6.62973833084106,
-38.6287918090820,
49.6804771423340,
-5.70657348632813,
-35.4496078491211,
49.6834716796875,
35.1991424560547,
31.7992286682129,
16.1369705200195,
8.87302398681641,
52.9109458923340,
-9.69332790374756,
-17.0280361175537,
16.1000118255615,
9.90702342987061,
21.3176822662354,
-16.0281429290772,
-4.86305475234985,
-12.5619735717773,
-46.0863304138184,
-27.7052078247070,
-10.9978752136230,
29.6742610931397,
-45.4104499816895,
-4.38236427307129,
36.0816345214844,
-57.7571601867676,
1.31620597839355,
16.0005798339844,
26.2185134887695,
48.1518135070801,
30.0971775054932,
-2.24221420288086,
6.69219350814819,
17.5066566467285,
-16.8458080291748,
43.8196411132813,
43.2188148498535,
-45.6290435791016,
25.0111579895020,
45.1161193847656,
-35.8247070312500,
28.5734729766846,
-9.37047576904297,
-12.6323442459106,
-9.80909538269043,
-12.7052707672119,
37.4333343505859,
18.8223018646240,
23.7188873291016,
-21.9280204772949,
42.4281158447266,
38.8919105529785,
-0.0496058464050293,
-12.5058631896973,
-34.9662628173828,
22.9836044311523,
-25.5721645355225,
-28.4639873504639,
41.3256187438965,
31.8037910461426,
-31.6811561584473,
-27.2767219543457,
26.8636360168457,
52.4389266967773,
-4.94940090179443,
-1.07172346115112,
65.4696960449219,
8.93780136108398,
7.47978687286377,
-39.3187713623047,
5.63259124755859,
36.4423904418945,
-57.1894950866699,
34.9943695068359,
-16.1291446685791,
-13.4775819778442,
33.8051948547363,
-23.3834457397461,
22.1311149597168,
31.0184288024902,
29.1212196350098,
5.81171226501465,
-23.4415340423584,
-21.3252887725830,
39.7728843688965,
2.29203176498413,
-40.6196975708008,
15.6563339233398,
1.30269467830658,
2.62851428985596,
17.1956329345703,
-1.68241691589355,
-29.8349533081055,
-36.7775459289551,
-34.2225189208984,
33.6902732849121,
8.94066047668457,
-10.5510864257813,
83.6522674560547,
-22.3197708129883,
-23.7545566558838,
53.2259902954102,
-51.2881011962891,
-11.0011997222900,
47.2961082458496,
11.0537958145142,
35.1753845214844,
0.200197696685791,
-41.6946945190430,
1.38725996017456,
4.91875553131104,
2.89971160888672,
67.0109100341797,
21.7984275817871,
-4.77406787872314,
69.5358734130859,
17.0870895385742,
-10.1046009063721,
14.5988092422485,
15.5969724655151,
43.3129615783691,
-17.6791458129883,
-25.5530624389648,
56.0552482604981,
5.91671371459961,
-26.8671607971191,
-10.4395637512207,
-5.19723463058472,
2.71302485466003,
-32.9780921936035,
-0.386070489883423,
51.9201049804688,
-16.0735893249512,
-50.5345993041992,
65.1207733154297,
16.1350479125977,
-32.3882293701172,
41.8539886474609,
32.7158699035645,
22.7353534698486,
-10.4106550216675,
39.8439979553223,
47.0311203002930,
54.4189338684082,
-2.09766197204590,
-15.6906366348267,
35.2957458496094,
-35.3464088439941,
8.69425296783447,
-6.73689079284668,
43.0277862548828,
36.7174682617188,
2.24901342391968,
22.3083209991455,
19.1250209808350,
42.8372611999512,
-5.42066192626953,
21.0939750671387,
20.2454204559326,
18.8475475311279,
-9.34567832946777,
51.0002288818359,
45.1840476989746,
-20.9764518737793,
57.4931602478027,
5.85666418075562,
11.0402412414551,
0.948605537414551,
18.8627243041992,
10.3870487213135,
-34.3439178466797,
44.1856651306152,
-2.70464944839478,
33.4339561462402,
-6.43335247039795,
-37.9258728027344,
8.35618495941162,
-26.7173385620117,
-3.50009226799011,
-12.8531532287598,
-13.4093189239502,
5.39047479629517,
7.77633571624756,
-47.6046600341797,
34.3876953125000,
72.0615539550781,
-17.4303607940674,
-46.7327957153320,
41.2638282775879,
41.8210983276367,
-21.7355880737305,
60.2426452636719,
-10.1876373291016,
-44.0113983154297,
-8.76082897186279,
40.9966697692871,
-16.8305206298828,
-18.4187164306641,
38.7665710449219,
-51.6292343139648,
4.48070907592773,
19.0664272308350,
25.0986042022705,
27.5778484344482,
-7.74623394012451,
47.3902587890625,
49.1472930908203,
5.27078151702881,
54.2017440795898,
33.1658287048340,
-23.4021797180176,
63.6156196594238,
16.6113967895508,
-13.8679866790771,
70.4353637695313,
22.9966430664063,
39.0726242065430,
51.2945060729981,
13.6082677841187,
55.4456710815430,
46.2638740539551,
-7.20980072021484,
-9.76392555236816,
53.9376831054688,
21.1671047210693,
21.6927680969238,
36.8711547851563,
-19.4153137207031,
34.7526855468750,
-17.1878871917725,
7.93175983428955,
73.2648925781250,
32.9361495971680,
45.2659416198731,
5.12647533416748,
8.79265022277832,
32.7777404785156,
4.53604888916016,
-38.5095596313477,
37.1947708129883,
53.7970771789551,
-29.3087425231934,
-15.5127077102661,
-10.2348842620850,
-16.7217483520508,
0.950193405151367,
33.8161849975586,
-14.8562994003296,
10.8370962142944,
14.7048273086548,
-48.2131233215332,
26.0844764709473,
6.67209243774414,
-11.3451528549194,
6.94752311706543,
10.6132316589355,
38.6074600219727,
2.13016891479492,
-12.5925025939941,
-28.5573654174805,
-2.37694740295410,
8.03195953369141,
13.1112575531006,
51.0539131164551,
25.7120323181152,
-23.2648048400879,
-23.1119480133057,
-0.977668762207031,
-2.72268295288086,
50.6936187744141,
50.5209426879883,
43.3818168640137,
5.69845867156982,
-36.2351112365723,
24.8699283599854,
34.6513023376465,
16.6899700164795,
36.0284805297852,
48.2251739501953,
6.48870134353638,
39.1423835754395,
52.6516914367676,
-33.6400413513184,
22.1059532165527,
33.6349639892578,
-43.1280326843262,
1.38159179687500,
24.0881576538086,
67.5968933105469,
9.47059822082520,
-6.62977504730225,
42.2480049133301,
-26.6829452514648,
54.5231552124023,
25.0675182342529,
-0.176129639148712,
39.9046020507813,
-40.4878921508789,
-4.30345439910889,
29.5376358032227,
-15.9537391662598,
-4.94413566589356,
38.7175750732422,
-1.77544188499451,
32.5214958190918,
59.3161888122559,
-6.15424060821533,
35.2800025939941,
12.2036323547363,
-5.60568571090698,
40.8065948486328,
55.2572860717773,
15.9868822097778,
47.1271095275879,
45.2364120483398,
-18.9786338806152,
52.5781707763672,
-0.220096826553345,
27.3119640350342,
34.9029846191406,
22.8239078521729,
33.1704406738281,
-48.7181701660156,
21.7251586914063,
-10.5268049240112,
35.0093269348145,
-0.666564941406250,
-54.4827003479004,
67.2018203735352,
-0.670614242553711,
-34.4071998596191,
-27.7207851409912,
10.1966381072998,
-16.3683509826660,
-46.9835700988770,
2.14401817321777,
22.9594669342041,
46.5915298461914,
-27.8281345367432,
13.8620681762695,
-4.69113779067993,
-1.05364418029785,
79.0726470947266,
8.09546184539795,
20.8242912292480,
47.8506164550781,
46.9380073547363,
-4.20839786529541,
30.5376434326172,
38.4871902465820,
-29.4254264831543,
33.0238533020020,
9.53599643707275,
11.2445964813232,
23.6928672790527,
9.76167297363281,
-2.17687034606934,
-40.6910552978516,
-26.6786727905273,
-35.1892471313477,
34.0795631408691,
51.3305282592773,
-18.4318408966064,
-13.0082540512085,
-5.88296651840210,
-37.0143089294434,
-8.19658374786377,
25.7029762268066,
-28.7115879058838,
-33.7669486999512,
33.3858566284180,
52.8655014038086,
-9.57608032226563,
42.9893531799316,
8.69801139831543,
-37.0400238037109,
38.7710494995117,
35.0067367553711,
46.1757698059082,
-6.83017921447754,
-23.1171703338623,
1.23937892913818,
39.0521354675293,
45.9353027343750,
5.00652456283569,
-10.2864637374878,
-37.8458061218262,
-34.3167266845703,
-35.9523429870606,
0.559070587158203,
43.9147682189941,
8.81673431396484,
-22.5521526336670,
5.94503021240234,
30.2959327697754,
34.0964355468750,
21.0528545379639,
7.45712804794312,
11.3182582855225,
46.0913925170898,
34.1084175109863,
20.1074161529541,
67.0075149536133,
-10.6011142730713,
0.919088363647461,
59.4041328430176,
24.7660713195801,
23.4125194549561,
-5.34056854248047,
45.4354896545410,
33.9383201599121,
5.14908790588379,
65.0487442016602,
58.5172729492188,
-12.1907176971436,
-28.3061790466309,
45.2224464416504,
-12.4331226348877,
-5.08529949188232,
43.5446281433106,
12.3803853988647,
-10.6722984313965,
-27.9704456329346,
59.8112945556641,
-3.19122409820557,
-7.10615539550781,
78.4850311279297,
-15.8818101882935,
-41.9408416748047,
26.8049201965332,
68.9892883300781,
29.9128341674805,
40.2283248901367,
20.9671516418457,
-35.3272895812988,
53.8951950073242,
29.3639869689941,
-16.3961429595947,
68.9847412109375,
0.681946516036987,
1.42568063735962,
48.2430915832520,
3.73453593254089,
59.8029708862305,
-15.3718490600586,
-41.5743484497070,
56.7182922363281,
-18.6742134094238,
-5.31731891632080,
11.6189479827881,
-35.3951568603516,
67.1862106323242,
8.91701316833496,
-14.9919815063477,
22.5331020355225,
-36.4238929748535,
31.1627311706543,
0.558357715606690,
26.5124015808105,
17.0783290863037,
-65.2401199340820,
35.8839950561523,
35.9206314086914,
52.1187248229981,
13.1430454254150,
-6.72651958465576,
6.53946018218994,
-6.48669338226318,
68.7490463256836,
-7.39745712280273,
-28.4581413269043,
-1.51850390434265,
53.0550994873047,
5.86784458160400,
28.0084648132324,
32.7883300781250,
-38.5117111206055,
58.6123390197754,
-39.5493240356445,
31.3806953430176,
27.4668674468994,
-53.1909103393555,
44.2191467285156,
16.3746166229248,
-25.8053016662598,
-3.99779891967773,
47.3226928710938,
7.91476535797119,
-22.5335521697998,
-27.9675464630127,
23.9700393676758,
-5.10155248641968,
-27.3765144348145,
34.6436729431152,
-14.4234886169434,
27.5869560241699,
-16.1134624481201,
-22.3764610290527,
74.2950820922852,
9.55790805816650,
20.4153118133545,
49.2782516479492,
-13.2509088516235,
-27.7368011474609,
45.5941505432129,
32.8955192565918,
-3.55688023567200,
15.9986057281494,
17.1735877990723,
3.64660310745239,
9.65944480895996,
48.9840965270996,
-0.303276538848877,
36.6923522949219,
16.2793960571289,
-51.4734802246094,
23.4733867645264,
52.2272224426270,
24.3415660858154,
-59.5544281005859,
16.9514846801758,
63.4017944335938,
-43.3391723632813,
11.0401058197021,
-7.63754034042358,
-53.1227722167969,
8.96214580535889,
-14.3307485580444,
-3.89960384368897,
62.2878913879395,
16.4153633117676,
24.4921455383301,
35.3108596801758,
-8.65531539916992,
43.1780776977539,
19.1292381286621,
38.7909774780273,
9.63329601287842,
-49.1624374389648,
12.6399040222168,
-28.8926029205322,
5.78558588027954,
-6.56059074401856,
-36.4224090576172,
-26.2398376464844,
-49.9756927490234,
39.8974037170410,
20.0138206481934,
37.5929756164551,
2.55577898025513,
-46.2115516662598,
58.4708251953125,
-12.2441425323486,
-23.8547191619873,
29.8682670593262,
-4.35075092315674,
-13.7161035537720,
1.57400989532471,
41.7677650451660,
22.1876525878906,
-33.5084686279297,
-5.45807838439941,
-1.20670604705811,
-51.5747947692871,
2.07226181030273,
0.958442687988281,
-39.6073455810547,
13.0883769989014,
16.3686561584473,
-26.7634124755859,
-29.2357921600342,
42.7832794189453,
42.9316329956055,
-2.87229347229004,
-1.96754026412964,
-33.0975723266602,
3.92315292358398,
51.1563568115234,
46.3062477111816,
15.0648145675659,
-17.0414123535156,
-20.7484607696533,
-5.61027526855469,
43.5716438293457,
41.2575073242188,
8.13238716125488,
-5.23770141601563,
23.4465847015381,
1.54947948455811,
-23.9052238464355,
60.6476554870606,
1.97566080093384,
-63.2581367492676,
29.4439754486084,
46.1890068054199,
31.0562286376953,
14.3044147491455,
47.6570472717285,
42.7421340942383,
-49.0473976135254,
37.8936500549316,
79.2672805786133,
8.11417007446289,
3.06665396690369,
-22.9352855682373,
-27.6915893554688,
10.4781360626221,
28.1136398315430,
1.66779518127441,
-42.5520744323731,
-34.5336227416992,
-18.9881858825684,
37.3935394287109,
33.3348045349121,
-45.8430099487305,
-3.79301166534424,
-0.583800315856934,
23.2153759002686,
16.5764522552490,
-5.19871425628662,
34.9315490722656,
-23.1686401367188,
46.1027526855469,
48.9019508361816,
18.3416233062744,
56.9624214172363,
-9.03030776977539,
25.1844329833984,
21.6901435852051,
10.2911977767944,
10.8108501434326,
-28.4327487945557,
64.6276016235352,
43.9088859558106,
-48.3801956176758,
46.8867073059082,
48.0876731872559,
-24.2247676849365,
38.0593566894531,
64.9973907470703,
34.8822326660156,
-0.871964454650879,
2.47253966331482,
7.67946290969849,
-11.1236190795898,
43.4503593444824,
49.1222190856934,
-9.35067844390869,
-16.6777801513672,
-20.2659587860107,
-4.24927234649658,
0.0512204170227051,
17.3743782043457,
34.4693298339844,
12.7329349517822,
-8.24698448181152,
-3.01785612106323,
28.7349319458008,
-16.6474895477295,
32.8745765686035,
44.6197509765625,
9.22344970703125,
69.1224441528320,
1.76472091674805,
28.5524253845215,
33.9312210083008,
27.1539802551270,
30.5118503570557,
-35.1748313903809,
62.0358123779297,
23.6890525817871,
27.6632843017578,
11.8351030349731,
-20.6472415924072,
27.1541099548340,
3.30979394912720,
0.204575538635254,
-18.8036708831787,
22.9318141937256,
-39.7635231018066,
34.3872604370117,
21.9177055358887,
3.73379421234131,
43.5245819091797,
-16.6789207458496,
33.1516189575195,
-32.8514328002930,
23.9300308227539,
51.5294647216797,
45.8805236816406,
-17.8892211914063,
-19.8186035156250,
40.1836624145508,
-27.6785583496094,
68.3150100708008,
-3.44859313964844,
-33.2994537353516,
41.6813278198242,
-26.2436618804932,
-21.7440338134766,
-3.25857639312744,
-1.52920520305634,
-48.5856933593750,
0.522900581359863,
77.0061492919922,
19.4359130859375,
34.9065513610840,
12.0451507568359,
14.4452476501465,
45.0512924194336,
-7.35769462585449,
-26.2838573455811,
16.2066612243652,
69.3776626586914,
-23.5424690246582,
3.93860244750977,
76.8784179687500,
-4.43324470520020,
-17.5776596069336,
49.6587944030762,
55.1207122802734,
5.33726501464844,
27.1505374908447,
20.1135368347168,
45.9379043579102,
13.9799156188965,
14.1104946136475,
35.7953414916992,
21.3593254089355,
45.8815231323242,
-32.7457809448242,
21.5654735565186,
4.97779560089111,
23.4215965270996,
76.4994049072266,
-39.4774856567383,
17.9805374145508,
62.5997390747070,
26.2072868347168,
38.2969169616699,
66.1519622802734,
44.8098831176758,
-43.1791687011719,
-5.94615554809570,
66.1038360595703,
19.8758563995361,
23.7209300994873,
9.87470817565918,
-57.7822837829590,
41.7881317138672,
25.7405300140381,
-26.2827243804932,
23.4365005493164,
-46.5643157958984,
-1.21471214294434,
33.7807998657227,
-1.02219414710999,
18.8733577728272,
49.5163536071777,
-9.72574996948242,
-7.33913421630859,
34.9441223144531,
-46.5676956176758,
30.2170791625977,
57.3119392395020,
22.4771804809570,
15.8106451034546,
-32.7629165649414,
-21.8309974670410,
-30.7730045318604,
-13.0020246505737,
30.4108695983887,
3.37870788574219,
4.49949550628662,
32.5881576538086,
-27.5247859954834,
-4.74233818054199,
53.4114570617676,
11.2422256469727,
18.6267795562744,
26.0024967193604,
46.4288291931152,
47.3067131042481,
19.3244285583496,
20.6542854309082,
-29.6947383880615,
45.7771530151367,
48.4887199401856,
-23.5103111267090,
25.6054286956787,
-9.57889747619629,
16.2183055877686,
21.2408981323242,
-2.10682868957520,
77.5455627441406,
22.5562343597412,
-20.2173309326172,
29.2258872985840,
3.56586265563965,
-11.8081073760986,
13.0129661560059,
-1.49704015254974,
-4.70432710647583,
62.5607604980469,
1.67226409912109,
-41.8281936645508,
73.6653137207031,
15.5016899108887,
-22.7378997802734,
59.8064918518066,
8.93882369995117,
15.0858221054077,
16.6161289215088,
-36.1501922607422,
34.9408454895020,
53.9628906250000,
18.5223026275635,
25.1781463623047,
-14.8132781982422,
-16.2905235290527,
35.9323921203613,
-12.3225660324097,
-30.9139118194580,
28.7871360778809,
6.69270610809326,
-16.5169181823730,
25.8364219665527,
64.9354629516602,
30.6333522796631,
-7.22512340545654,
44.3883972167969,
65.6358642578125,
-11.2412471771240,
-14.8284568786621,
54.4116096496582,
-8.96797752380371,
-2.59150624275208,
41.3674087524414,
-0.533206939697266,
-31.0625000000000,
-18.0252780914307,
47.6906089782715,
-25.3412170410156,
-38.4693756103516,
-3.90723514556885,
-33.2929191589356,
6.22623729705811,
1.06069147586823,
-9.95345306396484,
16.1630249023438,
-17.7309722900391,
-21.1461219787598,
12.3602428436279,
-16.4009552001953,
-13.0715255737305,
18.5338745117188,
32.0844001770020,
-3.68469715118408,
24.0960426330566,
34.9193687438965,
-38.6449203491211,
-37.5645294189453,
11.6627368927002,
38.6841812133789,
-4.13636207580566,
29.1156997680664,
56.2090682983398,
16.1100616455078,
21.8883686065674,
43.5481834411621,
61.7974967956543,
9.07717323303223,
-43.1156845092773,
7.31922245025635,
22.9220886230469,
19.1467800140381,
20.3458404541016,
-29.0853557586670,
26.3978023529053,
17.8528385162354,
-28.8001384735107,
48.6037635803223,
49.7818489074707,
18.3345184326172,
-21.4909477233887,
7.84826660156250,
59.8901481628418,
-33.1635284423828,
-46.3471755981445,
20.4321899414063,
25.3193912506104,
27.1786079406738,
14.8709497451782,
50.0759658813477,
46.3501319885254,
-22.5943546295166,
-2.93515825271606,
-9.08122634887695,
2.26440668106079,
-0.315131425857544,
-48.9308090209961,
17.1978073120117,
27.7306270599365,
4.15889596939087,
33.1488075256348,
-7.75908613204956,
63.7675514221191,
41.6003494262695,
-55.4131698608398,
65.4773406982422,
33.8892364501953,
23.3280067443848,
53.5403594970703,
-37.6673851013184,
-0.533667325973511,
-15.9626512527466,
-34.2882385253906,
11.5890445709229,
-37.4827461242676,
-43.9777717590332,
17.5938034057617,
-26.8719253540039,
-55.3641586303711,
19.2664375305176,
23.7092971801758,
21.6354122161865,
4.82086944580078,
-14.8453073501587,
6.80096673965454,
25.5713920593262,
27.1357021331787,
-32.8022575378418,
35.2863121032715,
38.0516052246094,
-50.4696235656738,
-18.9417533874512,
-13.7400531768799,
-2.97347140312195,
-34.5056800842285,
8.77089500427246,
29.4137401580811,
-15.7309131622314,
10.6571607589722,
7.21659374237061,
47.6520957946777,
-23.0806961059570,
21.1601791381836,
45.7514495849609,
-14.6521511077881,
73.6640090942383,
2.75685310363770,
-2.58855295181274,
-22.6940383911133,
-49.0958938598633,
48.0249748229981,
48.7406425476074,
-8.18308353424072,
20.7229080200195,
52.3411254882813,
-9.76980209350586,
61.0013694763184,
45.9532737731934,
-12.9173870086670,
51.9469146728516,
9.14140510559082,
-24.1873321533203,
7.84670591354370,
35.8592414855957,
54.8289031982422,
25.6780414581299,
1.33589935302734,
18.1425476074219,
12.1612405776978,
3.18468189239502,
-17.6719970703125,
-30.1687488555908,
-9.25534820556641,
-45.5513534545898,
-4.46217775344849,
1.55977189540863,
-14.1685981750488,
43.0673217773438,
8.19922924041748,
52.9846076965332,
41.1153564453125,
-18.3104648590088,
-12.7585115432739,
-17.7081069946289,
1.72345685958862,
-32.6528854370117,
-20.6818428039551,
33.4272460937500,
44.9749031066895,
-5.63909149169922,
-24.0101184844971,
13.2659120559692,
25.0292968750000,
36.5051612854004,
-20.0486679077148,
4.22525978088379,
38.3140602111816,
10.8768291473389,
20.6021137237549,
6.16461658477783,
8.56363010406494,
6.99049854278564,
52.2879638671875,
-8.72557830810547,
-22.8862476348877,
75.7036132812500,
-19.5157508850098,
-1.85667443275452,
22.4632396697998,
-59.4430389404297,
8.49427413940430,
-2.86550140380859,
-33.3041458129883,
43.7227630615234,
35.8826637268066,
5.58998203277588,
20.5990867614746,
28.5934219360352,
-7.55905342102051,
-43.8796157836914,
-15.5352325439453,
18.0954723358154,
30.5836334228516,
-20.7677230834961,
9.05750274658203,
55.0445365905762,
-2.00533986091614,
37.2473793029785,
34.0620040893555,
37.4505577087402,
19.7226982116699,
34.6929473876953,
39.1859626770020,
-21.0328292846680,
59.8901748657227,
29.3202247619629,
-22.9035720825195,
6.74755811691284,
46.9987945556641,
21.6068134307861,
-12.3127994537354,
-25.2152767181397,
-14.5038242340088,
-33.0948867797852,
-15.1754570007324,
53.3630371093750,
-30.0449333190918,
26.1226711273193,
-27.7258758544922,
-0.104113578796387,
72.5097808837891,
-67.6374435424805,
32.4507904052734,
36.0399742126465,
11.7181606292725,
42.4294586181641,
-18.6075286865234,
54.3204803466797,
43.4607124328613,
-2.03293943405151,
57.8018646240234,
64.8224945068359,
25.7236289978027,
23.5465183258057,
36.3917198181152,
11.3267660140991,
40.0915336608887,
55.0242271423340,
48.0543327331543,
15.4767704010010,
-18.4594707489014,
2.69425487518311,
-33.5557289123535,
21.8944797515869,
80.8610687255859,
11.0348320007324,
7.44283103942871,
20.9191894531250,
-9.52897644042969,
43.3842811584473,
60.3402481079102,
28.0881919860840,
50.5491714477539,
-6.67421627044678,
26.8058300018311,
30.9402389526367,
7.67501497268677,
48.6838417053223,
-33.6371383666992,
-12.3405351638794,
17.2394199371338,
46.5985565185547,
47.2346839904785,
-41.9025077819824,
-2.21247863769531,
59.8582687377930,
14.9391765594482,
-31.9985237121582,
-14.7126979827881,
-7.43136453628540,
-20.4928169250488,
6.17703151702881,
-8.63527488708496,
-21.9726867675781,
10.0019588470459,
-17.0531921386719,
27.3383159637451,
-24.4564037322998,
-7.44286537170410,
54.4843444824219,
-25.4399261474609,
6.78189182281494,
5.47746133804321,
23.0752525329590,
34.7367362976074,
29.7744178771973,
37.7151374816895,
33.4743309020996,
54.1998252868652,
45.2409820556641,
40.2655258178711,
51.1916961669922,
40.7567863464356,
-24.2326145172119,
10.7055892944336,
11.2594041824341,
-15.2210206985474,
-5.33771848678589,
-49.5898742675781,
22.3686218261719,
-8.51998233795166,
-39.3272895812988,
33.3188934326172,
31.4926700592041,
11.7051486968994,
3.82144021987915,
57.6180305480957,
25.0950088500977,
7.62207555770874,
-10.5859336853027,
-8.07970142364502,
47.1950416564941,
27.3739929199219,
19.7235050201416,
14.2146234512329,
6.04112911224365,
30.0570507049561,
45.2106781005859,
-34.8210182189941,
16.5922508239746,
56.1454887390137,
-17.7794513702393,
10.1549520492554,
20.5448188781738,
-7.13297843933106,
-7.77843284606934,
62.1733016967773,
44.8940315246582,
-13.7993583679199,
44.9208984375000,
19.4767799377441,
-28.7644863128662,
34.8604583740234,
48.3585433959961,
31.6624507904053,
30.4820919036865,
49.0098114013672,
49.0822067260742,
-25.9302635192871,
20.2956657409668,
47.5577697753906,
5.96700429916382,
28.1724243164063,
9.35272884368897,
17.9223022460938,
31.4364700317383,
-6.25086021423340,
-13.5614595413208,
-28.4071369171143,
-17.8644142150879,
19.7705230712891,
-38.9437561035156,
-16.5417709350586,
37.8118667602539,
33.3944816589356,
34.4367027282715,
-6.56452131271362,
-13.9455785751343,
35.7527656555176,
52.2748870849609,
37.2673492431641,
48.1128578186035,
-1.12750256061554,
32.2610244750977,
65.4748916625977,
-17.9730758666992,
9.33943843841553,
64.9568328857422,
-1.76871490478516,
18.5973072052002,
60.4836387634277,
-23.0378704071045,
-33.9794769287109,
19.1989936828613,
55.9334182739258,
11.2149724960327,
9.52898597717285,
-11.1970605850220,
19.8074054718018,
40.2613105773926,
0.713790893554688,
12.0478134155273,
-26.3844928741455,
44.0466461181641,
-1.92913842201233,
9.38090515136719,
13.4370822906494,
-7.98223066329956,
62.3053970336914,
-24.4466533660889,
7.98552322387695,
35.5461845397949,
38.1460075378418,
-6.14835596084595,
0.720708847045898,
64.4953384399414,
-3.80755424499512,
-22.1567802429199,
-10.7548952102661,
69.1312561035156,
7.64360427856445,
-46.5342636108398,
37.0795288085938,
-41.9292716979981,
-46.1109886169434,
-18.2028255462647,
3.72073268890381,
24.4167671203613,
11.2185363769531,
48.6458244323731,
-56.8924942016602,
20.0494308471680,
51.4258804321289,
-53.5691223144531,
8.80028152465820,
-22.9145164489746,
36.2123603820801,
-16.7173500061035,
-72.8107681274414,
48.2020645141602,
45.0084571838379,
-3.13679003715515,
-1.44803905487061,
48.7907638549805,
1.69333839416504,
-25.9486522674561,
59.8269729614258,
63.5102310180664,
3.18497252464294,
8.81231975555420,
-12.5652332305908,
0.251135826110840,
71.2254486083984,
8.62833404541016,
-47.8955612182617,
46.4870376586914,
45.2842407226563,
-23.6344184875488,
60.4536476135254,
7.55669307708740,
-49.5965995788574,
23.5517444610596,
3.04586696624756,
0.582013130187988,
-11.9522123336792,
-17.4087009429932,
-12.3342952728271,
-44.9684028625488,
-18.1937103271484,
34.5323028564453,
41.6575202941895,
19.9231243133545,
52.1273422241211,
19.7898960113525,
-18.7834129333496,
54.3028030395508,
-1.38719558715820,
-16.4626998901367,
34.3833007812500,
36.9589118957520,
34.3630332946777,
-36.3588142395020,
12.4548959732056,
37.5838012695313,
24.2159271240234,
28.0724334716797,
49.7440986633301,
38.5549354553223,
13.0324192047119,
55.1488075256348,
14.8054084777832,
16.7205829620361,
-15.6214637756348,
-1.21651518344879,
12.8792018890381,
11.8781490325928,
0.816776514053345,
22.3003158569336,
41.5918579101563,
-31.5605697631836,
-13.1562404632568,
-24.5460472106934,
22.1162071228027,
-24.2969570159912,
14.3803138732910,
57.1918067932129,
-15.2304325103760,
48.1153221130371,
52.8393592834473,
-6.03092575073242,
-23.0815544128418,
45.3726539611816,
-23.9899330139160,
-19.8722076416016,
64.3046340942383,
-0.643688082695007,
0.790420532226563,
16.6712703704834,
26.9468097686768,
54.7408599853516,
37.6770401000977,
41.0112686157227,
16.1822414398193,
1.59670925140381,
67.4060592651367,
12.3814001083374,
-20.8781547546387,
8.51226615905762,
-27.1057891845703,
2.82887554168701,
34.1047744750977,
46.8371276855469,
4.33054351806641,
-7.34173774719238,
27.6808147430420,
-29.1390514373779,
18.5457496643066,
64.5800704956055,
-12.8270788192749,
-26.2596530914307,
13.6186962127686,
27.9282264709473,
34.6405029296875,
43.0665359497070,
32.1056938171387,
-27.1194114685059,
-10.5035505294800,
13.9365053176880,
-29.9217681884766,
40.5666923522949,
-13.5811233520508,
-30.1842460632324,
39.4906349182129,
-12.4369983673096,
0.373558044433594,
1.54225361347198,
-11.0389785766602,
-6.93689441680908,
50.5693092346191,
15.6415843963623,
22.3673248291016,
58.4242095947266,
-36.3664665222168,
6.63181495666504,
54.9495849609375,
19.0369186401367,
-26.1319751739502,
14.1247482299805,
19.9955921173096,
-32.0605506896973,
-10.4795398712158,
-4.43298244476318,
0.753297090530396,
-19.3851814270020,
-31.1235198974609,
8.46734809875488,
24.2503452301025,
47.0099983215332,
35.2432441711426,
24.4219245910645,
59.6844329833984,
-12.9309062957764,
-36.2045593261719,
-13.9404067993164,
-18.3140983581543,
-4.33967447280884,
18.0619487762451,
16.5977401733398,
-44.8924407958984,
-21.5653514862061,
-22.2863864898682,
21.1209468841553,
64.8028106689453,
-40.5141830444336,
-20.4498863220215,
63.1729583740234,
42.3414459228516,
35.1717071533203,
25.4271087646484,
35.9440917968750,
58.4797897338867,
-2.31940460205078,
47.0938224792481,
30.6533241271973,
-58.0104598999023,
31.7671222686768,
48.0825729370117,
34.4581451416016,
30.8587551116943,
-2.00681400299072,
28.2301712036133,
-37.3719024658203,
-19.4748611450195,
19.6563282012939,
-42.8699340820313,
31.0763530731201,
-0.400282859802246,
-29.2956619262695,
-30.2614860534668,
-12.8242130279541,
51.0061569213867,
-34.3359603881836,
-5.11381340026856,
30.7993736267090,
23.8842468261719,
-20.8206863403320,
-43.1398925781250,
-12.2732028961182,
-5.46668243408203,
60.2907028198242,
21.8279933929443,
-35.3565826416016,
-8.52018165588379,
56.7227973937988,
2.11518287658691,
-6.84371757507324,
59.9753684997559,
-25.8851718902588,
-24.6054687500000,
-4.75694942474365,
12.4616079330444,
48.4847602844238,
-36.7909469604492,
17.1217842102051,
61.1040344238281,
-13.2678041458130,
31.5485572814941,
59.4675331115723,
14.2594614028931,
-53.9258956909180,
27.6509990692139,
49.6670227050781,
-40.1248130798340,
12.9426460266113,
-5.60318565368652,
-44.7949676513672,
14.0106077194214,
50.7911109924316,
-23.6436119079590,
-43.7131462097168,
-16.3830471038818,
9.68836116790772,
4.61610174179077,
-1.82843589782715,
31.2740745544434,
-17.6219749450684,
-1.27095079421997,
-0.870524883270264,
3.92289447784424,
45.4055480957031,
-6.83769893646240,
-64.5386199951172,
28.2682323455811,
32.6269493103027,
-31.2061614990234,
42.8224334716797,
28.5641784667969,
36.4683303833008,
-33.1523094177246,
17.0104770660400,
89.7084655761719,
5.53977537155151,
45.1025581359863,
-7.23501110076904,
9.73323631286621,
9.32654190063477,
-9.20322608947754,
62.6094818115234,
35.1121673583984,
25.5534286499023,
-11.7612142562866,
-15.3009119033813,
3.47292637825012,
13.6887998580933,
21.8985748291016,
-15.1437911987305,
19.8866081237793,
20.1019897460938,
14.1710872650146,
25.6430988311768,
29.4088020324707,
32.0494155883789,
12.6431694030762,
50.0945854187012,
15.3199234008789,
-24.1702861785889,
-9.22607421875000,
-18.2305278778076,
10.4229707717896,
34.2457389831543,
35.6874885559082,
-7.93816471099854,
13.2348337173462,
55.0933456420898,
-50.1545639038086,
16.9544601440430,
59.8516311645508,
-27.7868289947510,
-6.27330017089844,
36.3143234252930,
52.8370056152344,
24.1107769012451,
49.8989868164063,
24.3773727416992,
27.7770786285400,
22.7855587005615,
-19.4696826934814,
7.63687896728516,
47.4289245605469,
24.3563632965088,
-4.42355537414551,
47.7600784301758,
-11.2809762954712,
-17.8680381774902,
21.1292037963867,
26.7950725555420,
-0.0148687362670898,
-21.9323062896729,
-0.946601867675781,
-29.0047779083252,
27.1504497528076,
42.8161621093750,
-31.3707447052002,
-42.5607872009277,
31.4789600372314,
9.84222698211670,
-52.8885345458984,
-1.08956718444824,
-1.52236139774323,
-7.24215459823608,
-17.5236968994141,
8.08820533752441,
52.6900329589844,
22.1002349853516,
6.30830335617065,
-22.4058551788330,
38.7581596374512,
70.9670028686523,
-27.0572948455811,
-22.1603507995605,
13.2746496200562,
-35.4878616333008,
-42.2080116271973,
12.9644546508789,
-0.368837118148804,
13.0887985229492,
39.5213050842285,
-10.6263542175293,
-41.5314407348633,
1.05742740631104,
41.5352554321289,
-11.0012331008911,
63.9918136596680,
34.4432296752930,
-49.9410514831543,
12.7983951568604,
26.0188789367676,
55.6607017517090,
8.92905807495117,
32.1962966918945,
-5.69888210296631,
0.223193168640137,
27.5475769042969,
-20.3449859619141,
29.5493125915527,
-5.47372150421143,
-5.53629875183106,
-21.3097724914551,
26.4076728820801,
15.4219551086426,
4.18757009506226,
50.3021697998047,
-0.614621162414551,
-10.8132801055908,
15.4531002044678,
57.0082397460938,
-12.9575462341309,
-17.9012603759766,
-9.92193698883057,
-41.6474914550781,
-11.8658237457275,
17.6610126495361,
22.0139884948730,
-27.1131649017334,
41.4175605773926,
9.79935646057129,
-50.4512786865234,
39.4364318847656,
24.8463859558105,
30.7059478759766,
1.96633672714233,
-29.3412132263184,
31.8031311035156,
23.9666500091553,
6.63282299041748,
0.0667052268981934,
-9.71616077423096,
-10.2858667373657,
-12.8643989562988,
-6.89707851409912,
46.3849334716797,
-3.89079713821411,
-65.1452789306641,
17.7541465759277,
47.4974517822266,
14.5437364578247,
-40.5023422241211,
23.6343460083008,
-1.19586753845215,
-16.6992340087891,
66.7268142700195,
-0.105172634124756,
27.9368782043457,
-17.8789367675781,
26.3393650054932,
46.2816162109375,
-4.85692691802979,
25.5230636596680,
-52.9320411682129,
44.3249816894531,
48.5656127929688,
10.1917400360107,
56.5428009033203,
51.6674118041992,
39.3551445007324,
-35.1736984252930,
20.6932334899902,
83.7960968017578,
-0.920650482177734,
-45.4403610229492,
38.9673233032227,
-3.14798927307129,
-19.9765529632568,
67.4660644531250,
4.62960624694824,
44.4509811401367,
8.37374210357666,
-9.55284118652344,
56.0351867675781,
16.7075595855713,
13.3410024642944,
-47.6831169128418,
-21.6381969451904,
-25.0524711608887,
14.8759737014771,
59.9318275451660,
-6.50629854202271,
51.4321670532227,
1.29604578018188,
2.14540672302246,
60.8994369506836,
25.5320777893066,
42.8450164794922,
-18.1449146270752,
64.4693832397461,
48.3552856445313,
-45.2170181274414,
50.8313827514648,
4.51039028167725,
44.0586433410645,
-4.59625339508057,
2.16967868804932,
43.1574363708496,
-21.5142478942871,
57.9124374389648,
-13.1037731170654,
26.9406661987305,
16.7466945648193,
-4.67778873443604,
67.6291046142578,
-14.6488714218140,
-30.3772392272949,
-14.1897792816162,
65.8403091430664,
25.4549655914307,
-26.6413116455078,
-18.7019309997559,
-26.3598651885986,
-0.502101182937622,
-29.7952995300293,
45.2867279052734,
-9.33099937438965,
-60.6916198730469,
-22.1994380950928,
-2.31771659851074,
39.2553749084473,
22.4599895477295,
1.32079982757568,
-45.4733505249023,
55.0906333923340,
46.1888656616211,
25.5939655303955,
43.9823455810547,
-44.7155342102051,
38.1918792724609,
4.88164901733398,
-38.3626861572266,
-2.65673470497131,
-37.4178848266602,
-31.1928138732910,
12.8703403472900,
51.3299140930176,
-13.6000738143921,
-54.6145820617676,
2.56269836425781,
23.4485473632813,
13.3033456802368,
-20.2562599182129,
7.38021183013916,
44.3540649414063,
-4.58274888992310,
-16.8650970458984,
12.1286716461182,
24.5762958526611,
-25.6516723632813,
-20.8505096435547,
-6.45365619659424,
33.6429443359375,
30.2050170898438,
-28.0915832519531,
6.12241935729981,
18.4206428527832,
50.6282501220703,
-24.3262901306152,
-47.6710090637207,
5.62451744079590,
-2.91339850425720,
-5.40395069122314,
14.0161056518555,
33.2813568115234,
-37.4309158325195,
-22.3154277801514,
-2.92964887619019,
-11.9683713912964,
-19.7580509185791,
8.56958389282227,
2.78009271621704,
-32.8553543090820,
20.6683311462402,
-22.5523109436035,
11.8331089019775,
0.204375267028809,
-33.1499404907227,
36.0869827270508,
-27.9390106201172,
9.43754386901856,
31.7575397491455,
-12.9493770599365,
16.3569946289063,
35.1292228698731,
21.3460826873779,
-1.47469472885132,
35.2901191711426,
-17.8859348297119,
-6.86169052124023,
60.9084205627441,
26.4994487762451,
24.4585647583008,
25.7729206085205,
8.94201755523682,
21.6203250885010,
25.5111007690430,
25.5891666412354,
12.6233310699463,
22.1575908660889,
26.4849052429199,
-34.1236457824707,
3.03052067756653,
2.86770248413086,
7.71129322052002,
2.95969963073730,
-8.69814586639404,
72.9798126220703,
12.4766254425049,
-3.37984752655029,
16.1162910461426,
-33.5208663940430,
-21.4035034179688,
8.26937484741211,
-0.669481992721558,
-21.7734794616699,
20.5299186706543,
45.4091606140137,
-4.31701660156250,
-26.7479972839355,
23.4671936035156,
5.82605838775635,
4.64036655426025,
-18.1833496093750,
-56.1421127319336,
52.3710479736328,
-11.5857009887695,
-12.6856994628906,
28.4192943572998,
-2.04249286651611,
47.9259109497070,
-51.5759887695313,
10.6550931930542,
36.2142944335938,
-42.2069854736328,
10.1211328506470,
-0.871856987476349,
17.9006080627441,
-12.3479614257813,
3.69496726989746,
16.5994415283203,
-26.5083484649658,
35.7858390808106,
23.6368732452393,
-5.51133394241333,
24.2238769531250,
-4.37109851837158,
-42.6640586853027,
17.2476367950439,
25.4231491088867,
22.3202590942383,
22.1073474884033,
-0.596682071685791,
36.7612686157227,
35.2984390258789,
44.9178657531738,
-8.05918312072754,
-37.6794929504395,
21.4147167205811,
50.7990760803223,
-12.5712451934814,
-9.68972301483154,
39.2510910034180,
-13.7465896606445,
26.0767364501953,
-15.9606552124023,
-4.12428569793701,
69.0596237182617,
-46.2055892944336,
13.0485868453980,
90.4702377319336,
5.28845214843750,
18.8170089721680,
16.5798301696777,
7.71073389053345,
6.92190742492676,
20.5362739562988,
19.3327198028564,
-26.2087917327881,
40.4548568725586,
18.8405780792236,
7.60119962692261,
-13.9794158935547,
-7.78939914703369,
59.9610061645508,
-67.7059173583984,
10.7866363525391,
54.5120353698731,
-35.9146003723145,
51.1077346801758,
40.4336013793945,
21.2638626098633,
24.4406051635742,
26.8323383331299,
19.6611976623535,
-52.6443519592285,
12.9173793792725,
49.2652778625488,
-54.7791709899902,
-23.0933227539063,
53.6349220275879,
15.6833591461182,
-38.0546035766602,
11.5153045654297,
61.8394393920898,
27.3506622314453,
33.5459899902344,
13.0270023345947,
24.8259887695313,
-3.34717845916748,
-34.9949378967285,
63.7915840148926,
21.2858772277832,
8.07678318023682,
11.5309085845947,
2.51036834716797,
47.4639434814453,
38.5038490295410,
22.3041191101074,
-20.2915134429932,
50.5293807983398,
39.4152679443359,
-43.8540458679199,
17.7397689819336,
44.4931907653809,
-2.07839012145996,
-7.03676891326904,
-13.6494846343994,
3.02548027038574,
38.0289764404297,
-19.8041210174561,
-3.77928256988525,
27.5566692352295,
-29.1081924438477,
-15.0800027847290,
50.1724929809570,
24.2807369232178,
21.6222057342529,
42.3683586120606,
-21.5925827026367,
-26.1347351074219,
-17.3976745605469,
14.3858089447021,
-16.0663604736328,
-40.4210624694824,
36.3077545166016,
-41.0885467529297,
-11.7576045989990,
36.1175003051758,
-27.0475616455078,
-55.9970054626465,
-5.45334434509277,
37.8596420288086,
-52.8236045837402,
25.6489181518555,
12.9811773300171,
-50.4881095886231,
9.99714946746826,
20.9775390625000,
54.3441009521484,
33.1613159179688,
13.1149997711182,
3.25841474533081,
2.33563661575317,
38.8307075500488,
23.7870883941650,
-9.89874839782715,
-17.2349643707275,
-42.5037727355957,
4.66424846649170,
15.7283535003662,
-5.03549909591675,
9.74240875244141,
34.3867950439453,
42.0137672424316,
-46.0738372802734,
-13.5811634063721,
-8.75077819824219,
-54.9420089721680,
-19.8068542480469,
30.9462966918945,
44.0370483398438,
17.7360420227051,
59.8349914550781,
9.02443313598633,
-33.1365928649902,
68.3200378417969,
20.6285953521729,
-21.4454727172852,
60.9352035522461,
-6.61354541778564,
5.76613855361939,
38.2047882080078,
-14.7270193099976,
13.1807632446289,
-3.94426107406616,
-13.9983148574829,
12.4888162612915,
35.2124023437500,
17.6948051452637,
-29.4611129760742,
25.1126480102539,
85.6463012695313,
-39.9007835388184,
-0.262851715087891,
57.6186523437500,
-60.1067237854004,
26.2975616455078,
40.0309906005859,
-14.0443801879883,
-31.6512889862061,
15.5148344039917,
55.1586685180664,
-20.5638084411621,
37.0485496520996,
8.00028991699219,
-33.6420822143555,
8.46243286132813,
19.6298179626465,
58.4064826965332,
17.7355060577393,
-1.95026230812073,
34.2515602111816,
13.8913688659668,
-11.5368986129761,
15.7461681365967,
16.1130542755127,
34.4843444824219,
26.8025360107422,
-13.7339534759521,
67.1436538696289,
42.8905143737793,
31.1430969238281,
35.7050704956055,
-17.5756855010986,
25.2988433837891,
6.19832611083984,
19.3864879608154,
5.87014484405518,
-25.0603790283203,
27.8978691101074,
17.9420852661133,
-46.6790199279785,
-11.3599281311035,
56.1499099731445,
-4.80255365371704,
31.4393234252930,
33.8153762817383,
-22.4485511779785,
56.9305381774902,
34.9848709106445,
-15.1166229248047,
54.2557487487793,
56.6421318054199,
32.4877204895020,
11.7625398635864,
-36.1515502929688,
20.5304126739502,
-5.67723083496094,
16.9972934722900,
4.60546875000000,
-13.8702096939087,
36.1545104980469,
-42.1888236999512,
47.0970039367676,
-19.8888359069824,
9.98881149291992,
84.8599700927734,
-54.3457565307617,
29.3026199340820,
55.5097503662109,
3.97153282165527,
-35.4999618530273,
-2.48853111267090,
55.1644897460938,
30.2265586853027,
-38.2424163818359,
12.2034282684326,
75.6660156250000,
-41.6661224365234,
38.7509918212891,
22.9113197326660,
-34.2728729248047,
80.8408660888672,
43.2247200012207,
44.6922149658203,
-18.9814796447754,
-43.8134841918945,
57.1721954345703,
50.7887153625488,
6.19629478454590,
6.08303356170654,
25.9634456634522,
45.0133514404297,
29.2601585388184,
-19.8450698852539,
73.6147003173828,
-2.51275634765625,
2.57146167755127,
94.8821640014648,
-28.4954700469971,
51.1105461120606,
8.00879287719727,
-15.1914339065552,
10.1953783035278,
-5.21877479553223,
32.5284919738770,
-47.2885398864746,
39.7344818115234,
-17.9973831176758,
-16.7618370056152,
40.5150451660156,
0.949840545654297,
65.5769729614258,
-12.7674160003662,
-9.29890251159668,
-26.9290390014648,
16.4521694183350,
-0.0969991683959961,
-41.8676261901856,
50.1077919006348,
-18.1735324859619,
37.6299667358398,
11.0139636993408,
-6.18987131118774,
14.3836498260498,
-7.42069149017334,
46.0654067993164,
9.51627635955811,
30.1627941131592,
-20.0043430328369,
36.2612304687500,
49.6376380920410,
-49.2603530883789,
-11.4941539764404,
-8.81587696075440,
14.8641519546509,
20.5003280639648,
41.0060348510742,
16.2688388824463,
-19.7299480438232,
21.9624748229980,
18.7735328674316,
-17.6125469207764,
23.1829185485840,
27.8135032653809,
-51.1465034484863,
50.4001693725586,
19.3208370208740,
-37.6103515625000,
61.6657791137695,
18.2166576385498,
33.2781829833984,
36.1902122497559,
31.8087120056152,
49.7525939941406,
-0.0649156570434570,
21.9712409973145,
46.0112533569336,
2.74699211120605,
12.8734273910522,
18.7438220977783,
-23.2525138854980,
20.6954689025879,
2.82586860656738,
-43.2385368347168,
-39.2253341674805,
29.0824851989746,
46.0597610473633,
-31.3892002105713,
-5.78099441528320,
-2.07354378700256,
15.3325862884521,
10.5270528793335,
-30.4815139770508,
-20.7514553070068,
-13.2488851547241,
-4.33557415008545,
-22.9301490783691,
14.7492389678955,
30.7424240112305,
-31.3683643341064,
-21.7635765075684,
33.4871940612793,
-16.0007743835449,
-47.3084335327148,
31.8528919219971,
39.9531593322754,
14.2223358154297,
10.7048940658569,
0.972815036773682,
-34.8108482360840,
8.65187263488770,
40.6982192993164,
-24.9871692657471,
14.8808488845825,
18.6847572326660,
15.3794202804565,
-3.53443336486816,
14.5204257965088,
82.6591491699219,
-11.2786388397217,
-16.6015281677246,
-15.3256959915161,
-24.2335987091064,
-6.23132276535034,
-11.2854185104370,
-9.25022411346436,
-33.5762100219727,
11.5539503097534,
6.74048328399658,
7.39416265487671,
-15.8025341033936,
49.0111122131348,
7.33247184753418,
-39.0175819396973,
46.8202209472656,
-21.6246128082275,
14.6093120574951,
5.47735309600830,
38.6343002319336,
20.2422122955322,
21.4142551422119,
17.6650772094727,
-10.3279018402100,
40.2393989562988,
-48.4296226501465,
-33.6907691955566,
3.65317344665527,
44.4610404968262,
-40.0283088684082,
2.64518642425537,
84.0111694335938,
-2.62505817413330,
-31.9049148559570,
25.5814952850342,
70.9737777709961,
28.5190048217773,
49.4521713256836,
-18.2030849456787,
-14.4596643447876,
-5.76837921142578,
-38.0228042602539,
-20.4422779083252,
-12.6950435638428,
-49.7964668273926,
-14.6629734039307,
32.5104064941406,
10.5012292861938,
53.7052192687988,
2.39960861206055,
-38.1593322753906,
-27.2342090606689,
39.6995086669922,
26.6750221252441,
-4.96085357666016,
-13.8962144851685,
-37.8244895935059,
-26.5281276702881,
-11.0944242477417,
21.5932044982910,
-30.1154270172119,
24.5546817779541,
37.2070503234863,
13.3466348648071,
1.89496326446533,
3.31762123107910,
18.7589988708496,
-41.7224578857422,
25.6116504669189,
27.5804862976074,
23.1723613739014,
-13.1317501068115,
-37.9549560546875,
-9.51313304901123,
-58.8601913452148,
47.7688331604004,
6.94078302383423,
-9.93437194824219,
67.5303039550781,
23.9789390563965,
26.2282161712647,
-10.7947711944580,
3.16568994522095,
-21.2706184387207,
-8.22236156463623,
-16.3113479614258,
-31.4498748779297,
36.4097671508789,
-27.3909988403320,
-22.4665393829346,
-5.29740238189697,
22.9254188537598,
43.3288803100586,
-53.6546134948731,
11.9021654129028,
59.3627662658691,
-43.3112754821777,
28.0585765838623,
69.1345214843750,
-21.6984138488770,
-13.9144582748413,
-17.0104770660400,
19.7654762268066,
20.6706962585449,
-44.9124565124512,
-12.4955816268921,
-23.0905342102051,
-48.2718467712402,
-33.6587066650391,
-6.39070463180542,
8.30290508270264,
-33.6156959533691,
-50.2597007751465,
11.0473423004150,
10.8143768310547,
-53.8154487609863,
0.828751206398010,
41.2326660156250,
-3.84484577178955,
-19.7886123657227,
-6.73123168945313,
-14.8996725082397,
23.5628356933594,
39.9406852722168,
2.04561066627502,
18.8279113769531,
-7.13355016708374,
-17.0353527069092,
36.8139953613281,
67.7057418823242,
-25.3781280517578,
-9.78456497192383,
44.1107864379883,
-57.7908172607422,
9.06251716613770,
40.1576576232910,
10.5520076751709,
42.5144386291504,
-17.0115833282471,
38.2235755920410,
39.3868408203125,
-44.4515457153320,
34.7320938110352,
9.34212493896484,
-36.2440528869629,
42.0021095275879,
47.0739364624023,
12.2765102386475,
57.2522468566895,
60.1583595275879,
-31.9082679748535,
26.3360691070557,
40.9379272460938,
-6.16408061981201,
11.5147638320923,
7.93341302871704,
-4.94315528869629,
-37.0716629028320,
40.9023666381836,
-3.58478450775147,
-56.5567092895508,
56.6301994323731,
20.3252582550049,
-12.1646938323975,
42.6181221008301,
-13.3002815246582,
-4.31057357788086,
48.5265274047852,
-27.8139266967773,
21.7584304809570,
60.2448501586914,
27.4539031982422,
46.0574798583984,
-19.7437438964844,
37.9971389770508,
36.2307281494141,
-7.29389715194702,
36.8204612731934,
-44.4070281982422,
-2.78779029846191,
40.1235008239746,
29.7420234680176,
45.5859985351563,
3.63214755058289,
35.8181571960449,
48.8099784851074,
24.0700626373291,
10.1208171844482,
23.4257335662842,
61.8413696289063,
-34.8693237304688,
-16.3605480194092,
79.6540451049805,
-1.93491363525391,
-9.06051349639893,
33.8748626708984,
9.49768161773682,
-35.9521408081055,
16.8924732208252,
19.5617218017578,
-22.8164520263672,
2.37054562568665,
-31.2436466217041,
43.0630645751953,
-1.45133495330811,
-30.4372520446777,
55.4290313720703,
-39.4507560729981,
32.9339256286621,
26.4449920654297,
-49.6935577392578,
53.0568428039551,
30.7122917175293,
-0.722547054290772,
34.6059570312500,
53.6859436035156,
12.8336362838745,
-15.8508567810059,
-27.5851173400879,
28.1134719848633,
64.6286315917969,
-37.9559936523438,
-20.8134956359863,
42.0081481933594,
13.0925531387329,
-49.7384185791016,
0.592236518859863,
71.0671997070313,
-28.2458934783936,
-13.2448835372925,
21.5241889953613,
-31.5271377563477,
14.6307201385498,
0.0787469148635864,
15.7828989028931,
16.7352313995361,
-41.3768424987793,
-5.21040058135986,
36.6728553771973,
55.4012565612793,
-7.52489423751831,
4.95865249633789,
51.1641159057617,
34.0315856933594,
13.8034238815308,
18.1419792175293,
64.5881729125977,
0.862535476684570,
-41.5555953979492,
-17.9717235565186,
1.50344729423523,
2.18736863136292,
-10.6135311126709,
-39.8392562866211,
-8.27308845520020,
72.1236038208008,
21.2435264587402,
14.7519683837891,
14.9411964416504,
29.9905548095703,
30.7177944183350,
-13.8377017974854,
41.4652938842773,
9.16294765472412,
28.7770576477051,
38.6470260620117,
-24.3636817932129,
-0.856274127960205,
-28.0779037475586,
7.48615550994873,
-22.2110939025879,
-48.4974937438965,
10.6830406188965,
-14.3413572311401,
45.5469703674316,
8.22393035888672,
-14.5890235900879,
8.15916633605957,
-5.40555381774902,
28.4987373352051,
29.1551399230957,
62.8358840942383,
-22.1392421722412,
-29.1140918731689,
1.43242728710175,
15.9607906341553,
45.5370254516602,
-40.1163940429688,
11.7512111663818,
-18.1668224334717,
-33.8954086303711,
51.0241317749023,
-37.0499076843262,
-48.0056648254395,
6.70803833007813,
15.3155155181885,
-12.8682012557983,
-22.1693229675293,
51.2356872558594,
1.18197441101074,
-5.68165111541748,
17.9665813446045,
15.8258705139160,
54.7279777526856,
-17.8318214416504,
-23.9709644317627,
2.99144363403320,
32.5005035400391,
13.8260402679443,
25.5953330993652,
42.4144401550293,
-32.6591644287109,
38.6947097778320,
37.3240623474121,
5.86909723281860,
-18.5106525421143,
-27.3812713623047,
49.0708198547363,
-14.8921184539795,
-52.0914878845215,
22.5822048187256,
3.13776969909668,
-45.4964294433594,
29.0085029602051,
20.0632934570313,
0.327191829681397,
-2.56660890579224,
-6.40806388854981,
74.4889984130859,
-16.5135898590088,
-0.571554183959961,
11.9628543853760,
-14.5341281890869,
64.1897125244141,
-21.2392559051514,
-34.9193725585938,
-6.51141262054443,
-20.4903316497803,
-30.8280696868897,
21.1778507232666,
-3.38932418823242,
-69.0297698974609,
6.13657569885254,
27.9006710052490,
-11.8734111785889,
-35.3937683105469,
-1.10658931732178,
-5.54900693893433,
34.1070022583008,
30.6563816070557,
-23.2973098754883,
11.0393819808960,
21.8527984619141,
46.8262939453125,
23.3658275604248,
1.55902385711670,
-11.1599760055542,
-15.3648910522461,
3.88727259635925,
-6.86826419830322,
-18.2039794921875,
-22.3238029479980,
23.9639797210693,
-12.2193765640259,
2.49053573608398,
69.1488037109375,
22.2388229370117,
46.8114700317383,
17.9350223541260,
6.55266046524048,
21.7683620452881,
-5.57957601547241,
40.4451980590820,
-7.27605438232422,
-27.7208557128906,
15.6252470016480,
19.7035102844238,
17.0151557922363,
-3.72815132141113,
-22.1791706085205,
-1.27913522720337,
54.2506256103516,
-4.90791034698486,
-42.0169181823731,
39.1728057861328,
28.0893440246582,
-16.8088283538818,
20.5177879333496,
59.1916046142578,
19.2058410644531,
10.3768062591553,
-23.2191925048828,
-32.1590042114258,
51.2851066589356,
-12.6037359237671,
-45.7060356140137,
-26.0818462371826,
6.29955863952637,
33.1760292053223,
4.48768424987793,
35.4290962219238,
-22.6313056945801,
11.4559173583984,
41.5883216857910,
-27.1093788146973,
9.54780769348145,
-3.69010138511658,
8.51460266113281,
22.1941204071045,
9.57376956939697,
0.934843957424164,
7.99510955810547,
39.2904968261719,
33.8699645996094,
40.4073028564453,
6.80523490905762,
18.3935718536377,
12.4237079620361,
-19.7812919616699,
-10.1601390838623,
-11.7862472534180,
-32.1190109252930,
-41.7138824462891,
-4.51780414581299,
-25.3185958862305,
-21.0805435180664,
-7.31149482727051,
-0.480260848999023,
14.0277652740479,
35.7799568176270,
-10.9890918731689,
-30.1716156005859,
44.8495178222656,
-53.4184532165527,
-22.9966220855713,
57.0568199157715,
23.6736335754395,
43.5040054321289,
16.3654098510742,
52.6240081787109,
30.0042304992676,
13.9198169708252,
31.9077777862549,
21.9342117309570,
38.8546791076660,
26.9407482147217,
51.9253196716309,
25.7657737731934,
51.5491943359375,
24.8779602050781,
-21.4007606506348,
15.1505470275879,
41.2051086425781,
12.8719100952148,
-48.1365966796875,
-3.02943515777588,
4.24140501022339,
38.1484680175781,
50.4330482482910,
21.1125488281250,
29.1232910156250,
22.2172756195068,
30.7085609436035,
31.1614303588867,
15.9505176544189,
18.3754673004150,
9.13725566864014,
-6.26403236389160,
38.2880020141602,
6.54563713073731,
29.5667667388916,
61.6442756652832,
-36.1942291259766,
10.9167461395264,
59.1608924865723,
1.20231246948242,
-32.3386688232422,
45.2198486328125,
54.4841270446777,
-5.97797107696533,
29.7276191711426,
-14.6141138076782,
30.5984687805176,
33.6716575622559,
16.7182102203369,
38.1662406921387,
-5.19602489471436,
52.3816184997559,
59.1836547851563,
45.1736450195313,
41.7755012512207,
-1.84827041625977,
-17.3452167510986,
45.5868339538574,
12.7900800704956,
-31.1978054046631,
72.0931320190430,
11.4390754699707,
-45.6099014282227,
8.24260997772217,
-8.20462799072266,
13.3159961700439,
7.31838417053223,
13.6658763885498,
25.6642017364502,
-10.7280998229980,
31.2254352569580,
48.9686203002930,
23.1863002777100,
56.1964492797852,
58.9720230102539,
24.4166393280029,
19.0545635223389,
69.6971359252930,
43.9400291442871,
-29.7731246948242,
7.34640884399414,
-14.7728223800659,
21.3844261169434,
2.52505302429199,
-10.2783784866333,
56.1749114990234,
-42.5701675415039,
8.10345554351807,
31.8154964447022,
-43.6394386291504,
10.9912681579590,
30.4884262084961,
-21.6157283782959,
1.94122886657715,
16.5865154266357,
7.29614019393921,
29.5573654174805,
-43.6608848571777,
-29.7594184875488,
-17.0047626495361,
4.02199077606201,
51.7551078796387,
0.844780862331390,
29.2682971954346,
19.1852302551270,
-2.86462402343750,
-9.37039852142334,
41.5496292114258,
53.9161376953125,
-14.8740653991699,
7.18344640731812,
22.9865207672119,
68.3278961181641,
4.24263572692871,
20.7909927368164,
64.2964324951172,
-4.88857269287109,
6.80981731414795,
-14.0024232864380,
32.9671821594238,
-33.2476196289063,
-56.4513244628906,
8.44196605682373,
-33.5458183288574,
9.49459171295166,
-4.55922508239746,
17.0929508209229,
20.2334613800049,
-54.4085235595703,
-20.2724208831787,
45.9269714355469,
50.4345550537109,
7.96858406066895,
-0.981654524803162,
-15.2014656066895,
-24.9345531463623,
-26.0641784667969,
48.9428863525391,
30.1825599670410,
-61.5030670166016,
17.1525974273682,
27.7254924774170,
-21.9223899841309,
38.2810401916504,
55.5816650390625,
-41.9814414978027,
2.81908798217773,
53.4546546936035,
45.4483108520508,
4.26594352722168,
-16.4965324401855,
73.3382492065430,
-13.6527194976807,
-9.74408817291260,
57.9159355163574,
26.1038589477539,
-26.4660301208496,
-16.0686817169189,
51.9710502624512,
-17.0820941925049,
38.7822036743164,
25.8176212310791,
-25.3316955566406,
38.0419883728027,
-40.6530075073242,
-28.2768993377686,
7.72751379013062,
7.85278463363648,
44.3105545043945,
13.4844303131104,
16.9826164245605,
5.25738334655762,
-24.7969474792480,
24.1827678680420,
56.8665122985840,
-22.1108379364014,
-35.3398742675781,
-6.18181610107422,
-11.5663852691650,
13.9272327423096,
-27.4033966064453,
34.4198532104492,
3.07509231567383,
-42.3397064208984,
23.7345123291016,
-35.4254951477051,
28.7086639404297,
56.5897636413574,
-14.9230670928955,
-24.5120468139648,
13.5296792984009,
-17.0861034393311,
-43.2025985717773,
-10.4477863311768,
0.331210136413574,
13.0826454162598,
-46.9742050170898,
-35.2533836364746,
7.13265180587769,
39.9499359130859,
-1.54238128662109,
-41.4959144592285,
-8.99327468872070,
6.39560794830322,
6.06289100646973,
-30.8041095733643,
-25.8742027282715,
-33.3943939208984,
1.76291966438293,
-24.2360725402832,
-47.7620010375977,
-19.6608695983887,
-5.94807434082031,
35.3467636108398,
-44.6812362670898,
-31.3503036499023,
59.1341857910156,
18.6135330200195,
2.29477953910828,
58.0818977355957,
11.0657529830933,
-53.6064720153809,
46.1295127868652,
17.2113285064697,
4.99671745300293,
65.1665039062500,
-10.7353630065918,
10.1019735336304,
1.47765779495239,
31.5999908447266,
11.7953548431396,
-51.8739814758301,
60.5787277221680,
5.55742549896240,
15.7939090728760,
20.4994354248047,
-17.0600051879883,
73.3148880004883,
22.6636505126953,
40.6288032531738,
-8.78744316101074,
-18.9544925689697,
37.9813880920410,
-29.9338912963867,
41.8118553161621,
6.80202198028564,
5.96698379516602,
41.3994941711426,
-27.4938964843750,
36.2896080017090,
-5.35425949096680,
-42.9612731933594,
33.9152069091797,
29.0506649017334,
-17.4399604797363,
-26.5972232818604,
30.5698966979980,
34.5448570251465,
-61.5045928955078,
-0.108009338378906,
47.7063522338867,
-15.2400188446045,
53.0295410156250,
48.1842994689941,
44.4790573120117,
-12.0448341369629,
-52.8622627258301,
7.01900053024292,
-12.6770439147949,
28.6561279296875,
-44.5211486816406,
-8.89335823059082,
38.9451293945313,
-29.4184474945068,
54.5064468383789,
-15.4010219573975,
17.0762252807617,
15.0873069763184,
-47.6397552490234,
89.7644729614258,
4.75665855407715,
-22.9369087219238,
48.6848907470703,
9.55476570129395,
13.9714603424072,
13.0775403976440,
21.2261047363281,
42.5461997985840,
-17.9772605895996,
7.62342643737793,
85.3603515625000,
-15.2652492523193,
12.4545001983643,
66.0465850830078,
-18.2823886871338,
-5.26905059814453,
43.7967872619629,
53.4904899597168,
-19.4300880432129,
0.182807922363281,
59.4629211425781,
22.9770946502686,
20.5474033355713,
-6.95803546905518,
40.4504241943359,
23.7597026824951,
-21.1991996765137,
30.5577430725098,
18.0134983062744,
8.85300827026367,
-8.64997577667236,
47.7760734558106,
20.0663146972656,
-43.5962791442871,
-9.57552528381348,
-11.8273458480835,
-15.3644361495972,
-40.2027435302734,
55.9900817871094,
48.7732734680176,
-55.2142295837402,
42.2536621093750,
30.1394481658936,
-3.51513671875000,
58.5623664855957,
30.8045673370361,
19.0036087036133,
50.4640998840332,
62.2327613830566,
18.1969795227051,
-39.0417823791504,
45.6545104980469,
62.7385292053223,
-23.7240085601807,
61.9628181457520,
31.7793121337891,
-62.5092163085938,
-12.2177352905273,
38.4525604248047,
42.1707382202148,
-22.9124145507813,
8.42746067047119,
31.6039104461670,
-22.0946197509766,
26.8109626770020,
46.9804534912109,
-12.7524547576904,
25.4002876281738,
27.9096717834473,
-26.8833332061768,
3.54973983764648,
-2.88611912727356,
-10.9125041961670,
3.01057744026184,
-11.1792802810669,
-39.4174499511719,
-13.7657537460327,
12.4819021224976,
8.43483924865723,
14.8136959075928,
55.1918258666992,
40.8564910888672,
-45.7197532653809,
58.5710449218750,
66.1783370971680,
-54.7633666992188,
16.9620704650879,
34.0170059204102,
-78.3001708984375,
10.8518199920654,
36.2892761230469,
-20.1792259216309,
30.1777839660645,
-16.3816661834717,
35.0141029357910,
-16.1490802764893,
-8.53889942169190,
67.7136840820313,
10.0296764373779,
7.54119253158569,
9.59908485412598,
14.8800277709961,
21.0900325775147,
58.9821701049805,
25.2112159729004,
11.4535093307495,
0.703738570213318,
27.8603725433350,
42.0829353332520,
7.09297084808350,
0.488538742065430,
-41.3932952880859,
3.01266670227051,
8.32756614685059,
-2.80050945281982,
43.6520423889160,
-4.61621379852295,
-55.2281265258789,
37.1916885375977,
16.7505149841309,
-11.5099639892578,
78.3819122314453,
-15.1215667724609,
-29.3115158081055,
61.6439895629883,
42.0367279052734,
-27.7431297302246,
-41.3930015563965,
65.7091674804688,
-5.76788902282715,
-73.4889373779297,
51.9202499389648,
57.8724441528320,
6.08107662200928,
-14.1826038360596,
7.31831789016724,
5.38604974746704,
18.2877063751221,
35.2211418151856,
-35.2179298400879,
10.4716396331787,
68.5773162841797,
-1.63174057006836,
-56.0424194335938,
13.5738162994385,
-19.6100540161133,
-42.2235069274902,
-11.9201469421387,
-38.3475494384766,
52.7159957885742,
-7.76360702514648,
-10.4363031387329,
10.4765892028809,
-38.7827339172363,
-25.3673381805420,
-20.3054542541504,
52.1262893676758,
14.3314762115479,
-35.9456672668457,
-30.4816684722900,
0.979497313499451,
11.6134576797485,
12.3070831298828,
0.350970983505249,
2.93408846855164,
9.98533821105957,
-31.9187774658203,
-13.0755920410156,
21.1092529296875,
46.2167243957520,
-46.1795921325684,
-38.4247665405273,
39.1830368041992,
-20.1927471160889,
-49.5058822631836,
-12.0884418487549,
49.6756248474121,
33.3617935180664,
15.6758365631104,
-5.01810932159424,
-23.0268058776855,
31.7081794738770,
-21.4996929168701,
-42.1165084838867,
3.76549124717712,
-46.4230041503906,
-15.4815464019775,
13.4012670516968,
10.9031572341919,
-1.78951358795166,
9.45510864257813,
30.5081863403320,
17.9289646148682,
61.2307357788086,
12.1427021026611,
25.3210258483887,
-4.80126762390137,
-27.3556747436523,
33.2897148132324,
18.6526832580566,
18.3023681640625,
-43.6380081176758,
30.6056499481201,
59.1875152587891,
8.01007652282715,
48.7126083374023,
19.6675910949707,
9.63242912292481,
13.7900257110596,
-9.87167072296143,
-15.6506175994873,
30.5430889129639,
-18.6497306823730,
-37.9806060791016,
-16.3403797149658,
-21.0326271057129,
22.2545547485352,
-34.4693794250488,
24.8797225952148,
4.03220272064209,
-43.0695419311523,
47.9649887084961,
33.1089553833008,
27.9380950927734,
-22.8361587524414,
7.70532035827637,
-10.1445741653442,
13.8031787872314,
58.9396209716797,
-22.4513092041016,
31.2613677978516,
-6.81676340103149,
15.6284809112549,
22.4777069091797,
-8.43040084838867,
46.3468513488770,
-25.5355625152588,
0.667093038558960,
39.1316337585449,
29.0443840026855,
23.7513370513916,
-17.5204601287842,
16.7500743865967,
24.5393886566162,
13.1914463043213,
57.2267036437988,
40.3113670349121,
-12.8858318328857,
6.79195451736450,
-6.06453943252564,
-29.6059150695801,
13.8064994812012,
39.4204025268555,
19.5444107055664,
-16.4324512481689,
-22.0899353027344,
-15.1690063476563,
-5.52465534210205,
24.0494995117188,
17.8446521759033,
-27.7821674346924,
-12.1818408966064,
7.58147430419922,
31.5875720977783,
32.1406021118164,
35.7787322998047,
43.7649421691895,
-22.6905555725098,
30.3173141479492,
73.0273666381836,
-16.7231979370117,
-28.1764831542969,
3.79624319076538,
-12.6454257965088,
-16.9229412078857,
-45.6089401245117,
3.96176338195801,
-0.650495052337647,
-16.7686882019043,
45.7324790954590,
-19.5663433074951,
46.1095542907715,
16.4791831970215,
-22.5823841094971,
53.0878601074219,
-18.8989715576172,
-25.5487899780273,
-34.1921386718750,
1.93277740478516,
45.0136451721191,
25.7219944000244,
-14.8624916076660,
-20.6891880035400,
59.9229354858398,
-12.9186220169067,
-20.6659069061279,
50.8843803405762,
46.5957794189453,
24.7014598846436,
11.3670005798340,
22.4460239410400,
-25.6602039337158,
38.0839920043945,
36.2446632385254,
7.15591573715210,
6.40036296844482,
7.01644134521484,
83.7018051147461,
-46.2957687377930,
11.4069843292236,
55.8887290954590,
-37.0105667114258,
53.8594131469727,
-7.66095542907715,
38.5510864257813,
84.3635101318359,
-36.4595718383789,
-18.3610229492188,
9.45268630981445,
-14.0116386413574,
29.4297943115234,
-19.8885173797607,
-33.3405761718750,
52.2029228210449,
-35.9062652587891,
-31.6954860687256,
-6.33040618896484,
30.9230766296387,
25.5972290039063,
-13.1316251754761,
78.6556854248047,
1.76746559143066,
-29.0504493713379,
-7.57153511047363,
56.6755905151367,
20.3850326538086,
-60.4053192138672,
23.9794750213623,
-12.3485221862793,
40.6654052734375,
-19.3036308288574,
-10.3947162628174,
39.9467811584473,
-37.9805679321289,
58.4914779663086,
18.6572227478027,
-29.2435874938965,
-11.4520235061646,
36.0546531677246,
-8.20750808715820,
20.0023651123047,
34.8410758972168,
-12.0272560119629,
42.6696701049805,
-35.1044540405273,
64.4406738281250,
25.9495086669922,
-17.3100204467773,
29.0307521820068,
-2.22363805770874,
66.1115264892578,
-26.7454795837402,
12.8449983596802,
16.8705482482910,
-15.5558395385742,
55.9127120971680,
21.4095649719238,
-12.1377305984497,
-23.5291080474854,
-5.00334405899048,
-22.8123855590820,
50.9766464233398,
-2.67600631713867,
-9.53998756408691,
16.3076019287109,
-41.9888572692871,
25.5686035156250,
-25.0718936920166,
30.4145603179932,
47.2586517333984,
24.4259414672852,
-15.8678007125855,
-42.8532371520996,
13.5617389678955,
-30.1171302795410,
-0.0949401855468750,
14.3400859832764,
14.5203361511230,
52.8322181701660,
35.8040161132813,
-9.24380779266357,
21.5375232696533,
2.95759701728821,
1.50041770935059,
40.2098083496094,
31.5971012115479,
51.4152488708496,
-35.6415252685547,
-12.6688346862793,
42.3356971740723,
-2.57164621353149,
56.1391296386719,
-11.7110729217529,
-34.3425254821777,
43.6527214050293,
1.98082828521729,
-11.6689186096191,
-3.63314342498779,
41.8648147583008,
17.7628154754639,
-37.3921089172363,
30.6601715087891,
44.4870185852051,
-31.0441169738770,
-49.1562347412109,
29.2786903381348,
35.2734756469727,
-40.4009628295898,
34.3616790771484,
47.3481864929199,
-7.80751562118530,
25.0741806030273,
17.6849842071533,
53.0805282592773,
24.0543918609619,
22.2964859008789,
72.2829284667969,
25.3624458312988,
28.8034839630127,
22.1430778503418,
11.5839443206787,
30.5719146728516,
13.9508457183838,
7.48474311828613,
14.9577226638794,
39.5639801025391,
0.315278053283691,
-31.1980667114258,
55.3992462158203,
17.5432815551758,
-23.5113697052002,
25.6301593780518,
-35.6562881469727,
5.03618431091309,
19.9017696380615,
16.5953025817871,
51.3202056884766,
-31.6290359497070,
11.4241428375244,
-19.7506675720215,
6.03123664855957,
76.2747039794922,
4.51276779174805,
44.3501205444336,
62.0516853332520,
22.2685947418213,
-7.30582380294800,
8.47667694091797,
-20.1080493927002,
-8.97680187225342,
-10.1860466003418,
-33.4935150146484,
26.6016960144043,
-41.8753890991211,
-3.19132041931152,
56.0102462768555,
-23.7671279907227,
-5.94136142730713,
30.2247066497803,
25.2901229858398,
1.24192333221436,
24.5270042419434,
33.9056930541992,
30.0278186798096,
11.6495227813721,
-32.9525222778320,
65.1820831298828,
19.8448562622070,
-55.7873535156250,
-9.83528995513916,
-18.2635021209717,
59.4236145019531,
-19.2169494628906,
-2.20944404602051,
66.5398712158203,
-65.4273529052734,
-19.6077194213867,
-4.48384332656860,
-25.4968986511230,
17.1890010833740,
48.2724876403809,
51.9009628295898,
-8.20364952087402,
-34.5140075683594,
2.13577079772949,
32.4897384643555,
12.9511184692383,
17.3297672271729,
48.8714141845703,
39.5585136413574,
-40.5390815734863,
-2.91640257835388,
32.5145072937012,
-46.3070259094238,
-8.10695648193359,
3.65522646903992,
6.02210950851440,
11.7771444320679,
-10.5619029998779,
-37.9323654174805,
-16.2590293884277,
58.1228828430176,
-12.1871767044067,
-21.5551681518555,
-16.6602745056152,
-20.2067813873291,
21.4286499023438,
28.8425483703613,
17.0126914978027,
-45.3309745788574,
12.5650243759155,
55.6025238037109,
-12.2719020843506,
2.96038103103638,
66.4010772705078,
-26.4540157318115,
-33.4613952636719,
45.6531906127930,
-33.3741340637207,
-22.5768775939941,
20.7725257873535,
-2.45992755889893,
-8.75305843353272,
51.9929237365723,
7.99501800537109,
-48.3564949035645,
63.9885597229004,
14.5966434478760,
-11.4433345794678,
49.4478607177734,
15.1500558853149,
36.5691146850586,
17.0446414947510,
-19.5678863525391,
26.7814216613770,
54.2900466918945,
9.64300823211670,
-7.16867399215698,
-20.6619091033936,
18.3014526367188,
54.3237152099609,
-24.9230594635010,
41.3335800170898,
-8.59810733795166,
-38.1148757934570,
56.7470245361328,
-36.0111427307129,
20.5891551971436,
24.0098762512207,
-44.2292861938477,
44.6187248229981,
47.9751014709473,
-25.2545013427734,
-22.4869689941406,
-1.89902853965759,
10.4187946319580,
12.5064001083374,
-33.6931571960449,
45.2097816467285,
3.33386802673340,
-23.1271209716797,
42.9844093322754,
-33.2817077636719,
0.750371932983398,
-1.31514668464661,
21.0454635620117,
23.9502868652344,
-1.40753340721130,
10.8785820007324,
-36.1906738281250,
33.9226913452148,
52.4517211914063,
41.4887466430664,
22.5580368041992,
55.8133850097656,
35.1772766113281,
-29.9874916076660,
41.5172080993652,
16.6912841796875,
10.4484777450562,
-18.8729553222656,
22.1722316741943,
-0.550384521484375,
-34.6575508117676,
38.2850646972656,
-23.7828540802002,
-12.3278656005859,
-36.8504295349121,
-21.1310462951660,
43.5333480834961,
18.1777839660645,
-2.96533393859863,
-19.3655052185059,
0.374233245849609,
64.3721618652344,
-0.0606002807617188,
-5.46936035156250,
23.8419609069824,
-32.8359298706055,
50.2892379760742,
22.4591236114502,
19.8418712615967,
-5.51439857482910,
-61.4138717651367,
15.9840259552002,
-1.81886577606201,
-13.2241497039795,
38.1992950439453,
-12.7262535095215,
17.9970722198486,
42.0080413818359,
-26.8206920623779,
63.0871391296387,
0.992663860321045,
-6.89114522933960,
35.9086761474609,
10.6754121780396,
35.0752410888672,
21.5625305175781,
48.7091102600098,
55.6530189514160,
21.5382633209229,
2.50154876708984,
64.9480972290039,
0.644436836242676,
16.6075744628906,
48.5062179565430,
-36.0864410400391,
-13.9677877426147,
4.75631380081177,
17.6570396423340,
-23.6686859130859,
-22.3514118194580,
13.6539726257324,
26.4072895050049,
5.70113515853882,
-5.33356714248657,
50.0592231750488,
23.8596725463867,
-6.59862804412842,
20.5496635437012,
33.2125930786133,
1.53898084163666,
33.1687850952148,
21.6187229156494,
-16.6974697113037,
61.3512725830078,
10.4830827713013,
-32.6897964477539,
33.0992164611816,
52.2373962402344,
32.6808128356934,
-1.36523342132568,
28.1308727264404,
36.5622100830078,
-27.4860286712647,
-31.5559463500977,
6.13312244415283,
-16.5491313934326,
13.2934665679932,
5.08467960357666,
-35.7357559204102,
7.86369132995606,
-11.3207464218140,
0.803871154785156,
-9.59871482849121,
-27.7541618347168,
5.30563735961914,
-28.6139011383057,
-5.49802684783936,
-8.63078022003174,
-2.89985275268555,
84.9175262451172,
-2.16072082519531,
-37.5677528381348,
53.1084747314453,
5.66489219665527,
27.9437389373779,
16.3734550476074,
-37.0447120666504,
-19.0851955413818,
-41.1932525634766,
-7.34792423248291,
-33.0814170837402,
38.0569190979004,
16.1591930389404,
-32.4323577880859,
48.0631866455078,
-35.4111328125000,
47.3528709411621,
14.9853706359863,
-26.0932044982910,
76.4735488891602,
13.7709960937500,
26.9421424865723,
28.1601181030273,
36.4787445068359,
54.2112045288086,
16.0055484771729,
42.9003829956055,
43.1249008178711,
-2.23687076568604,
37.7195243835449,
54.7580261230469,
52.9971923828125,
11.7666664123535,
-21.0486469268799,
46.4143371582031,
30.6149864196777,
20.1524353027344,
7.01649951934814,
2.94306826591492,
46.6932640075684,
60.3487663269043,
7.54521369934082,
-33.9327354431152,
-19.3920421600342,
-3.44193840026855,
43.8590545654297,
43.8848381042481,
-3.83427286148071,
-22.9753913879395,
33.3722114562988,
5.91334819793701,
-32.0116767883301,
15.3345870971680,
2.20530557632446,
17.6598815917969,
10.6479816436768,
-11.6543598175049,
-11.7954196929932,
22.0396842956543,
42.9782447814941,
-31.9652519226074,
0.427701473236084,
38.9142112731934,
15.5075054168701,
-22.0569267272949,
-0.132557868957520,
26.7968597412109,
-40.3701362609863,
15.6125125885010,
67.1614074707031,
44.3468475341797,
-36.9003715515137,
-45.5619888305664,
14.2901697158813,
15.7222108840942,
66.9792404174805,
23.8404731750488,
-18.7769145965576,
-16.1929550170898,
11.5605678558350,
9.71964836120606,
-36.5362777709961,
39.9413642883301,
-22.7546920776367,
-46.0942039489746,
27.1485195159912,
-43.3051567077637,
-8.85359096527100,
6.15334892272949,
-57.4469795227051,
-20.7463111877441,
-18.9176864624023,
-30.1383533477783,
18.1248970031738,
-1.63933908939362,
-16.3519077301025,
22.6344909667969,
15.1604804992676,
-19.7221679687500,
-13.3276882171631,
12.2182464599609,
19.5345191955566,
39.5607719421387,
4.52664947509766,
-22.6121139526367,
38.2463836669922,
8.24575424194336,
-40.6765785217285,
-5.47738933563232,
-8.03812599182129,
62.5459365844727,
18.4611301422119,
-41.4220199584961,
73.2268295288086,
34.1453781127930,
32.2788276672363,
26.4616069793701,
-20.8654365539551,
13.2462463378906,
0.869947433471680,
-22.6899032592773,
-8.12642955780029,
-5.55626153945923,
-47.5742111206055,
-36.8806686401367,
23.6318550109863,
39.0489730834961,
-11.6818876266480,
-7.10817527770996,
38.0371627807617,
66.9502792358398,
10.9368801116943,
9.73084926605225,
43.0862197875977,
-31.0623340606689,
38.2909240722656,
51.4125556945801,
18.4314212799072,
-14.2126760482788,
3.65031623840332,
99.1259460449219,
-21.1065883636475,
-5.14787244796753,
10.6410961151123,
-42.8918266296387,
20.7835044860840,
13.1891117095947,
21.9709339141846,
-8.14703845977783,
-4.35244417190552,
-0.0881843566894531,
-22.5758533477783,
-17.1168956756592,
-4.11221122741699,
11.4328289031982,
8.04073143005371,
58.3274116516113,
24.5858345031738,
-39.1403732299805,
1.98210763931274,
35.1835823059082,
27.1508560180664,
60.2481765747070,
18.9730777740479,
-21.0894317626953,
-35.1616668701172,
1.46266174316406,
62.7299880981445,
17.6299133300781,
39.9066543579102,
-26.8642559051514,
-45.2391586303711,
-6.44915819168091,
10.8834009170532,
7.35559320449829,
-46.2594261169434,
17.6976165771484,
54.0058593750000,
39.1770095825195,
25.6817684173584,
54.7091979980469,
-0.671254634857178,
-21.7188529968262,
28.5877838134766,
-14.8591499328613,
-23.4266510009766,
-2.32798457145691,
-3.40315723419189,
-60.9776458740234,
-31.4649543762207,
7.57855892181397,
-7.66076612472534,
-15.3965425491333,
-2.98878860473633,
27.7057838439941,
-35.0746231079102,
17.1698799133301,
17.3488121032715,
-6.55108308792114,
-4.93531799316406,
-33.5807723999023,
55.6004257202148,
34.5711975097656,
27.6630668640137,
43.7934494018555,
60.1016044616699,
-10.4327239990234,
15.2959232330322,
42.8491630554199,
-29.6253738403320,
6.90779781341553,
-19.2664813995361,
42.4785270690918,
-24.8554992675781,
-20.1433105468750,
55.7588348388672,
-10.1967353820801,
-36.5230407714844,
-14.9830255508423,
17.6325492858887,
-26.7671966552734,
7.43287420272827,
-6.53819799423218,
-17.5861396789551,
-31.3943538665772,
-25.4679756164551,
49.7207450866699,
4.23790025711060,
7.42348718643189,
4.51271724700928,
12.2315711975098,
38.0471229553223,
-0.287051200866699,
25.2315864562988,
4.85562849044800,
-20.1809520721436,
14.4259567260742,
10.2519674301147,
-8.48547744750977,
32.1806678771973,
17.3295974731445,
-38.7840347290039,
28.3066463470459,
-8.29131221771240,
-22.4356842041016,
44.2576942443848,
-47.9568099975586,
22.9040336608887,
36.7746810913086,
-69.6593399047852,
35.7901840209961,
27.4806118011475,
18.4456977844238,
-29.0059051513672,
22.5495853424072,
48.5310287475586,
-48.9009819030762,
52.1075057983398,
-19.8701457977295,
17.6440086364746,
14.5466022491455,
-34.4048652648926,
-22.0155105590820,
-12.8960189819336,
34.4508590698242,
-14.2089939117432,
-8.38347244262695,
-33.1308059692383,
39.1167488098145,
-24.9246425628662,
13.4467811584473,
15.9286117553711,
-54.0501556396484,
86.7507247924805,
5.77596569061279,
43.5784568786621,
31.4316921234131,
-25.2577362060547,
25.6316871643066,
10.5294675827026,
24.4954013824463,
-17.1913948059082,
28.4270591735840,
33.0554351806641,
22.7907066345215,
34.5744705200195,
8.39726829528809,
45.8068466186523,
6.59843444824219,
-26.6974277496338,
17.2931385040283,
52.8140449523926,
27.4542922973633,
-7.63315773010254,
-3.79469680786133,
41.6549682617188,
29.7177314758301,
2.43452620506287,
34.6165275573731,
-28.4390563964844,
-21.4473304748535,
63.3871917724609,
45.4579811096191,
-4.68706226348877,
-21.9181461334229,
19.7720565795898,
52.4844512939453,
-24.6507415771484,
9.51382541656494,
61.5388488769531,
-44.2968444824219,
18.7021713256836,
12.0618162155151,
-11.0831661224365,
17.6216735839844,
-60.6199760437012,
35.4575691223145,
2.83522796630859,
-26.1209430694580,
11.1887559890747,
-0.429985046386719,
52.4082908630371,
-32.6162605285645,
38.7130241394043,
71.1366653442383,
-5.85675573348999,
10.9017696380615,
-22.3493881225586,
43.8248939514160,
25.5794258117676,
32.0130920410156,
12.2473773956299,
-33.4201660156250,
55.9116668701172,
36.0595512390137,
-8.63056278228760,
13.2225923538208,
14.5387325286865,
-72.7163162231445,
40.4699211120606,
7.01304054260254,
-2.71441268920898,
35.8734359741211,
-49.6143379211426,
36.7241249084473,
-34.5608139038086,
44.1837234497070,
-6.55388927459717,
-26.5840892791748,
25.1120777130127,
-4.91767120361328,
72.2216720581055,
12.3831110000610,
-5.07466506958008,
7.09819507598877,
57.3631706237793,
2.56679940223694,
12.6512203216553,
33.2410430908203,
42.3587570190430,
21.9629898071289,
-21.1985607147217,
18.7624778747559,
-12.2239274978638,
47.2738494873047,
-16.8118667602539,
4.50478792190552,
31.7222118377686,
-55.0546646118164,
23.3786296844482,
52.2097129821777,
28.8966751098633,
-11.3575906753540,
2.79763936996460,
-1.88057136535645,
-15.2996969223022,
28.6159553527832,
-9.39226055145264,
-0.0157973468303680,
-30.7440681457520,
-10.0309019088745,
75.1652908325195,
17.7259559631348,
27.2733001708984,
-4.18418502807617,
5.10827827453613,
53.0383033752441,
-5.71471357345581,
-12.5761890411377,
13.6367454528809,
8.31330490112305,
-52.6184158325195,
19.5872268676758,
6.55011558532715,
-38.7786521911621,
74.1821746826172,
4.69456481933594,
-31.6935653686523,
12.8513774871826,
6.75061845779419,
-19.0846042633057,
-10.3612155914307,
63.9132041931152,
9.57910442352295,
-33.0803413391113,
-21.1502304077148,
38.7981948852539,
23.0461273193359,
-40.9742469787598,
35.5728874206543,
3.45276689529419,
-34.2812156677246,
34.5863876342773,
11.4204654693604,
-41.2094116210938,
42.8580055236816,
-2.66937065124512,
-0.00417900085449219,
35.8949317932129,
-44.2989578247070,
77.4172363281250,
44.7438850402832,
-39.4322891235352,
11.6205253601074,
31.8966331481934,
27.0114669799805,
30.7846031188965,
-7.51689147949219,
-29.2972698211670,
-4.10405063629150,
-50.4760284423828,
5.25603294372559,
48.7162895202637,
31.9604759216309,
15.6327857971191,
5.51057243347168,
12.8426570892334,
18.1847667694092,
46.7113571166992,
-3.99744319915772,
3.70127964019775,
21.8112812042236,
-28.2879905700684,
51.4853820800781,
55.1948471069336,
21.6762485504150,
21.0988121032715,
11.3437690734863,
45.2660751342773,
-46.1891555786133,
14.3393545150757,
27.1436843872070,
-33.3991279602051,
6.95340442657471,
-35.6395988464356,
15.3501586914063,
2.39472508430481,
33.6586990356445,
8.39846897125244,
-25.3149013519287,
21.3300323486328,
-17.4138011932373,
60.3884162902832,
46.4438362121582,
21.3510322570801,
-3.18190002441406,
-35.8198928833008,
21.4394245147705,
54.7224769592285,
17.9385719299316,
-15.6269054412842,
61.4009552001953,
-3.59214019775391,
-17.1835670471191,
72.8125915527344,
43.0580177307129,
-45.6321678161621,
-28.1207790374756,
56.7233390808106,
-36.1413269042969,
10.7843170166016,
59.2008857727051,
-6.99437427520752,
-32.5784378051758,
2.28882598876953,
70.9466400146484,
42.4279251098633,
40.6808357238770,
18.8750534057617,
47.3283348083496,
56.2482566833496,
54.7703628540039,
-3.75041580200195,
-5.23051071166992,
10.6520566940308,
-16.5539512634277,
43.9661750793457,
16.7000141143799,
53.1851158142090,
11.2392091751099,
39.8539962768555,
30.8283004760742,
-27.5280666351318,
-0.0245256423950195,
-43.7049331665039,
-12.7651052474976,
-25.8894462585449,
82.5075759887695,
10.0074100494385,
-41.1486930847168,
77.3958053588867,
-19.2043323516846,
42.9920730590820,
-7.98612880706787,
7.42513275146484,
55.9486770629883,
7.40340948104858,
61.1814804077148,
-22.4750366210938,
29.5016746520996,
-10.3187789916992,
-44.8147468566895,
52.8656654357910,
32.3055877685547,
-13.7024888992310,
-18.4161396026611,
49.2616882324219,
59.8056793212891,
11.0337209701538,
27.0852890014648,
52.9574661254883,
-28.1533088684082,
-35.7360496520996,
12.4072036743164,
5.66245651245117,
-13.7329568862915,
-0.797314167022705,
7.06495237350464,
12.5838756561279,
-2.51922369003296,
-30.2478027343750,
-13.5703516006470,
-11.0924968719482,
31.6616115570068,
43.9569778442383,
38.7732696533203,
35.6313476562500,
45.6573791503906,
50.5391693115234,
3.15631294250488,
10.6311073303223,
45.1890296936035,
1.21829700469971,
9.47292709350586,
69.2674636840820,
26.8501720428467,
5.59191036224365,
27.0242462158203,
12.8822174072266,
-59.5642127990723,
18.0360107421875,
24.4347457885742,
-50.4586601257324,
47.7542114257813,
-31.5884857177734,
-27.9071846008301,
55.5930519104004,
19.7560462951660,
-2.19186973571777,
-35.0794372558594,
-21.6674270629883,
2.47430801391602,
46.5374412536621,
-28.2258071899414,
-18.8801860809326,
65.9510726928711,
23.8617877960205,
22.0835018157959,
-16.5961437225342,
14.7897768020630,
36.7617645263672,
16.2999191284180,
47.2225341796875,
8.27114105224609,
-26.1382942199707,
-32.9041633605957,
13.5436763763428,
-15.6243677139282,
-38.7341346740723,
44.9361495971680,
46.2557220458984,
19.6527252197266,
28.7070693969727,
39.5023612976074,
-14.2476902008057,
8.83574008941650,
19.3575000762939,
3.11763453483582,
49.7184753417969,
-13.2509193420410,
38.8570365905762,
37.2081985473633,
-26.0645408630371,
56.3165740966797,
15.2909898757935,
8.10293865203857,
10.7764034271240,
-37.9796524047852,
-12.5249013900757,
15.4826021194458,
36.4883460998535,
7.81368017196655,
-36.4020652770996,
-0.534532546997070,
47.1989402770996,
-29.6223106384277,
41.6004028320313,
22.5034122467041,
-36.4383163452148,
42.8891754150391,
-20.9711780548096,
52.0005950927734,
2.69573020935059,
0.187061309814453,
36.2476730346680,
-25.2919883728027,
-6.43366050720215,
3.15944576263428,
68.7787017822266,
-25.4369850158691,
-2.15654945373535,
70.0425186157227,
-15.7955341339111,
-13.9331493377686,
-12.4622325897217,
-39.4853134155273,
17.5793075561523,
10.8518171310425,
20.3153858184814,
47.1979789733887,
-38.5267105102539,
-17.7701244354248,
36.2743988037109,
43.3893127441406,
0.852092623710632,
28.7498092651367,
28.8475513458252,
-30.4930763244629,
36.3434791564941,
33.9074516296387,
5.03273868560791,
31.0414829254150,
-0.0778491497039795,
-20.2553863525391,
53.0375251770020,
65.6403350830078,
-24.2863807678223,
-39.4470825195313,
36.3632316589356,
21.2532672882080,
23.6106986999512,
56.3661956787109,
38.3279571533203,
48.9236450195313,
35.0140571594238,
27.4900207519531,
-4.50802803039551,
27.4918746948242,
-10.0069942474365,
-10.9396238327026,
87.4479827880859,
-11.4066429138184,
-45.2855987548828,
-19.6076145172119,
2.08344006538391,
24.1230278015137,
15.5330333709717,
-25.6207427978516,
-42.3953628540039,
3.17624855041504,
-52.9503097534180,
42.1565361022949,
21.7746753692627,
-37.6222381591797,
63.9243431091309,
-5.47830390930176,
53.6055793762207,
65.2004852294922,
-20.0356712341309,
-3.43672704696655,
37.6853790283203,
-19.3965663909912,
-10.9097366333008,
50.4740524291992,
-32.9485664367676,
2.98761940002441,
51.6421203613281,
19.9829788208008,
-5.39308929443359,
54.7391700744629,
21.2048320770264,
11.1920051574707,
23.8441734313965,
-59.3015480041504,
3.37220191955566,
37.6726455688477,
-8.67206382751465,
-33.0172271728516,
-27.7727413177490,
-34.5473365783691,
34.5929603576660,
-12.3054981231689,
-37.0931205749512,
72.4101104736328,
12.0088710784912,
23.0352001190186,
56.0658149719238,
45.8219871520996,
46.4198493957520,
-34.4161529541016,
-28.8052883148193,
48.7593078613281,
13.9401531219482,
0.973476409912109,
18.2246265411377,
-32.2839050292969,
-14.5634374618530,
-45.3479003906250,
0.802691459655762,
54.2313880920410,
-53.0981292724609,
23.1881942749023,
21.0963134765625,
1.46447086334229,
51.6310424804688,
-7.95106697082520,
7.82512187957764,
-37.1956291198731,
-16.2519226074219,
23.3727092742920,
1.05101740360260,
17.2915611267090,
-22.6489181518555,
26.8175239562988,
16.5607051849365,
-8.02772712707520,
52.2998504638672,
5.03875732421875,
32.1643943786621,
-6.11444997787476,
-3.61247348785400,
67.9643630981445,
6.16745805740356,
29.5203781127930,
3.74097299575806,
-15.7159051895142,
-26.7170448303223,
-15.9718933105469,
46.6589889526367,
38.2070312500000,
27.2283153533936,
39.9319381713867,
49.6523818969727,
36.9349403381348,
14.0632343292236,
-5.61486291885376,
65.2734985351563,
-5.41209411621094,
-14.1762647628784,
52.1428527832031,
12.4210395812988,
31.0953502655029,
13.4968070983887,
42.0402030944824,
-11.6687030792236,
39.4859580993652,
56.5528106689453,
3.97301435470581,
74.0119476318359,
-5.29617309570313,
2.00172424316406,
33.5798988342285,
54.3765640258789,
33.3776855468750,
20.8768711090088,
9.18632316589356,
-25.9472141265869,
68.3609008789063,
-2.19580459594727,
21.9570350646973,
29.6875000000000,
-16.8787498474121,
10.6618194580078,
-44.4618034362793,
24.4409580230713,
44.8491439819336,
12.4220256805420,
-0.562357604503632,
15.5537042617798,
7.36073112487793,
55.5461616516113,
1.71018600463867,
-19.4780521392822,
52.5082130432129,
-39.5884399414063,
62.9826049804688,
48.8187828063965,
-7.98062705993652,
-0.238776206970215,
-26.2842826843262,
27.3791790008545,
-20.1830081939697,
-31.2936019897461,
-0.570426464080811,
-19.9951877593994,
-51.5654373168945,
-20.6799697875977,
-29.6191577911377,
-12.8219070434570,
51.7230300903320,
-19.4512577056885,
7.23759078979492,
67.6808471679688,
-13.6178607940674,
-23.1141948699951,
35.5142936706543,
-14.8332366943359,
-31.5417251586914,
23.1861648559570,
-13.5206270217896,
45.1368484497070,
0.710266113281250,
-63.7628173828125,
39.4026641845703,
-32.4789619445801,
-29.8817825317383,
13.5313911437988,
10.2540016174316,
16.4701232910156,
7.91399765014648,
44.5368309020996,
-27.2485389709473,
-15.1250143051147,
8.70686244964600,
31.0001945495605,
36.1903800964356,
-32.7746047973633,
47.7774887084961,
35.0727958679199,
52.1614990234375,
53.9889831542969,
-3.13437557220459,
53.9756050109863,
12.0223999023438,
-10.6696853637695,
-6.34760379791260,
-20.4611911773682,
-30.9776496887207,
49.1069564819336,
10.0599174499512,
-44.7688140869141,
-6.94418478012085,
-25.1213283538818,
51.2915840148926,
-44.4779624938965,
27.7338428497314,
31.1496887207031,
-22.7343082427979,
61.9155883789063,
-59.4576187133789,
46.0848808288574,
13.0331544876099,
-51.8865051269531,
53.2298889160156,
17.3608703613281,
31.8012771606445,
44.2784347534180,
8.27722740173340,
4.53514051437378,
61.3886032104492,
30.5352840423584,
-43.7541351318359,
0.390757560729980,
37.5852279663086,
10.3111114501953,
-42.3599777221680,
-25.7192459106445,
39.4219741821289,
-20.5079784393311,
-19.6815376281738,
64.7061233520508,
-13.4145679473877,
-29.2053318023682,
57.7568359375000,
22.0525436401367,
32.4327049255371,
62.9734077453613,
37.7961349487305,
51.1947326660156,
28.4369544982910,
70.8124465942383,
9.36156082153320,
-19.1349678039551,
90.4926452636719,
43.2515182495117,
42.6649551391602,
-0.948599100112915,
-23.9913101196289,
18.3342323303223,
19.0576057434082,
62.7695503234863,
20.2839012145996,
35.1102790832520,
-18.7296657562256,
-9.61527252197266,
74.7066726684570,
-31.3439617156982,
33.9694213867188,
60.0140762329102,
-30.0810317993164,
-18.2972240447998,
-9.15104675292969,
-32.8763771057129,
-24.5907135009766,
-5.02876567840576,
47.6360092163086,
-6.84045934677124,
-46.1218261718750,
48.8110809326172,
-26.6746120452881,
2.99651575088501,
-14.7728977203369,
5.92126083374023,
41.0998420715332,
-13.6638832092285,
21.8102416992188,
-42.6357955932617,
2.52974033355713,
45.2191352844238,
28.8111019134522,
-4.63700723648071,
21.3593845367432,
61.3858032226563,
17.6863632202148,
-17.0319004058838,
35.8282318115234,
26.3212852478027,
-38.8131141662598,
58.7869377136231,
-15.4450778961182,
-34.7781524658203,
43.0761909484863,
-31.4570579528809,
-7.29603862762451,
5.45226573944092,
-32.9567871093750,
18.7608432769775,
-7.62386131286621,
-23.5545730590820,
33.9576225280762,
-29.0062274932861,
-31.9205474853516,
31.8778896331787,
41.1395339965820,
-17.5455169677734,
-56.5975952148438,
9.71665191650391,
39.8952255249023,
-2.31094169616699,
-44.4589614868164,
14.7616167068481,
-14.0059547424316,
-35.1409606933594,
51.8646125793457,
-13.7024087905884,
17.4918022155762,
12.6008014678955,
-20.6205101013184,
53.1775588989258,
26.6848716735840,
53.6681251525879,
-10.4619264602661,
-37.6311416625977,
-2.24955391883850,
11.9212265014648,
27.3305969238281,
-52.2235565185547,
23.0394744873047,
38.2337493896484,
38.5502281188965,
23.1530952453613,
-44.5863418579102,
9.90741729736328,
16.5399398803711,
33.3197669982910,
14.2803077697754,
21.9610099792480,
-23.3548049926758,
-0.371202468872070,
18.3593082427979,
-53.5899505615234,
3.49637603759766,
-30.3319339752197,
-0.643348693847656,
-2.90954136848450,
7.14117860794067,
66.6960906982422,
-41.2368850708008,
-51.1201248168945,
16.4703540802002,
50.0670089721680,
14.9352836608887,
48.2048339843750,
26.5479660034180,
-13.6798143386841,
58.1321945190430,
16.3120651245117,
28.6657180786133,
5.34193754196167,
-12.4932441711426,
32.8587989807129,
33.7530479431152,
-30.3071556091309,
-0.295465469360352,
56.8641700744629,
-49.8993797302246,
35.2523536682129,
52.1834907531738,
-27.3557415008545,
-22.1528205871582,
-16.5039520263672,
52.6583786010742,
48.7328033447266,
9.56237697601318,
3.35758495330811,
35.0399208068848,
53.3454437255859,
20.0824527740479,
-31.1705036163330,
-32.7822799682617,
38.0514411926270,
-6.93294525146484,
-38.0435791015625,
38.3615150451660,
-11.5836696624756,
-44.6180267333984,
-42.5004806518555,
-8.60659503936768,
38.2808456420898,
-41.9814071655273,
29.7386188507080,
74.3948287963867,
6.95183753967285,
27.1478900909424,
24.4494857788086,
60.6619262695313,
21.5290699005127,
42.6770362854004,
18.2918701171875,
-25.0364418029785,
66.8683929443359,
22.6081161499023,
48.4546127319336,
8.36963939666748,
15.6432971954346,
59.5092163085938,
-12.2695636749268,
12.3346509933472,
1.28368186950684,
-1.55151081085205,
-44.0106964111328,
5.68800354003906,
53.6947288513184,
2.41512966156006,
16.4547443389893,
-7.13803625106812,
-5.34280967712402,
-19.8239955902100,
19.6984405517578,
60.5359115600586,
-23.2953758239746,
-25.8414516448975,
38.5434722900391,
33.0559730529785,
-36.9537277221680,
-34.9853897094727,
60.6815605163574,
9.91533851623535,
-45.3505363464356,
43.4890213012695,
-0.362816810607910,
16.7481555938721,
48.4840736389160,
-18.9031543731689,
40.4408988952637,
34.9909629821777,
33.6529388427734,
4.54942989349365,
-0.634710311889648,
74.8273544311523,
-0.154485702514648,
49.7220611572266,
36.7912025451660,
-22.0899906158447,
54.3248596191406,
-30.0971527099609,
-46.0769958496094,
-16.2521972656250,
-30.1042327880859,
-32.2615394592285,
-34.1612663269043,
39.7989273071289,
22.6773376464844,
8.31641101837158,
12.9878149032593,
-21.7014522552490,
6.92462825775147,
13.8997116088867,
15.9903450012207,
-27.8312835693359,
-3.78975677490234,
76.2260589599609,
30.0265560150147,
29.1593818664551,
30.7433509826660,
-19.5385837554932,
27.0350589752197,
53.1807937622070,
-34.6899337768555,
-3.05463981628418,
66.0678405761719,
2.26490020751953,
-59.5872726440430,
6.26393318176270,
66.5684509277344,
-56.7903594970703,
-30.4548530578613,
40.1958160400391,
-46.5608444213867,
25.0265254974365,
76.7759704589844,
-13.4903392791748,
-37.2857589721680,
20.0785179138184,
56.3483085632324,
24.8947315216064,
43.5810699462891,
63.6199188232422,
11.0929021835327,
-10.7303705215454,
40.5959548950195,
54.5166816711426,
-12.0021581649780,
24.5798969268799,
59.1069831848145,
-27.6800632476807,
7.45683956146240,
-3.00845336914063,
-34.7015419006348,
37.3801116943359,
-34.1037712097168,
-47.7474975585938,
-18.6658744812012,
-46.7095222473145,
-22.7205505371094,
34.7046928405762,
24.7271728515625,
31.0857276916504,
37.9286346435547,
-4.14416408538818,
13.2799072265625,
-23.2130489349365,
37.7560577392578,
22.4658241271973,
-4.16509246826172,
65.4473114013672,
-10.5562458038330,
-13.3673257827759,
51.3626022338867,
40.7392044067383,
-33.8233184814453,
2.41821861267090,
0.569947242736816,
-17.9353904724121,
14.5352687835693,
-42.3444366455078,
46.7861518859863,
10.6205043792725,
-43.7203979492188,
38.1852416992188,
19.3833293914795,
32.0165100097656,
-22.5753269195557,
-4.81531906127930,
37.6030883789063,
-12.2721195220947,
9.50699424743652,
18.1721267700195,
-26.0763549804688,
-19.2130222320557,
13.7181072235107,
-48.9355812072754,
-4.22925567626953,
14.9411859512329,
-6.89974164962769,
59.8492889404297,
-25.8300628662109,
17.5342025756836,
45.5222549438477,
-40.1446723937988,
32.6844787597656,
-2.88664197921753,
-8.42265129089356,
31.7228221893311,
-0.135906860232353,
26.3242092132568,
13.1559076309204,
5.36271619796753,
20.1257743835449,
5.02039670944214,
-0.488026857376099,
13.1959400177002,
1.37157618999481,
29.4831962585449,
48.3143348693848,
-42.1926727294922,
9.09118843078613,
52.9254150390625,
-39.6436042785645,
-13.9332380294800,
-0.473022460937500,
-47.0996284484863,
0.475250244140625,
47.8659706115723,
-6.26073646545410,
0.603926837444305,
32.5293998718262,
5.40081357955933,
14.2449579238892,
-9.61326599121094,
-17.4065971374512,
-15.2772932052612,
-21.9286746978760,
4.12288379669189,
-14.3472661972046,
-44.3122825622559,
-34.5111808776856,
-30.6875724792480,
14.3539505004883,
57.2376899719238,
-8.35751342773438,
-0.979270935058594,
21.3486595153809,
23.8143749237061,
56.6580657958984,
45.4519920349121,
23.7956066131592,
-21.4542160034180,
56.7522506713867,
64.3101501464844,
-11.0718269348145,
-7.66575813293457,
-35.0232543945313,
-10.6946792602539,
-49.4741821289063,
-4.65221977233887,
23.7376327514648,
-69.1720275878906,
11.0762434005737,
16.9254570007324,
-26.6409893035889,
-21.7415981292725,
32.8380279541016,
54.1147193908691,
-47.7621536254883,
-7.52862548828125,
-21.0130634307861,
-8.73612403869629,
39.3376083374023,
11.6505947113037,
4.76897287368774,
-46.0137901306152,
21.7458915710449,
-25.8036918640137,
-5.94349288940430,
83.4870147705078,
21.1643600463867,
20.8538532257080,
14.3611469268799,
-9.23662662506104,
-20.8528652191162,
54.4459800720215,
47.4449462890625,
34.1673278808594,
33.0324935913086,
20.2593059539795,
73.0495300292969,
8.30389404296875,
-37.6051559448242,
-11.7539072036743,
1.98615288734436,
-43.4085998535156,
-43.0327682495117,
51.3868026733398,
51.6519432067871,
-16.3080272674561,
-6.28934288024902,
41.4844512939453,
50.3456115722656,
10.8869876861572,
14.6771640777588,
63.7767486572266,
-33.5406723022461,
25.8602275848389,
80.9646148681641,
-45.0321121215820,
47.1091079711914,
-2.13003540039063,
-19.8392486572266,
38.7585334777832,
-39.4454650878906,
55.1069602966309,
11.0469875335693,
-4.46796369552612,
70.2733688354492,
-21.4773941040039,
32.5807418823242,
37.2367210388184,
-38.5102157592773,
23.9027423858643,
13.3703184127808,
16.4835815429688,
40.9890747070313,
-14.2778015136719,
-8.66870403289795,
-25.0674247741699,
-2.05811405181885,
40.1817283630371,
-0.0442290306091309,
29.0951042175293,
39.5925979614258,
47.2881355285645,
38.5919151306152,
23.4686737060547,
40.7645416259766,
3.10760068893433,
48.7010688781738,
29.7902030944824,
-25.6128997802734,
-2.77946901321411,
16.0744590759277,
49.8974342346191,
-43.3972511291504,
-5.83632469177246,
50.8523483276367,
-23.9693489074707,
-17.9442062377930,
-14.3423318862915,
58.9714317321777,
-16.1765441894531,
-25.2111549377441,
43.5145111083984,
-44.5500602722168,
41.6275291442871,
20.2259769439697,
-50.1816291809082,
34.0495033264160,
-7.87063503265381,
6.77744436264038,
42.2947959899902,
-10.2891254425049,
38.8826942443848,
0.852749824523926,
-3.52370262145996,
62.5221900939941,
-9.47899627685547,
26.4942646026611,
32.6396942138672,
9.06642055511475,
24.2417240142822,
-1.02466177940369,
55.4324188232422,
23.6473617553711,
3.54494905471802,
26.1636562347412,
3.38430976867676,
-47.3013648986816,
6.28187322616577,
12.6751880645752,
-39.5872955322266,
55.2886199951172,
-40.9617691040039,
-3.38004302978516,
85.0200653076172,
-5.29747676849365,
4.30525112152100,
55.5704574584961,
7.18205070495606,
-7.88472604751587,
24.2860679626465,
-30.2275943756104,
23.2112693786621,
-23.5838508605957,
-52.9509468078613,
33.6718139648438,
58.9451522827148,
-18.1716461181641,
-22.1743640899658,
52.3735275268555,
-33.6087150573731,
26.4846744537354,
63.6016540527344,
-15.3199157714844,
6.52515697479248,
20.1399765014648,
-17.3991050720215,
-39.2080307006836,
30.5553474426270,
60.9258537292481,
-20.3459682464600,
-16.4359016418457,
67.0590820312500,
29.5965442657471,
12.2026824951172,
41.2554512023926,
-14.1432094573975,
-10.2373838424683,
24.8253707885742,
6.90668153762817,
27.0553779602051,
-1.20622444152832,
-17.7882728576660,
34.5505790710449,
-44.9364776611328,
5.88997745513916,
78.3458480834961,
-55.9749832153320,
24.3820476531982,
39.1803703308106,
-52.7964591979981,
28.1380863189697,
15.9965982437134,
7.28347492218018,
-5.24520874023438e-05,
2.44548082351685,
58.5624580383301,
7.58866310119629,
-28.2416610717773,
44.5398178100586,
62.1558799743652,
-32.0196037292481,
14.6253070831299,
8.38657760620117,
-34.4373435974121,
21.3296699523926,
-16.0315799713135,
49.2380104064941,
-21.7039813995361,
-55.0331153869629,
79.3292083740234,
4.97198486328125,
-8.96997642517090,
-32.8391342163086,
-7.68074798583984,
42.7522773742676,
6.45490646362305,
43.0290031433106,
43.9114227294922,
50.8724479675293,
-36.7254791259766,
32.9467391967773,
72.2646942138672,
-15.1704168319702,
78.3201675415039,
12.2911367416382,
31.8516921997070,
52.0541534423828,
-23.5670471191406,
48.1957817077637,
-6.16744613647461,
-42.7458686828613,
38.7667655944824,
42.0307350158691,
43.6992645263672,
28.3268089294434,
-13.2669076919556,
67.8993377685547,
30.6442985534668,
-50.2960700988770,
0.0873841643333435,
-24.5153713226318,
-14.0108776092529,
-24.1749763488770,
7.56577682495117,
22.5447044372559,
-9.94483184814453,
32.7992095947266,
-2.60120487213135,
-17.7933158874512,
37.7446327209473,
49.6396789550781,
5.15791130065918,
37.4896278381348,
1.71164512634277,
21.1382808685303,
47.5519371032715,
-39.3178901672363,
30.2061119079590,
31.8443679809570,
-42.0756301879883,
11.0382404327393,
24.7708206176758,
-39.8482551574707,
-4.29037094116211,
39.3930015563965,
-2.42351150512695,
-68.7966308593750,
16.8314933776855,
9.78877258300781,
-41.6970252990723,
43.2509613037109,
-36.4400100708008,
-30.6162548065186,
33.8881721496582,
25.6235694885254,
0.808606982231140,
8.28084373474121,
4.58792114257813,
16.9293842315674,
55.3445625305176,
-12.3806886672974,
-12.3232793807983,
-2.73931694030762,
18.6195030212402,
35.9051666259766,
26.4373512268066,
-10.1325864791870,
1.41694450378418,
73.6630706787109,
16.4445533752441,
42.7449264526367,
45.4452705383301,
-21.0216140747070,
40.6261672973633,
59.2742843627930,
6.59646368026733,
-3.08896303176880,
-8.98358535766602,
-17.4028282165527,
31.0415687561035,
27.8298950195313,
-6.05901908874512,
-50.9151763916016,
-23.2293663024902,
44.3111991882324,
27.8584785461426,
25.0539703369141,
12.2990989685059,
31.9335613250732,
-22.0221366882324,
-6.36846923828125,
32.2563133239746,
-10.2829551696777,
27.4562625885010,
-14.5529279708862,
37.2259407043457,
11.5798339843750,
-53.2106628417969,
53.1499137878418,
58.0661087036133,
9.93860721588135,
-26.3779296875000,
12.9463729858398,
56.5926818847656,
41.2321395874023,
31.5722732543945,
12.2718734741211,
34.4815101623535,
40.5347671508789,
10.8310031890869,
31.1033020019531,
4.05751228332520,
-28.6999740600586,
6.97675275802612,
-12.0452985763550,
-15.8655729293823,
11.6122531890869,
-36.8416481018066,
-7.16117382049561,
43.3490715026856,
-14.7664127349854,
-14.2988662719727,
-2.17771005630493,
-2.16675543785095,
-17.7538070678711,
-18.3226165771484,
36.5393066406250,
26.9790534973145,
-42.9626655578613,
-19.0290641784668,
70.7698059082031,
-15.9901628494263,
-21.9042358398438,
46.9495277404785,
-7.89014720916748,
12.0773735046387,
18.8268222808838,
60.8727569580078,
12.3581733703613,
-20.0102863311768,
6.63863277435303,
-31.4128112792969,
57.1502037048340,
-25.6599025726318,
2.44600677490234,
51.4555740356445,
-58.5830459594727,
-13.0644302368164,
46.0562591552734,
24.7848815917969,
-34.8827667236328,
54.8959465026856,
-10.1959037780762,
-54.3768310546875,
19.5572185516357,
11.9776630401611,
6.93077039718628,
-61.0096511840820,
3.51494979858398,
62.5551300048828,
5.75577545166016,
-2.44276189804077,
63.6260643005371,
50.9855957031250,
26.0536155700684,
44.4988708496094,
11.0520935058594,
42.8785781860352,
41.0787544250488,
17.4143371582031,
-15.8991670608521,
-8.73325061798096,
44.1313896179199,
23.9367942810059,
13.4466571807861,
6.23530912399292,
-2.18952274322510,
-19.0042705535889,
62.8088340759277,
9.18682289123535,
-13.0960474014282,
19.8888530731201,
-39.5132064819336,
48.3556175231934,
-0.906830787658691,
-11.9099407196045,
7.92272424697876,
-29.7498836517334,
6.80413055419922,
73.3303833007813,
-17.7199020385742,
-6.36035156250000,
56.9595260620117,
-56.1044235229492,
24.3276271820068,
16.1315250396729,
37.4315528869629,
-8.49294471740723,
-60.6843261718750,
-6.28747320175171,
-24.7153091430664,
25.7702369689941,
-42.7413139343262,
-7.86991405487061,
42.0550003051758,
-33.4701957702637,
-25.6408863067627,
-2.12179160118103,
-27.4394893646240,
16.9409885406494,
52.8690452575684,
23.3502998352051,
59.2500534057617,
17.6759147644043,
14.6795635223389,
39.8547439575195,
18.1913757324219,
34.2678680419922,
17.3235473632813,
-8.56800079345703,
15.7770261764526,
51.5631408691406,
-16.2027702331543,
-8.16879177093506,
-31.8770446777344,
0.502490997314453,
20.2716045379639,
-30.5508403778076,
45.0104675292969,
-28.5775833129883,
13.9921493530273,
35.2070999145508,
9.85597801208496,
-4.98117494583130,
27.6230335235596,
29.8096961975098,
-42.9511642456055,
56.1249771118164,
-24.3211822509766,
10.0471897125244,
21.7940349578857,
-3.59499645233154,
-3.59946250915527,
-37.9339637756348,
62.1346054077148,
1.59973621368408,
10.7052850723267,
4.36821651458740,
-1.50428676605225,
40.7116889953613,
31.8988685607910,
57.1227302551270,
26.9049644470215,
5.46215438842773,
-16.9542350769043,
31.8118591308594,
11.7673435211182,
-37.3107872009277,
27.8841857910156,
32.7862777709961,
-30.2771301269531,
-15.4783773422241,
58.0489273071289,
40.5601692199707,
16.6547164916992,
-19.8195476531982,
42.6383132934570,
20.7755126953125,
-28.3089561462402,
39.2761001586914,
24.2874050140381,
41.8355178833008,
47.6801338195801,
57.2555618286133,
-14.9610385894775,
46.1210708618164,
42.8870544433594,
9.06472015380859,
46.6953620910645,
-8.01142883300781,
69.9789199829102,
-60.5917625427246,
-7.90622568130493,
66.3150329589844,
-62.6046981811523,
15.6946945190430,
38.0355339050293,
15.1172561645508,
-6.31462860107422,
-10.0477619171143,
4.14579677581787,
38.2283325195313,
12.2628526687622,
-1.07930302619934,
45.8750190734863,
8.83399295806885,
29.0982589721680,
-9.88755798339844,
21.7651653289795,
66.1857299804688,
-4.58570766448975,
39.8821640014648,
13.7958021163940,
-4.51390409469605,
28.3173904418945,
-10.5141801834106,
-38.6068763732910,
39.7475547790527,
4.07935714721680,
-23.6594390869141,
86.8379211425781,
-11.5767250061035,
-4.68504619598389,
0.186466693878174,
2.49040770530701,
50.1861305236816,
-29.5835819244385,
51.4830436706543,
32.8502807617188,
5.28242254257202,
16.7093811035156,
-13.7055301666260,
-27.2310562133789,
-19.0586624145508,
-12.1074562072754,
-39.6957054138184,
-9.79982852935791,
-37.4180679321289,
16.8210182189941,
-22.2713203430176,
-54.2396583557129,
-26.7531852722168,
-7.65318679809570,
42.5414390563965,
4.99512338638306,
20.4038734436035,
-9.04498767852783,
33.1942672729492,
20.1418056488037,
27.9924316406250,
57.9694175720215,
-48.3690071105957,
17.7256164550781,
30.4027309417725,
-11.6599712371826,
24.1588649749756,
-15.3228187561035,
-9.26505279541016,
14.8399562835693,
-2.30404853820801,
-10.0702304840088,
-39.1175842285156,
-14.9486503601074,
0.297442078590393,
-36.2078399658203,
-7.16926765441895,
31.6358547210693,
9.62985324859619,
1.37944376468658,
57.7093772888184,
40.5001411437988,
-32.1684494018555,
5.74004077911377,
9.02994251251221,
12.2619562149048,
65.2378158569336,
23.1267814636230,
-17.5207881927490,
-28.5307483673096,
-10.0515613555908,
8.33635044097900,
-17.7262096405029,
-4.20966339111328,
24.5932598114014,
6.89366722106934,
6.38217353820801,
23.6455459594727,
31.5446090698242,
9.44609069824219,
-13.0946464538574,
43.9342269897461,
62.0979309082031,
34.7643165588379,
50.3047637939453,
-1.08681106567383,
1.02048015594482,
48.4553489685059,
-20.5277214050293,
-1.88287270069122,
6.20572566986084,
-14.3646717071533,
-24.9246959686279,
-34.9405822753906,
55.8517227172852,
8.96819877624512,
-47.8204803466797,
-3.81609249114990,
-13.9618225097656,
-49.9734420776367,
10.3034696578980,
22.7483768463135,
-22.3837814331055,
2.41521120071411,
-31.6369762420654,
-7.83692836761475,
-26.5973415374756,
-32.2293014526367,
-2.52667331695557,
-11.2271881103516,
57.8510246276856,
18.0356140136719,
26.6807289123535,
3.91783857345581,
-29.4631099700928,
45.7212753295898,
7.81591749191284,
-13.3397321701050,
-27.1560745239258,
10.6904582977295,
1.47758865356445,
-10.2429695129395,
64.2927780151367,
35.6787986755371,
0.683951854705811,
-41.9802780151367,
18.3695621490479,
59.3341941833496,
4.23539352416992,
47.3272171020508,
50.9533958435059,
-16.9056205749512,
-34.5305252075195,
41.2799110412598,
50.6938438415527,
34.3744850158691,
17.1717128753662,
-23.5206031799316,
11.2350311279297,
52.7068405151367,
65.9984207153320,
-9.53205680847168,
20.7638549804688,
71.7770080566406,
-12.3714122772217,
-23.9736003875732,
12.0621109008789,
18.6909141540527,
18.3045120239258,
-4.16358566284180,
-24.2137718200684,
54.1789665222168,
32.7304725646973,
-14.5582065582275,
27.3641433715820,
21.1227741241455,
37.3715782165527,
-5.38302803039551,
-25.7779159545898,
18.2387847900391,
-11.5115947723389,
14.6914157867432,
47.2682037353516,
-17.0041484832764,
-40.0962066650391,
-2.75173950195313,
30.9205017089844,
43.2605476379395,
20.0496330261230,
10.5589923858643,
43.7084732055664,
-19.3435859680176,
-36.3677215576172,
41.9924850463867,
-25.3491477966309,
10.2498073577881,
25.4292125701904,
4.49791049957275,
52.7683639526367,
-40.5804214477539,
49.1389236450195,
54.4101219177246,
-53.8632774353027,
36.0935783386231,
-12.6975841522217,
-21.6617164611816,
46.4564590454102,
-11.9886913299561,
18.7111797332764,
52.2631416320801,
20.6568279266357,
-3.07811951637268,
17.6497383117676,
61.0418739318848,
0.167764663696289,
-26.7595367431641,
31.7814140319824,
53.3331069946289,
-13.4730472564697,
4.16577148437500,
23.3334465026855,
17.2401943206787,
37.5371475219727,
-15.9717979431152,
15.0346622467041,
51.0956535339356,
38.0448608398438,
-12.2498769760132,
11.1885128021240,
54.2228698730469,
19.8788909912109,
40.1024703979492,
60.6668624877930,
39.6972427368164,
20.0215244293213,
44.6414070129395,
18.2719097137451,
47.3508453369141,
49.6432800292969,
-5.81956195831299,
40.1951637268066,
-15.4934711456299,
-19.8412151336670,
17.3586521148682,
19.3649578094482,
54.0169906616211,
-7.90540170669556,
33.5855026245117,
45.7275695800781,
-38.1795578002930,
15.8607225418091,
0.344692230224609,
-20.5832977294922,
-10.7072687149048,
-37.5921058654785,
-14.1998138427734,
-19.2525405883789,
10.5053310394287,
14.9982881546021,
-34.0773353576660,
21.1873092651367,
67.6774826049805,
-20.5349922180176,
-20.2361202239990,
7.16465663909912,
2.72274351119995,
49.6996612548828,
6.14445209503174,
-9.95526409149170,
37.8496017456055,
23.2299079895020,
-26.3931045532227,
-13.9122295379639,
-15.7524852752686,
-10.5245389938355,
-9.88188552856445,
-37.0771255493164,
-26.9685630798340,
29.0335445404053,
13.2391967773438,
-34.1211967468262,
42.8688964843750,
4.18993520736694,
31.4317855834961,
-4.71021080017090,
-11.9450988769531,
78.5832138061523,
-12.0581569671631,
-6.02549409866333,
-8.46936798095703,
18.2504653930664,
-30.9386520385742,
17.4858741760254,
71.1955947875977,
-38.1828613281250,
46.9437370300293,
15.9196014404297,
-28.5256118774414,
-16.2128505706787,
2.93330121040344,
54.8353805541992,
18.2426815032959,
48.6431999206543,
15.2280044555664,
-22.8518447875977,
-8.80481624603272,
-25.8870162963867,
24.0797901153564,
10.2608203887939,
-48.5677757263184,
-25.1225490570068,
47.0194854736328,
-19.1677932739258,
-41.4555892944336,
-7.19482040405273,
-70.0932006835938,
36.7416839599609,
16.2286262512207,
-21.6878852844238,
-0.558053016662598,
-17.7233734130859,
-3.01842164993286,
-37.1032257080078,
62.6856460571289,
19.3798999786377,
22.3590316772461,
60.6354446411133,
37.0266838073731,
12.6032142639160,
-10.0780086517334,
46.6671524047852,
-40.1785392761231,
77.2188568115234,
43.1620292663574,
-67.2040176391602,
53.3260841369629,
3.65511941909790,
30.6900253295898,
6.39356708526611,
-22.6032829284668,
47.3899803161621,
36.3132171630859,
23.5337638854980,
33.7684898376465,
43.7007598876953,
-42.9641342163086,
6.36988067626953,
28.4659252166748,
-12.3323907852173,
20.7103748321533,
-43.3633804321289,
-3.01361083984375,
-1.41540670394897,
39.8974990844727,
39.3991432189941,
-12.1620569229126,
54.1856918334961,
-3.09650206565857,
38.7765350341797,
35.4020805358887,
25.0862445831299,
67.9015426635742,
35.7830085754395,
-2.16954517364502,
-14.2345104217529,
68.2442703247070,
3.19167900085449,
1.14297056198120,
66.0236663818359,
30.9463367462158,
23.4572963714600,
-4.17574882507324,
-1.39844703674316,
69.6704330444336,
-9.62321090698242,
-30.0351409912109,
60.5336456298828,
24.3506946563721,
29.2727012634277,
-10.7492733001709,
-19.4065208435059,
2.14566135406494,
41.3360824584961,
-5.61878395080566,
-6.64312839508057,
45.3390655517578,
37.7182121276856,
14.9909219741821,
-17.6225948333740,
49.2982940673828,
-11.4405059814453,
39.8478088378906,
-7.46088600158691,
0.268075942993164,
33.7129859924316,
-72.2326354980469,
13.4945745468140,
15.1316652297974,
56.6217002868652,
23.6150436401367,
12.4557418823242,
32.4647903442383,
-43.5012969970703,
9.59316253662109,
56.5478172302246,
53.6722412109375,
20.9892539978027,
-24.2156887054443,
14.5666589736938,
50.3830413818359,
0.166639089584351,
-11.5676689147949,
14.0305299758911,
40.0753211975098,
-12.0708465576172,
-34.2615852355957,
-0.908643245697022,
-32.0766181945801,
-3.77562427520752,
-7.30662488937378,
34.1491279602051,
39.2474441528320,
-24.4045467376709,
7.88256549835205,
-10.2844200134277,
41.2469139099121,
43.2795333862305,
-14.5394315719605,
-1.66813445091248,
15.3674039840698,
5.28538894653320,
-43.6829910278320,
-0.889256358146668,
-4.48597908020020,
-22.7144393920898,
-19.0906467437744,
-24.8249759674072,
-7.75997495651245,
12.6171550750732,
20.6876525878906,
-46.1669692993164,
-12.6614465713501,
29.1894397735596,
-23.7489948272705,
-16.7260780334473,
37.0625839233398,
41.0012817382813,
-6.17725086212158,
12.2765731811523,
31.8569908142090,
-1.45195794105530,
17.0394668579102,
17.6451778411865,
-8.84281635284424,
-41.8516921997070,
-6.97704601287842,
14.8483524322510,
-46.0767898559570,
35.9238929748535,
30.0182304382324,
16.1734600067139,
37.4322776794434,
1.03505063056946,
60.9480667114258,
7.52219963073731,
-13.7039747238159,
-10.9897012710571,
12.1585397720337,
66.4733352661133,
4.94973564147949,
-12.2229251861572,
9.43649864196777,
48.4492416381836,
3.27764034271240,
-10.4379329681396,
18.4759445190430,
-6.85511779785156,
50.4113998413086,
3.36547422409058,
5.99974632263184,
61.6230392456055,
-3.79806995391846,
2.93717956542969,
23.5626659393311,
25.4963550567627,
35.1112747192383,
29.2387981414795,
-41.4573478698731,
-23.6567077636719,
-4.29820919036865,
-37.0268478393555,
-12.0729522705078,
-40.7132415771484,
42.0533294677734,
17.2030372619629,
10.5674772262573,
42.6962242126465,
-14.9034709930420,
33.6147727966309,
-17.0073585510254,
7.69874191284180,
36.0408821105957,
32.2382621765137,
46.1223831176758,
61.8036804199219,
11.5272216796875,
-25.2682037353516,
59.0549812316895,
0.505073547363281,
54.6262359619141,
38.9384117126465,
-17.0198364257813,
48.1843566894531,
12.8820190429688,
28.1990947723389,
51.2850112915039,
-12.6388988494873,
-35.5771255493164,
7.36762857437134,
4.75117349624634,
2.11906909942627,
8.41848278045654,
-8.65665912628174,
-33.7769622802734,
-15.4710912704468,
-2.64371109008789,
-11.9372997283936,
-34.7432899475098,
-20.8178100585938,
60.4712104797363,
0.617988348007202,
-39.5178337097168,
23.5764389038086,
15.7063760757446,
30.6871967315674,
14.6711616516113,
36.6848640441895,
29.1123905181885,
-65.1761627197266,
17.2831783294678,
-23.1384201049805,
-27.2799015045166,
34.7353286743164,
-26.5506801605225,
8.42971229553223,
-40.7642936706543,
13.2151584625244,
-7.71695613861084,
-25.6723556518555,
50.5709457397461,
-64.9269256591797,
-13.4820432662964,
23.7488536834717,
2.46204233169556,
36.6466827392578,
38.3526573181152,
-14.3658237457275,
-52.4386558532715,
36.1204643249512,
7.29307556152344,
-56.9271163940430,
-14.2452983856201,
11.0459499359131,
-18.1590175628662,
-22.7183570861816,
36.1443519592285,
29.6398010253906,
-10.2794113159180,
-9.55071544647217,
0.738215446472168,
34.6798248291016,
34.2615928649902,
53.6524467468262,
7.11969280242920,
-23.2966632843018,
45.9217910766602,
-33.2363243103027,
-29.8604679107666,
-5.97416019439697,
-44.4105262756348,
38.9597358703613,
14.1108341217041,
-55.7085914611816,
-11.5247039794922,
41.3049430847168,
-37.2046546936035,
-44.9656791687012,
23.7314624786377,
15.7554397583008,
21.1526489257813,
2.95313453674316,
57.9180107116699,
-11.8499565124512,
-20.9190711975098,
38.9309692382813,
-15.1925849914551,
-42.4719085693359,
-21.1561851501465,
51.9361534118652,
-45.3435859680176,
20.5039672851563,
20.0174198150635,
-29.2104988098145,
20.0312500000000,
-45.0646972656250,
-30.7954616546631,
-28.6244812011719,
-4.96050739288330,
-18.6091442108154,
0.710431098937988,
8.00843620300293,
-3.13265538215637,
-20.2117271423340,
-6.79306888580322,
-10.4471111297607,
19.3169174194336,
38.7183914184570,
17.0217475891113,
49.4938697814941,
-30.5651893615723,
58.3028030395508,
16.9212512969971,
-13.6609077453613,
48.2562828063965,
25.8699913024902,
9.51906776428223,
-50.3900260925293,
13.7646598815918,
15.7938766479492,
-39.6957015991211,
35.2031822204590,
55.5980186462402,
-60.9371795654297,
5.02631378173828,
-0.852302551269531,
-6.01531982421875,
52.4838256835938,
-34.2873268127441,
-31.9456520080566,
12.4339389801025,
52.1856727600098,
-15.4421472549438,
16.2738304138184,
55.1174583435059,
25.9313774108887,
12.6940040588379,
-42.1607208251953,
58.0806236267090,
7.46574020385742,
-26.8170871734619,
21.4817657470703,
-33.9222450256348,
34.3561058044434,
-27.4372253417969,
-24.4412555694580,
74.3348617553711,
0.571651458740234,
23.7039299011230,
7.24145698547363,
-28.2240295410156,
27.7118949890137,
-36.1059226989746,
-30.0788364410400,
17.9792041778564,
-45.9245223999023,
-48.3527603149414,
12.9879150390625,
49.2779388427734,
-35.9426002502441,
-7.72062301635742,
44.2627143859863,
-68.4912185668945,
-21.2829399108887,
-12.6457901000977,
18.4586238861084,
52.8295974731445,
-49.0592918395996,
10.1219959259033,
14.9462413787842,
20.5673999786377,
26.2207813262939,
-12.2933549880981,
81.9750213623047,
41.2768821716309,
-1.01050901412964,
1.53874111175537,
-9.58118152618408,
-13.3459119796753,
-27.3874931335449,
61.1988258361816,
-17.2245006561279,
-20.1966629028320,
30.4782562255859,
-50.6470375061035,
50.9970855712891,
18.2797508239746,
-36.6529655456543,
-4.98466444015503,
-7.30398416519165,
30.1641426086426,
8.57611465454102,
43.7655487060547,
15.9899559020996,
-11.0736484527588,
-9.90065383911133,
8.29669570922852,
-6.64432001113892,
-45.5251350402832,
31.0511627197266,
-28.7607803344727,
-16.5439872741699,
-8.21274280548096,
-4.81267929077148,
22.0162887573242,
-12.1986141204834,
44.9137496948242,
-14.1848926544189,
-23.1175003051758,
-18.7975234985352,
21.9675407409668,
54.4303512573242,
31.3315505981445,
62.8547363281250,
4.92932605743408,
11.1257228851318,
55.5017395019531,
2.22431850433350,
-30.5081043243408,
71.4795837402344,
32.1035804748535,
-2.83839821815491,
50.9213790893555,
30.1620159149170,
50.6723976135254,
-51.4257545471191,
20.9434204101563,
29.7811126708984,
-40.9890899658203,
77.4582138061523,
15.0407133102417,
20.7325553894043,
58.4902763366699,
23.3651237487793,
21.8485813140869,
51.1042938232422,
-18.1617393493652,
3.00655937194824,
77.0309448242188,
1.28707504272461,
19.1968288421631,
9.06449890136719,
-3.70057201385498,
-21.3506927490234,
8.50639343261719,
25.2692337036133,
26.3610458374023,
5.26911401748657,
-3.74435806274414,
95.7767639160156,
-7.80250740051270,
6.36827278137207,
59.7174377441406,
0.0151785016059875,
59.8542022705078,
-21.6414718627930,
-33.8546562194824,
41.4579277038574,
44.6052513122559,
23.8790740966797,
-43.3541259765625,
-8.83478450775147,
-6.49578475952148,
-3.35422611236572,
36.5490875244141,
16.0924129486084,
-11.3257656097412,
-36.2789192199707,
-25.7741508483887,
-19.3266162872314,
-11.1142139434814,
-5.40610122680664,
30.3933296203613,
23.8364276885986,
-20.0772075653076,
29.7185592651367,
64.0181427001953,
29.7335090637207,
-36.3110160827637,
-27.2428817749023,
38.3909606933594,
64.1088943481445,
-10.5472030639648,
-1.41755485534668,
58.6883239746094,
-45.4578628540039,
-0.335154533386230,
46.9155273437500,
-17.1671085357666,
-10.1737718582153,
-40.2443275451660,
-18.0378646850586,
40.8572387695313,
22.9782257080078,
21.1550655364990,
-12.9449748992920,
11.6719408035278,
55.0538864135742,
-11.9820022583008,
35.0673866271973,
65.4834442138672,
7.64607715606689,
-13.0834426879883,
16.3202476501465,
18.8708934783936,
50.4155883789063,
18.2318305969238,
30.7654876708984,
26.4517250061035,
-42.3118896484375,
67.9607620239258,
-17.0117683410645,
-2.08905220031738,
15.8068008422852,
7.12762928009033,
39.4089813232422,
-3.48019552230835,
66.3302917480469,
-15.2909650802612,
-21.6112155914307,
-10.5996570587158,
18.0285644531250,
40.8086776733398,
28.0824661254883,
29.2431335449219,
-12.8631381988525,
25.3658065795898,
-48.4265289306641,
-1.21865558624268,
71.1315841674805,
14.4501075744629,
-30.6410961151123,
-34.7014122009277,
15.5749206542969,
6.41911697387695,
48.3608665466309,
12.8067531585693,
27.8708419799805,
-3.68003082275391,
-27.4514808654785,
61.4807510375977,
-28.7158489227295,
16.7709503173828,
-0.841584920883179,
20.4963016510010,
43.8208999633789,
-13.4274578094482,
101.121688842773,
-19.7493648529053,
-26.8751945495605,
59.5849418640137,
18.8064765930176,
41.9382019042969,
18.6683464050293,
-28.0287857055664,
-14.9825611114502,
48.3762283325195,
-41.8445281982422,
15.9526252746582,
50.9305038452148,
-31.2655982971191,
54.8016281127930,
28.0279674530029,
47.4476699829102,
52.8559494018555,
20.7488059997559,
51.2871551513672,
39.4036140441895,
11.7993555068970,
8.41510105133057,
43.9813041687012,
48.6583900451660,
-5.03049564361572,
-8.91366195678711,
49.8005065917969,
29.6088771820068,
39.5255012512207,
9.27184963226318,
-9.33020591735840,
51.6073379516602,
-26.7527294158936,
-10.5440120697021,
83.0868835449219,
-3.29221057891846,
-0.143053293228149,
59.9168395996094,
18.9736785888672,
3.75962924957275,
-1.14029598236084,
23.4686107635498,
-11.3029117584229,
-48.9794387817383,
25.3662548065186,
40.0161972045898,
-25.4613494873047,
-4.20522975921631,
-8.55454063415527,
-20.1917839050293,
36.5768966674805,
-2.61530709266663,
9.93250942230225,
-25.8314437866211,
8.28170013427734,
67.2440338134766,
21.7616443634033,
36.0244407653809,
-6.79278993606567,
10.0632467269897,
6.20570945739746,
-8.10578346252441,
-2.59169197082520,
0.109176158905029,
15.6870489120483,
37.7852325439453,
14.2694683074951,
-5.95447015762329,
32.2352294921875,
-42.0951614379883,
-32.8678932189941,
36.1378097534180,
-12.7608499526978,
-35.0469322204590,
24.9263687133789,
27.6546020507813,
22.4708671569824,
-12.5799980163574,
-5.70275497436523,
17.6919746398926,
-27.5868415832520,
5.23037195205689,
-26.8706150054932,
6.52287244796753,
-16.8254776000977,
-45.0017585754395,
29.2693710327148,
-12.1150455474854,
31.6899642944336,
6.61652040481567,
-0.651583194732666,
30.3469638824463,
14.6325416564941,
23.9176254272461,
-37.2891960144043,
46.8914871215820,
37.8889045715332,
9.32285785675049,
65.7903747558594,
-3.41217994689941,
-3.33236360549927,
10.4638843536377,
-8.06269168853760,
7.61867332458496,
29.0413780212402,
-37.7328262329102,
-14.1280136108398,
29.6544742584229,
-41.4792442321777,
1.96800518035889,
5.58008909225464,
-29.4727706909180,
21.0608444213867,
-21.5399570465088,
37.7199058532715,
58.9105682373047,
-50.6276931762695,
12.2833919525146,
-19.9146575927734,
13.4718399047852,
59.8832168579102,
10.5273284912109,
-22.3820362091064,
-18.5038738250732,
31.1543159484863,
-5.61059761047363,
27.2470550537109,
53.6004638671875,
56.1341018676758,
-7.05980777740479,
22.5393867492676,
-3.71584224700928,
-3.05378532409668,
35.0813903808594,
-28.4835605621338,
19.9768962860107,
-7.25075101852417,
26.1858520507813,
-24.9344711303711,
3.55031108856201,
-0.308858871459961,
-54.9403152465820,
25.3947200775147,
33.8145256042481,
-7.11184024810791,
-29.7266578674316,
59.8116950988770,
-11.8485393524170,
-40.9404678344727,
41.2546043395996,
61.4079780578613,
3.92494869232178,
-5.08386421203613,
14.5293579101563,
18.5421066284180,
35.7678565979004,
26.7964553833008,
8.53739070892334,
-34.2629547119141,
7.43343782424927,
-35.9800148010254,
16.1507778167725,
21.4740619659424,
-26.3186168670654,
33.6065216064453,
42.4329681396484,
30.4216880798340,
-32.6961288452148,
54.8789939880371,
51.8341598510742,
-47.4480247497559,
22.7079410552979,
10.4865846633911,
-24.5294322967529,
55.6331329345703,
-8.44861984252930,
-17.1769371032715,
67.3121414184570,
-50.0504074096680,
-28.2701187133789,
17.3676986694336,
-15.6071805953980,
39.4983406066895,
2.82637071609497,
10.6843719482422,
2.42690849304199,
-25.1379203796387,
25.4387474060059,
30.6197071075439,
-5.13584184646606,
-28.9529323577881,
19.1627655029297,
31.3371143341064,
39.1024208068848,
-12.5694751739502,
-63.3389816284180,
41.7448120117188,
43.6523628234863,
24.0789966583252,
52.3167495727539,
12.2107725143433,
14.5624389648438,
-15.2023096084595,
-18.9466648101807,
73.5632476806641,
41.1077079772949,
18.0365295410156,
28.8977012634277,
-28.7597904205322,
26.4292831420898,
26.5086841583252,
-7.88343620300293,
19.7163677215576,
-20.2349395751953,
-27.6263675689697,
-19.9549732208252,
1.77148795127869,
-10.6910696029663,
-8.20855712890625,
5.73906135559082,
-53.5072059631348,
3.38081836700439,
28.3817501068115,
22.5541343688965,
45.8393249511719,
-8.04967117309570,
43.3196449279785,
-0.580659866333008,
-56.6925544738770,
44.3570671081543,
-8.96554756164551,
-2.17770481109619,
37.0277175903320,
0.281299740076065,
16.3502044677734,
27.3951454162598,
3.92763948440552,
-19.3254470825195,
43.6498565673828,
42.7640686035156,
30.7880687713623,
-5.95878744125366,
4.15773010253906,
37.5940284729004,
-13.1934633255005,
4.93120098114014,
43.4559516906738,
52.7258377075195,
-27.9012031555176,
13.3695964813232,
-6.76885986328125,
-27.4415740966797,
54.0637588500977,
-5.20655584335327,
-7.19747734069824,
34.6365547180176,
24.6147708892822,
-32.5442123413086,
28.5457477569580,
27.5558376312256,
35.2844200134277,
15.2483654022217,
-63.5779876708984,
71.8949508666992,
-7.22800445556641,
-18.8634166717529,
13.4583501815796,
-33.8838043212891,
61.9272193908691,
-40.4643859863281,
-38.8253631591797,
50.5402412414551,
-19.0713996887207,
-69.4647903442383,
27.1602210998535,
56.7431983947754,
-14.3205099105835,
33.0027542114258,
12.7034044265747,
23.3743476867676,
14.2592926025391,
19.1663837432861,
65.4763946533203,
-16.1953659057617,
-26.3719711303711,
-5.54941082000732,
-40.3308792114258,
-1.85971260070801,
72.6492462158203,
20.3487167358398,
-54.0595855712891,
41.0305366516113,
46.7879104614258,
-11.5148401260376,
55.3433074951172,
-16.6081657409668,
20.5840263366699,
49.1836585998535,
24.2097549438477,
19.7988624572754,
-27.4542827606201,
53.3619689941406,
2.34988403320313,
19.5098609924316,
-7.65693283081055,
-12.5639667510986,
45.5470657348633,
-27.5249309539795,
-26.1259021759033,
-42.4827995300293,
-22.1194114685059,
-31.0367202758789,
5.06190204620361,
56.6603279113770,
-43.6132812500000,
-17.2992248535156,
62.6578216552734,
-2.85422897338867,
31.5736827850342,
24.2967758178711,
-39.3397865295410,
50.5067749023438,
40.7633285522461,
-9.47541046142578,
39.9500923156738,
58.1048812866211,
-21.1058788299561,
10.8291168212891,
88.3154907226563,
14.7328395843506,
25.6967201232910,
46.3788146972656,
-16.7733192443848,
-30.3404159545898,
-11.8522214889526,
-16.0957984924316,
-32.0869674682617,
14.1616353988647,
10.0774250030518,
-11.4216918945313,
50.8002395629883,
38.5929183959961,
-22.9219818115234,
-25.7029247283936,
75.0924453735352,
36.9302444458008,
-57.8267097473145,
21.0756530761719,
14.5423774719238,
24.9573211669922,
53.6532135009766,
37.1717224121094,
7.21488285064697,
53.1872291564941,
47.8656005859375,
38.7694854736328,
42.1807670593262,
-30.7093162536621,
52.2368087768555,
-7.98585033416748,
30.6287708282471,
29.6575088500977,
-7.51071739196777,
32.6748275756836,
-62.5902709960938,
31.7958126068115,
58.7742080688477,
-26.5155448913574,
-36.5402565002441,
62.0278587341309,
11.9547309875488,
-66.2816925048828,
-1.38364863395691,
-24.1896896362305,
-42.6713447570801,
10.3353252410889,
36.1981811523438,
-39.0729446411133,
-29.1142749786377,
1.15723633766174,
-16.2349319458008,
-12.0871791839600,
1.15926170349121,
2.98512458801270,
0.419034957885742,
37.7635879516602,
-4.05006837844849,
1.34229326248169,
61.5929985046387,
-12.1428194046021,
5.26497650146484,
72.3338470458984,
-4.33470344543457,
5.94886779785156,
44.9328880310059,
9.44515132904053,
22.2913837432861,
62.8228454589844,
30.9417304992676,
-7.46039628982544,
62.3028564453125,
11.5408878326416,
-11.0461292266846,
40.1191864013672,
25.9627037048340,
76.8577041625977,
-22.3022994995117,
-0.107315063476563,
56.7240486145020,
-49.6139183044434,
3.75694656372070,
71.6309127807617,
41.7487716674805,
-4.63634252548218,
48.8727035522461,
20.5936203002930,
-32.7476577758789,
-32.6846694946289,
5.81407928466797,
20.6140289306641,
-44.5094490051270,
32.2065010070801,
43.2899093627930,
27.0757446289063,
20.2554798126221,
-28.7841377258301,
-16.7403030395508,
28.1984176635742,
-24.7026157379150,
-20.8210849761963,
46.5168685913086,
-36.6445388793945,
0.880334615707398,
25.8221054077148,
10.5746631622314,
-1.15816044807434,
9.29368495941162,
44.2373695373535,
-16.3952331542969,
15.4014091491699,
-30.1557197570801,
-2.94258022308350,
9.58894920349121,
-8.49825191497803,
57.3402099609375,
-26.1845645904541,
46.6140060424805,
-5.48389816284180,
-41.6608238220215,
54.9613037109375,
-0.598618268966675,
21.7689590454102,
19.7177581787109,
40.5969734191895,
30.4256134033203,
-44.9258193969727,
21.6116523742676,
72.9654922485352,
-40.0724563598633,
8.21716880798340,
45.1730346679688,
-31.3204879760742,
13.6241722106934,
-39.0822944641113,
-9.09269046783447,
1.96258163452148,
-19.5932846069336,
53.0242347717285,
-38.3502006530762,
-5.49081611633301,
20.9981346130371,
-48.6121673583984,
26.3867454528809,
18.0801734924316,
-0.940515995025635,
16.2456111907959,
14.5850152969360,
-12.5241994857788,
5.20542335510254,
48.2844924926758,
-31.4362888336182,
0.827085494995117,
17.0273590087891,
-9.59509277343750,
59.1932830810547,
-9.07495117187500,
22.4300823211670,
50.3071861267090,
-36.6134948730469,
35.9726333618164,
0.506084442138672,
-3.27420616149902,
70.4236602783203,
18.4850368499756,
14.7399120330811,
19.3050174713135,
16.6873798370361,
27.8347358703613,
-18.9438571929932,
-3.97566246986389,
45.8432884216309,
28.9535903930664,
12.2903270721436,
-0.997106313705444,
25.1747550964355,
14.1551942825317,
38.5171966552734,
-6.00951766967773,
-21.3925304412842,
78.6696929931641,
24.2563190460205,
30.9664230346680,
11.7618837356567,
-16.7543296813965,
25.2589988708496,
29.7648258209229,
64.6728363037109,
27.2962112426758,
-4.55389928817749,
44.0064659118652,
56.2836990356445,
35.2863464355469,
28.3039054870605,
23.2136688232422,
20.0746307373047,
43.9641227722168,
59.8526191711426,
44.8371849060059,
26.4124298095703,
-48.0638046264648,
6.94610452651978,
69.6779098510742,
-39.1921043395996,
-14.8753938674927,
36.4751510620117,
39.3339843750000,
-2.09023094177246,
-36.3542366027832,
-5.10976696014404,
-11.6314888000488,
-37.6777000427246,
-4.56389856338501,
65.0687255859375,
-25.7126121520996,
-45.8872375488281,
41.7473297119141,
-3.78791856765747,
-5.06432533264160,
63.1544227600098,
28.8043670654297,
18.4226951599121,
23.2820644378662,
10.8201198577881,
7.72042083740234,
-32.4341735839844,
19.9871368408203,
36.1760215759277,
14.0306091308594,
9.13432121276856,
22.6914825439453,
55.1642189025879,
-25.2905826568604,
-15.4827919006348,
41.5527725219727,
-25.3152160644531,
-41.5774497985840,
24.4452037811279,
31.9664230346680,
-41.8992767333984,
23.2578239440918,
61.4054412841797,
-49.4871253967285,
-10.0973339080811,
27.6529979705811,
17.5681533813477,
42.5351448059082,
16.6274509429932,
18.3156242370605,
11.3603105545044,
3.33495450019836,
-11.2755317687988,
-33.0885810852051,
34.3594093322754,
15.6281070709229,
-13.9022350311279,
2.66451549530029,
1.70642805099487,
3.21772670745850,
-3.43328905105591,
34.0804824829102,
30.3732547760010,
52.2644691467285,
-6.30099201202393,
3.35454750061035,
84.2614135742188,
19.7427864074707,
19.7459163665772,
33.2730979919434,
-20.7297477722168,
-27.6582946777344,
58.5082817077637,
22.5007858276367,
14.9644012451172,
32.7469635009766,
-32.8983039855957,
34.7746658325195,
23.2320137023926,
-34.2790107727051,
-13.8471670150757,
-43.2205047607422,
-27.4638824462891,
30.9636211395264,
-24.7217960357666,
-13.4554023742676,
56.5530357360840,
-28.7691497802734,
-7.32895851135254,
81.7321166992188,
10.5616588592529,
-4.32384538650513,
12.2910165786743,
48.6169548034668,
27.7276668548584,
-48.0763854980469,
60.3589439392090,
40.0743522644043,
3.50808143615723,
33.2250404357910,
8.28403377532959,
-55.2463684082031,
-7.59323835372925,
37.3041000366211,
-52.5265960693359,
42.9570236206055,
-32.3755531311035,
-7.59858322143555,
40.1386489868164,
-11.8631219863892,
54.5292282104492,
-6.82842350006104,
21.0338592529297,
36.3951721191406,
22.4658908843994,
4.34960412979126,
46.2944908142090,
-7.30145454406738,
-23.1138057708740,
58.6632537841797,
-27.4358978271484,
31.5137290954590,
30.5505676269531,
5.89905023574829,
42.9229202270508,
0.124514818191528,
15.9243526458740,
-6.65290021896362,
3.84617185592651,
-6.03913021087647,
5.45538902282715,
62.3526840209961,
-0.359631538391113,
-5.67345142364502,
43.5125007629395,
37.9641990661621,
-51.1377754211426,
-22.6523132324219,
75.4267807006836,
3.03421783447266,
-33.1468505859375,
37.9790077209473,
57.2347755432129,
29.3526821136475,
25.6100349426270,
-0.0851778388023377,
16.8962650299072,
58.8201446533203,
41.4808235168457,
43.7223777770996,
29.3445167541504,
-2.54551839828491,
32.6331520080566,
73.3312988281250,
33.6107826232910,
16.1631984710693,
-5.76197004318237,
-11.4143676757813,
63.4592285156250,
-25.8799781799316,
7.09429359436035,
59.4276046752930,
-35.2657814025879,
56.3179092407227,
8.57839584350586,
-46.5519905090332,
-22.6838932037354,
-4.11652946472168,
4.95827007293701,
-40.3073616027832,
-0.137218952178955,
-14.0460643768311,
34.5145950317383,
-10.8393020629883,
2.92891120910645,
39.1809349060059,
-72.5137481689453,
20.8456401824951,
53.5971031188965,
42.6299934387207,
24.1206359863281,
32.3752441406250,
61.5419273376465,
-24.0136489868164,
-13.3359918594360,
40.4600677490234,
-8.98395919799805,
-55.1904029846191,
45.3682937622070,
40.9250030517578,
-46.6409912109375,
28.7134742736816,
55.3046760559082,
11.4072093963623,
17.9528789520264,
34.4405593872070,
21.5085639953613,
17.0573883056641,
35.0346641540527,
-9.69735050201416,
-6.81134557723999,
24.2908248901367,
-12.4102182388306,
3.84121298789978,
-23.2356243133545,
-50.0001487731934,
44.9265060424805,
-13.4945878982544,
-27.9967613220215,
98.8722991943359,
-18.6657791137695,
-35.0740776062012,
39.9780311584473,
-13.5365638732910,
54.4957771301270,
23.8523502349854,
-49.6923217773438,
51.7305603027344,
23.1026878356934,
-70.6432876586914,
26.0405502319336,
56.9123649597168,
11.3827857971191,
44.2048568725586,
56.0974731445313,
3.91970634460449,
-35.1637954711914,
-11.6864070892334,
7.77621078491211,
44.1591339111328,
23.2844905853272,
37.3971824645996,
20.6462249755859,
-32.4699020385742,
25.7892627716064,
46.7262535095215,
46.4656372070313,
-18.9133625030518,
4.89031600952148,
54.2401275634766,
49.3794860839844,
30.1828117370605,
26.2545547485352,
21.0995521545410,
-35.3406143188477,
38.7987442016602,
-37.3499908447266,
-39.7405319213867,
71.6416549682617,
3.75271034240723,
-24.4194927215576,
-18.6407051086426,
15.3702669143677,
-16.5108871459961,
-43.3701019287109,
-36.8318557739258,
-8.82016181945801,
-6.83035659790039,
-53.8244857788086,
37.8048934936523,
15.9248304367065,
1.17774105072021,
16.3749485015869,
-2.12938499450684,
29.6445960998535,
-30.4658660888672,
-12.9196491241455,
15.4451780319214,
8.47016620635986,
-3.90487384796143,
26.5473346710205,
14.4601325988770,
-59.7584381103516,
34.2714042663574,
41.0920677185059,
-48.6533279418945,
-11.7514324188232,
2.59301471710205,
-36.7827339172363,
29.8794574737549,
31.1121711730957,
-52.4577789306641,
0.0478725433349609,
7.42291736602783,
2.94688415527344,
35.8976135253906,
15.7741327285767,
15.8401660919189,
15.2078752517700,
52.2011032104492,
14.6087961196899,
-41.0808639526367,
55.5841636657715,
69.8906250000000,
-25.5742588043213,
29.4840106964111,
81.9374465942383,
6.09481430053711,
7.56262588500977,
0.320747613906860,
-13.2456045150757,
-21.6466903686523,
-13.8807983398438,
9.17115211486816,
1.73463249206543,
40.6215324401856,
27.1411361694336,
34.0321693420410,
-12.9487419128418,
9.83961200714111,
47.8771209716797,
-14.0075855255127,
27.3283843994141,
47.4807128906250,
-5.99007034301758,
-45.2923431396484,
63.5695381164551,
-7.02519607543945,
-26.6078910827637,
12.1947002410889,
-38.5225448608398,
59.2098808288574,
44.0908279418945,
39.7650032043457,
10.5468730926514,
39.9328689575195,
-12.8756523132324,
-37.3008995056152,
26.4428920745850,
0.346770763397217,
52.0539169311523,
-25.7810401916504,
18.9541740417480,
44.6357192993164,
-47.6646347045898,
52.0374450683594,
37.8737564086914,
-34.5322341918945,
29.8836669921875,
24.6195240020752,
-10.6123876571655,
-30.9111309051514,
16.2174110412598,
38.1928138732910,
-26.6872463226318,
3.87988090515137,
13.0289297103882,
-17.6387882232666,
-38.2688026428223,
15.4752578735352,
46.6862525939941,
6.92827081680298,
7.66363096237183,
-16.1815261840820,
-1.50519728660584,
-14.8467035293579,
-28.5128021240234,
4.50375747680664,
-21.9310188293457,
8.92942047119141,
55.9808959960938,
44.3950042724609,
-0.373243570327759,
14.5975723266602,
66.7208480834961,
36.7530441284180,
18.0065898895264,
-27.7742900848389,
-20.4165153503418,
42.1890983581543,
43.3672676086426,
33.5668563842773,
11.9822473526001,
-10.5786895751953,
-26.4719142913818,
30.3581771850586,
32.9885330200195,
25.2368335723877,
47.9783401489258,
-23.3023490905762,
-8.25023078918457,
-12.2309885025024,
-0.452745437622070,
28.2947692871094,
-20.8540096282959,
18.9683494567871,
54.6590118408203,
38.7357215881348,
-3.37261486053467,
29.7855529785156,
12.9371309280396,
-20.8663520812988,
46.4237480163574,
27.9431552886963,
22.3203639984131,
-6.61664295196533,
22.0090370178223,
53.7376441955566,
-1.09214305877686,
52.8759002685547,
49.2035865783691,
9.17134380340576,
-23.7362022399902,
-33.5315246582031,
-0.858318924903870,
-24.2008399963379,
-11.9808759689331,
37.8538780212402,
13.2673206329346,
-44.4420471191406,
9.00532817840576,
5.47119808197022,
-10.3362436294556,
41.7601280212402,
50.0566825866699,
48.3234443664551,
6.55210542678833,
22.3077774047852,
42.9455490112305,
43.7782402038574,
47.5892524719238,
28.5527114868164,
52.9655418395996,
45.4076690673828,
15.1088018417358,
-5.71790695190430,
-16.5104598999023,
-20.7904415130615,
-29.3073673248291,
-8.64891147613525,
50.0034599304199,
7.77114152908325,
-20.9253520965576,
53.0013999938965,
-41.0462074279785,
-23.4471855163574,
67.2901687622070,
-14.4616632461548,
-13.5745649337769,
10.3991193771362,
-22.4335956573486,
-7.73892307281494,
49.8694992065430,
-6.77420949935913,
15.7295141220093,
59.6716728210449,
-16.0650024414063,
-17.0186843872070,
-26.9283695220947,
39.3078002929688,
48.3781166076660,
18.2464904785156,
36.9710693359375,
19.1431579589844,
22.1116161346436,
21.1124019622803,
47.0105895996094,
-8.95982170104981,
45.1506385803223,
48.5069923400879,
-27.6616744995117,
4.99511909484863,
-34.4568481445313,
6.40036106109619,
50.8830680847168,
9.50724315643311,
-43.2404251098633,
33.6369209289551,
32.0658378601074,
-60.7992477416992,
49.4412040710449,
34.3105659484863,
-49.0690536499023,
-32.7522239685059,
-20.6513767242432,
32.7843475341797,
34.4085845947266,
-38.4963340759277,
-18.5019149780273,
39.2078056335449,
43.3165168762207,
48.4532012939453,
16.0043334960938,
30.4277839660645,
7.24683094024658,
-46.5008392333984,
57.5887565612793,
45.5357017517090,
-12.2367010116577,
40.8712997436523,
-18.6256752014160,
-33.6578826904297,
60.0662155151367,
21.1093826293945,
13.4929533004761,
52.2453536987305,
0.910593986511231,
39.8562164306641,
7.43019151687622,
-6.26946449279785,
71.5851593017578,
-13.7879257202148,
-1.86419296264648,
38.8975524902344,
-28.3630943298340,
22.1187763214111,
43.0952796936035,
21.9538803100586,
16.5812435150147,
22.3335170745850,
58.6732826232910,
44.9948272705078,
5.63706970214844,
-18.4682636260986,
17.0254325866699,
23.9197998046875,
-16.9564476013184,
-23.2596111297607,
37.7083969116211,
-21.9942150115967,
-41.2145957946777,
35.8810119628906,
-35.7111129760742,
6.27051925659180,
-11.0973234176636,
-4.03592872619629,
37.2295608520508,
-51.5926437377930,
-20.7070007324219,
-28.5569496154785,
25.6991844177246,
42.7606124877930,
-29.9114799499512,
5.29405546188355,
-17.5896263122559,
21.3617477416992,
58.7425003051758,
35.1736793518066,
21.0195732116699,
3.61074709892273,
52.9645462036133,
-41.1511611938477,
-7.31180095672607,
69.9738769531250,
-2.47900724411011,
32.2651443481445,
-10.3209352493286,
-17.0467491149902,
-7.28778553009033,
47.0917053222656,
16.6414184570313,
-9.42317676544190,
44.9300308227539,
-17.9113883972168,
-25.7622814178467,
-30.3288307189941,
29.7809047698975,
-25.2874698638916,
0.883092880249023,
5.69635009765625,
-11.8453531265259,
39.2825164794922,
1.95521891117096,
39.8819580078125,
-46.5532341003418,
27.6724643707275,
70.1546325683594,
-25.0499496459961,
-25.6607456207275,
14.2751073837280,
54.4296188354492,
-23.0607585906982,
-35.1759643554688,
48.8591804504395,
10.6640920639038,
-52.6361923217773,
-28.6822433471680,
16.9446830749512,
36.5236473083496,
-42.5523643493652,
22.8148651123047,
44.1301002502441,
8.85560798645020,
23.8204116821289,
14.3526382446289,
22.9640674591064,
-38.9376716613770,
14.0647783279419,
19.2649307250977,
-2.39382934570313,
54.8910713195801,
20.4398651123047,
-39.7779312133789,
15.5576057434082,
73.4987716674805,
3.04709148406982,
-14.3500299453735,
29.5810470581055,
9.46125602722168,
39.6233711242676,
55.2513885498047,
2.13784456253052,
50.7863388061523,
-7.79604530334473,
-1.84948062896729,
44.2237358093262,
1.39024496078491,
33.7402076721191,
27.7338771820068,
-3.60660266876221,
-31.0715026855469,
-18.0214424133301,
-23.3628902435303,
27.0671024322510,
36.6348304748535,
5.56622409820557,
-51.6577835083008,
33.0270195007324,
34.0569763183594,
-39.3451385498047,
67.3388595581055,
-35.1646423339844,
12.1906719207764,
-11.4140281677246,
-33.2732810974121,
7.38326072692871,
-5.24898433685303,
11.4810667037964,
-53.4065475463867,
74.5093536376953,
39.6022529602051,
-60.7120971679688,
-16.6032485961914,
22.6814460754395,
11.9906511306763,
16.4587135314941,
17.3938903808594,
41.5815620422363,
7.10988330841064,
-30.6848583221436,
29.9724464416504,
18.7793178558350,
31.3942756652832,
-33.7831916809082,
17.3890247344971,
60.9836425781250,
21.5350933074951,
59.7491416931152,
-11.2103290557861,
-4.96688652038574,
69.5499572753906,
28.4872570037842,
59.3192520141602,
54.5827789306641,
-42.1038208007813,
9.38249206542969,
-2.31496429443359,
-16.4424858093262,
-0.699090719223023,
6.07057189941406,
21.3466720581055,
-1.35911488533020,
34.0068817138672,
52.5469932556152,
14.8864164352417,
-36.0508728027344,
30.5912303924561,
30.6231746673584,
31.3927497863770,
52.5741653442383,
-23.9289512634277,
17.7857627868652,
47.2881393432617,
55.6087455749512,
23.0195732116699,
-20.1677207946777,
66.8027877807617,
60.5386199951172,
-11.6738967895508,
29.5320987701416,
61.5922393798828,
-4.37220764160156,
-49.8614311218262,
71.5158386230469,
30.6880512237549,
-28.4060974121094,
18.3770389556885,
-22.2214889526367,
33.2532806396484,
-20.5094909667969,
-8.97421073913574,
61.1138038635254,
37.6087532043457,
-19.6638107299805,
-1.44222927093506,
44.2649002075195,
-9.96711349487305,
-26.8720798492432,
-19.4512786865234,
23.5677757263184,
-40.7872810363770,
5.67736625671387,
25.1441192626953,
6.52752685546875,
57.5754241943359,
29.5512351989746,
16.2911529541016,
-34.5566101074219,
7.74720859527588,
-25.7899169921875,
14.6102123260498,
19.6842365264893,
-48.8445129394531,
-6.99011850357056,
-27.0994300842285,
35.5250396728516,
19.9524078369141,
12.5737056732178,
-27.1294555664063,
-16.7905235290527,
65.6848068237305,
-41.1453704833984,
-5.09780883789063,
27.2026004791260,
-26.5608634948730,
-37.3918724060059,
-6.91716384887695,
-4.72616672515869,
-8.58181667327881,
16.3102664947510,
-34.2378005981445,
3.40787410736084,
2.21193695068359,
17.4250793457031,
19.6622867584229,
22.0789527893066,
46.9082832336426,
-18.5772075653076,
28.9949283599854,
37.0215377807617,
43.3094558715820,
46.0635414123535,
52.8646392822266,
20.6577167510986,
-37.4704322814941,
35.3291320800781,
8.36418056488037,
12.2736148834229,
-8.04839420318604,
-42.4441833496094,
-21.9127979278564,
-20.3112773895264,
58.0590896606445,
44.2170677185059,
-7.74696922302246,
-29.1264877319336,
-7.91122531890869,
-10.6192245483398,
-8.74070739746094,
12.5017518997192,
-20.1308708190918,
19.0950736999512,
25.1141872406006,
6.45578193664551,
-2.04285502433777,
16.3190593719482,
11.8080263137817,
-35.4492607116699,
14.2957248687744,
45.6158447265625,
35.4498023986816,
42.2528724670410,
-19.8911228179932,
-21.6447448730469,
-2.80485320091248,
-35.5614624023438,
23.8902778625488,
40.9279365539551,
43.3715934753418,
4.88344001770020,
-24.9075355529785,
-12.2579059600830,
-14.9352188110352,
8.27290248870850,
-15.4158143997192,
11.6623859405518,
6.94879436492920,
-1.87506437301636,
-7.87166118621826,
-20.1248683929443,
26.7703495025635,
11.4826259613037,
-12.1715822219849,
19.8927021026611,
-2.05228424072266,
36.1997871398926,
50.4532203674316,
-19.0185775756836,
61.8047752380371,
16.8841266632080,
-28.9801406860352,
-10.1534118652344,
3.88559103012085,
32.8923721313477,
-82.2652969360352,
-5.74609375000000,
56.5557098388672,
-26.2245101928711,
-35.2787055969238,
-7.47698879241943,
25.3414611816406,
-19.6805763244629,
15.0610141754150,
20.5869789123535,
-40.1929473876953,
2.66282749176025,
45.2191734313965,
16.8326225280762,
-28.7516517639160,
-15.5831613540649,
-32.5155410766602,
-14.5229349136353,
29.2870712280273,
-5.67757987976074,
-24.8518199920654,
-46.7674026489258,
-12.2782230377197,
31.7296676635742,
2.73726034164429,
-43.2862510681152,
-41.4330024719238,
-11.1660337448120,
-24.2478160858154,
20.7945594787598,
51.1944465637207,
-10.0054740905762,
-54.6869888305664,
-24.8100204467773,
-13.5563735961914,
-3.38672780990601,
-2.74564194679260,
-38.0716361999512,
39.8855857849121,
5.98938655853272,
-15.7241086959839,
24.5921478271484,
20.7465953826904,
38.0263137817383,
-14.3332099914551,
59.3653602600098,
37.8994750976563,
9.68983078002930,
44.0563049316406,
-10.8180379867554,
45.3685684204102,
3.96232032775879,
-34.3638076782227,
-19.5415248870850,
-27.2513732910156,
-1.08095514774323,
-10.1190967559814,
6.54419803619385,
47.1771163940430,
47.9079666137695,
19.2796382904053,
18.9355278015137,
-28.9723472595215,
-9.11608314514160,
43.2791824340820,
57.6452064514160,
-2.49715018272400,
-19.4218578338623,
45.0007362365723,
-46.1957817077637,
23.4811687469482,
24.9165515899658,
-47.8225746154785,
0.347217082977295,
-25.5584354400635,
9.13996028900147,
8.21214103698731,
19.2149868011475,
35.3764076232910,
9.79279136657715,
11.7619409561157,
-25.2491416931152,
2.17401695251465,
32.6098327636719,
-20.1708011627197,
25.2812690734863,
64.7072753906250,
21.9721145629883,
7.00500059127808,
-0.640753149986267,
28.7318534851074,
5.49736976623535,
-35.2881011962891,
-24.2226734161377,
-8.25057411193848,
50.0491867065430,
25.5861396789551,
25.4138946533203,
17.7070713043213,
-4.17616939544678,
61.5384330749512,
-53.3057594299316,
-8.73436832427979,
45.4813652038574,
-17.5203361511230,
54.1852951049805,
-6.01364231109619,
30.6469116210938,
10.7276430130005,
5.33828067779541,
30.0968704223633,
-29.6912002563477,
23.0134544372559,
-22.1187992095947,
-14.4453010559082,
-25.1374969482422,
19.4841880798340,
54.9197387695313,
-19.5857238769531,
-25.7100715637207,
-2.57569885253906,
40.7874031066895,
36.8422508239746,
30.5629005432129,
-39.9057846069336,
-27.7225818634033,
12.2768535614014,
-1.51932168006897,
-17.4591865539551,
-3.15920829772949,
41.1683387756348,
-10.6026878356934,
12.7262077331543,
21.0476913452148,
7.28248310089111,
59.0833663940430,
44.0218276977539,
-0.449029922485352,
-26.3757400512695,
10.6511535644531,
44.6289596557617,
-3.92520785331726,
11.1799621582031,
58.8528823852539,
-17.5426254272461,
-7.40977811813355,
70.3262710571289,
18.2354335784912,
-2.05910491943359,
-17.1378765106201,
29.2627964019775,
56.4440460205078,
-38.5668258666992,
19.9740734100342,
23.9468822479248,
-59.2362976074219,
-27.0887508392334,
-16.2542991638184,
-2.13619613647461,
52.3249931335449,
6.50627708435059,
-27.0251789093018,
12.0657062530518,
-7.82910442352295,
-28.5089416503906,
-19.6015739440918,
69.6262054443359,
25.7392120361328,
-54.7776718139648,
29.2778778076172,
-23.7771186828613,
22.7600708007813,
65.1880950927734,
0.448881149291992,
44.4450340270996,
34.2637901306152,
41.7827148437500,
35.4584083557129,
49.3450050354004,
47.4178543090820,
-43.9443664550781,
-6.20310783386231,
61.5546188354492,
11.3644695281982,
-40.0890197753906,
-20.1746368408203,
9.69016075134277,
-10.8363685607910,
34.3854064941406,
7.56265592575073,
-24.3516921997070,
53.3171272277832,
-25.7228202819824,
-15.5333337783813,
49.8782501220703,
14.6187553405762,
-21.4622917175293,
-3.81568598747253,
14.0494318008423,
-25.1781368255615,
-17.5425529479980,
-27.8173923492432,
42.4067840576172,
39.7411422729492,
-39.2916870117188,
14.9244184494019,
25.7359275817871,
30.9219017028809,
12.2515125274658,
-33.5292282104492,
57.0403213500977,
42.8771171569824,
-31.7222499847412,
7.45107316970825,
18.0422019958496,
44.2829895019531,
-20.5685062408447,
-39.3495788574219,
57.9460144042969,
-13.4875335693359,
-28.7903842926025,
61.0807991027832,
42.1164665222168,
34.1645202636719,
43.6034011840820,
-4.44820785522461,
-11.4069833755493,
-8.80320072174072,
-6.19982194900513,
-7.48100471496582,
-41.0636291503906,
15.4373874664307,
3.60091471672058,
-3.00476169586182,
52.4556999206543,
27.7381610870361,
29.1092643737793,
15.4379367828369,
37.7184600830078,
-10.1546955108643,
-1.13768386840820,
100.786247253418,
-2.35666227340698,
26.3065910339355,
42.9185523986816,
5.55133867263794,
45.6904754638672,
-23.8720493316650,
36.1022109985352,
14.4997367858887,
-39.6554260253906,
29.5850353240967,
50.4558448791504,
-1.44919013977051,
-2.02964615821838,
46.5577545166016,
29.6794414520264,
30.1583824157715,
-20.5801887512207,
41.1888008117676,
36.8248100280762,
-36.3382301330566,
-21.6746978759766,
26.7180995941162,
40.0848579406738,
-69.8903808593750,
47.3750915527344,
41.2530975341797,
-46.5886611938477,
59.7901115417481,
23.2888202667236,
23.5623245239258,
29.8983268737793,
47.8283882141113,
10.7982540130615,
-35.7358207702637,
79.5066909790039,
-20.4460029602051,
-40.3320846557617,
79.6464233398438,
-16.1784534454346,
-58.1364669799805,
28.1226997375488,
35.1835784912109,
-45.6202316284180,
9.59875011444092,
41.3804550170898,
-51.2314872741699,
-11.8588829040527,
51.8420486450195,
5.61360073089600,
-26.6739101409912,
-9.14432334899902,
-35.6811180114746,
0.159370422363281,
49.7285690307617,
47.1629600524902,
29.1486873626709,
-15.3985729217529,
-16.6149291992188,
22.8531684875488,
5.45054531097412,
-13.7804450988770,
52.2025222778320,
17.5690517425537,
40.9561767578125,
20.3294067382813,
-32.1672363281250,
12.0551137924194,
-0.287441372871399,
-0.622557997703552,
-30.6339035034180,
31.6431121826172,
20.6001777648926,
1.31036186218262,
60.2748641967773,
33.5856018066406,
-0.373056411743164,
-2.89575791358948,
37.6555709838867,
1.83558666706085,
-36.2143898010254,
6.86289072036743,
-1.09400224685669,
-31.1304588317871,
-5.01857376098633,
10.7479209899902,
38.7504005432129,
42.3359031677246,
30.5252819061279,
-35.9746017456055,
-4.05776071548462,
43.2389526367188,
-25.1255912780762,
45.4949493408203,
17.2543640136719,
4.91984415054321,
45.8326950073242,
20.9991912841797,
5.79475593566895,
-6.64613580703735,
0.659970521926880,
-7.55199146270752,
-44.3136367797852,
-25.0690917968750,
52.5223083496094,
-48.7291297912598,
-46.1985130310059,
-3.89432954788208,
-27.9561500549316,
-16.1285324096680,
-38.5734443664551,
41.5016479492188,
-32.9540519714356,
-38.9241180419922,
52.8050117492676,
15.7722654342651,
35.8424949645996,
23.3189525604248,
7.65399742126465,
-10.7094659805298,
18.9461688995361,
27.1061592102051,
-25.8728103637695,
3.85351610183716,
24.3369102478027,
-5.48351955413818,
7.26063728332520,
58.9694290161133,
5.56164407730103,
32.5792541503906,
23.9903697967529,
-31.0809402465820,
32.5533599853516,
10.3538799285889,
8.92954444885254,
52.7483787536621,
50.6787567138672,
-41.5558471679688,
-17.9239826202393,
42.8503379821777,
-8.33806228637695,
16.6233348846436,
21.8516044616699,
36.3010597229004,
8.07016181945801,
-15.3485517501831,
9.26313495635986,
-32.5093917846680,
-28.7843532562256,
2.73996925354004,
14.5099048614502,
-14.9185256958008,
18.9735317230225,
49.8952293395996,
-32.2963027954102,
-31.5582733154297,
-4.99210596084595,
-5.09338903427124,
38.6778182983398,
53.1702003479004,
-22.4506607055664,
-47.4071426391602,
-18.4781799316406,
-32.6751861572266,
30.6081809997559,
40.9798927307129,
-22.1602172851563,
36.2546958923340,
43.3770828247070,
18.2816886901855,
-8.54724693298340,
4.57962036132813,
48.8210716247559,
-31.1158790588379,
30.7675552368164,
1.31817054748535,
-1.65750646591187,
40.7678413391113,
-34.4471206665039,
41.4576072692871,
21.8297653198242,
-3.41599369049072,
1.88023519515991,
47.3987197875977,
4.83428573608398,
-52.7366256713867,
7.81322050094605,
-23.7786235809326,
-29.3468990325928,
7.63041734695435,
28.8604621887207,
38.5203399658203,
38.1384963989258,
0.269594192504883,
3.25003194808960,
-27.5066299438477,
15.3132238388062,
16.1895351409912,
-38.0462722778320,
5.17651176452637,
-20.6492443084717,
52.6345100402832,
30.1215896606445,
-37.4171905517578,
28.4946861267090,
21.4388046264648,
-20.6813468933105,
-26.4814491271973,
35.2342300415039,
54.7414474487305,
28.0159683227539,
49.1387062072754,
10.7351322174072,
-31.9027309417725,
11.0891513824463,
33.3665657043457,
18.4189109802246,
34.8340301513672,
64.4683837890625,
19.2955780029297,
-12.1776742935181,
-10.4556236267090,
5.31603288650513,
38.9080009460449,
25.1219024658203,
-6.77331066131592,
-24.4858093261719,
17.6279029846191,
15.1184234619141,
32.6389274597168,
64.9512939453125,
44.5229949951172,
39.8498268127441,
-31.0617752075195,
26.2842941284180,
64.2897338867188,
-43.2022018432617,
11.4467353820801,
71.7356109619141,
-2.43882751464844,
1.12650680541992,
78.1011962890625,
15.7428741455078,
-31.0044288635254,
-31.6913661956787,
-15.2529125213623,
-0.730920791625977,
-35.9342498779297,
-2.43591547012329,
-43.3964347839356,
-7.31820774078369,
-19.5032863616943,
-32.1708374023438,
32.2432785034180,
-27.7484188079834,
-22.2425231933594,
-3.06395649909973,
27.1105403900147,
-26.7682495117188,
-11.0650663375855,
19.8159942626953,
-34.2246551513672,
34.1769104003906,
14.9006586074829,
-25.7157287597656,
20.1786746978760,
13.0495204925537,
-16.7747478485107,
2.16755676269531,
31.2085113525391,
16.7075843811035,
-2.73909091949463,
43.6564178466797,
47.1519126892090,
5.75925636291504,
-12.3663606643677,
33.9297218322754,
51.1378784179688,
-48.3302879333496,
-25.8335666656494,
18.9711761474609,
-3.04012846946716,
34.8467483520508,
-9.17883205413818,
-12.1039743423462,
53.0048599243164,
-38.0794677734375,
-30.2431621551514,
-6.57283449172974,
10.1413269042969,
11.4685173034668,
-40.3311767578125,
28.6859798431397,
-19.4134216308594,
20.1303672790527,
55.7013778686523,
24.5629749298096,
27.2214660644531,
25.0979995727539,
57.9187583923340,
54.7796859741211,
55.2344970703125,
-27.0209331512451,
27.4120121002197,
46.9070434570313,
23.9939880371094,
23.0638599395752,
10.6778821945190,
31.8035163879395,
-60.1684837341309,
-10.1066751480103,
48.2828674316406,
-4.24017906188965,
-9.56375789642334,
-32.3960456848145,
-35.5748863220215,
53.3529663085938,
-3.05525016784668,
-28.2908382415772,
7.13923168182373,
-33.8189201354981,
14.5289793014526,
17.8729286193848,
37.5747070312500,
-2.92313003540039,
-0.750293731689453,
32.4377746582031,
7.99421310424805,
64.4319152832031,
-20.7839221954346,
-9.92793846130371,
31.3204193115234,
-42.4845962524414,
13.8069667816162,
23.5590705871582,
20.5812301635742,
-18.8628616333008,
-9.15630722045898,
64.6982421875000,
23.3026161193848,
0.412445545196533,
-33.7208747863770,
-8.95684814453125,
41.3921279907227,
40.0683517456055,
41.4174995422363,
54.3546524047852,
35.5147056579590,
10.1525058746338,
11.0133981704712,
-15.8399066925049,
32.0766601562500,
8.41359233856201,
-14.7462949752808,
21.1515407562256,
-11.1009874343872,
41.1074600219727,
-17.6578254699707,
-44.2928771972656,
30.1251926422119,
0.658679008483887,
36.2244644165039,
42.4085998535156,
46.7440567016602,
43.3420295715332,
-7.85645294189453,
3.55951976776123,
8.10078620910645,
31.8075256347656,
-3.79620552062988,
-39.9584197998047,
8.81000328063965,
-11.4670381546021,
33.1152267456055,
29.6306228637695,
-39.9928665161133,
32.7747840881348,
43.6360664367676,
-34.4377632141113,
0.998863220214844,
66.4792633056641,
-9.13138484954834,
-11.8141174316406,
15.2025470733643,
-0.0914516448974609,
57.4435806274414,
26.2476615905762,
5.61931228637695,
59.4584541320801,
-37.5062103271484,
-34.3644332885742,
67.9742202758789,
-1.30667209625244,
18.9086151123047,
-12.0869874954224,
-40.9287185668945,
31.4429454803467,
25.1480083465576,
48.9941520690918,
2.31072092056274,
-39.6284484863281,
54.9687805175781,
37.8536643981934,
-35.8209533691406,
14.1812133789063,
24.8354377746582,
48.0586585998535,
6.04167318344116,
2.32018756866455,
67.4648208618164,
39.1609230041504,
23.4689388275147,
5.99351167678833,
59.3390197753906,
-3.71826362609863,
24.5799274444580,
71.3677291870117,
-39.4653778076172,
-5.45800542831421,
-1.76957952976227,
22.2765045166016,
20.6152667999268,
-18.8945617675781,
24.8339710235596,
19.5839977264404,
-32.4231262207031,
-5.22080230712891,
53.4477424621582,
41.4215812683106,
26.4283676147461,
61.7755355834961,
36.7583427429199,
5.46934127807617,
44.9978637695313,
-2.01243972778320,
52.8662338256836,
43.7402343750000,
-33.1737060546875,
28.9327487945557,
-19.8891868591309,
22.3899726867676,
6.88466167449951,
-42.8793754577637,
7.01857280731201,
-37.9132385253906,
22.0062122344971,
44.8081016540527,
25.1840515136719,
18.2618484497070,
-27.6425704956055,
-16.7756195068359,
38.0109863281250,
9.14877891540527,
32.2529602050781,
50.1184425354004,
-48.3586120605469,
-3.01258087158203,
63.9568824768066,
66.5667114257813,
-35.8619079589844,
-7.86157703399658,
-4.12297821044922,
-24.3732757568359,
18.1094970703125,
-18.9836769104004,
62.4713172912598,
-27.1936664581299,
-51.3383178710938,
-10.2921714782715,
-40.3260192871094,
-16.7371921539307,
-39.3836669921875,
-35.0007781982422,
12.6833534240723,
6.20063972473145,
-33.9188728332520,
56.3022575378418,
25.1983070373535,
6.05976963043213,
38.7816390991211,
-34.1905708312988,
35.7374877929688,
45.6376075744629,
2.76993989944458,
-1.33663630485535,
-15.7362842559814,
11.7832050323486,
-3.70856142044067,
-13.0646753311157,
5.09534740447998,
24.2485523223877,
-28.1183872222900,
-52.9589347839356,
19.4604969024658,
11.2560768127441,
-12.4970169067383,
24.8405780792236,
-5.00059890747070,
-45.3774147033691,
7.17235660552979,
20.8719215393066,
35.2525177001953,
15.0997724533081,
-35.3139762878418,
22.8745040893555,
25.6450271606445,
-8.70435619354248,
17.2879352569580,
-5.48067569732666,
-41.5630378723145,
-22.1705207824707,
30.9009666442871,
26.2020225524902,
-29.3691120147705,
-26.6593570709229,
-6.33823966979981,
31.9675254821777,
-7.40383529663086,
-13.6956453323364,
42.2417259216309,
14.5570745468140,
7.67316150665283,
-9.23764610290527,
40.6126365661621,
36.2150840759277,
-9.47357368469238,
-3.61359500885010,
-46.0390777587891,
-5.79778003692627,
-5.47630643844605,
-38.6568946838379,
5.68320369720459,
50.7071418762207,
-13.9602937698364,
-50.7789726257324,
52.2680244445801,
48.2508583068848,
19.8151321411133,
5.45232248306274,
-30.0628776550293,
6.16795539855957,
60.7785072326660,
44.0185127258301,
25.3754348754883,
48.1332168579102,
-35.0048675537109,
-43.6619720458984,
7.14210128784180,
22.4193325042725,
67.1094131469727,
-1.33734869956970,
18.6875476837158,
22.6411991119385,
-13.9909782409668,
14.8886156082153,
-6.24066781997681,
44.9967956542969,
18.3420734405518,
17.0341644287109,
12.6634798049927,
-27.3130779266357,
28.2734146118164,
39.4502754211426,
18.0874938964844,
54.8010787963867,
49.1259536743164,
-15.7799949645996,
49.6651458740234,
37.5935516357422,
2.37938213348389,
11.4980001449585,
-8.22846508026123,
0.665745854377747,
0.566502451896668,
-3.16152882575989,
-39.8245201110840,
53.5880699157715,
23.5173950195313,
-60.0067367553711,
68.5100173950195,
23.3026714324951,
-43.4158096313477,
11.9772796630859,
-0.743375658988953,
19.2831993103027,
28.8940849304199,
-42.9943199157715,
-1.13611316680908,
27.6716194152832,
-52.9810905456543,
32.0620765686035,
57.0599517822266,
-25.2183208465576,
28.6475620269775,
14.1133613586426,
-34.5542907714844,
-2.84926295280457,
33.6109466552734,
-8.26820468902588,
-42.7250823974609,
6.77104187011719,
35.8831024169922,
25.8651599884033,
0.334486603736877,
23.0694751739502,
-37.1076736450195,
-14.6100673675537,
21.1280860900879,
-44.2384643554688,
59.3658523559570,
51.1321868896484,
6.52562713623047,
-9.89633178710938,
-39.5492019653320,
14.7181301116943,
3.71101188659668,
29.3127498626709,
31.5729179382324,
-28.9541358947754,
7.64500427246094,
8.36117172241211,
-0.969327926635742,
47.5482788085938,
11.2177858352661,
34.2892723083496,
-1.92180824279785,
-20.8064022064209,
66.7097244262695,
-24.3987331390381,
21.2942543029785,
2.21844720840454,
-2.47888946533203,
69.2185974121094,
-13.5340003967285,
59.8294219970703,
-26.6133441925049,
14.5495700836182,
28.0606079101563,
-41.3996124267578,
39.5804481506348,
-32.8981246948242,
51.2290496826172,
-8.63072395324707,
-3.71852493286133,
77.9914093017578,
-14.8134384155273,
-16.5480136871338,
-35.5829849243164,
-0.798828125000000,
-22.3611011505127,
18.3010101318359,
3.34786057472229,
-32.3716812133789,
64.7399063110352,
-37.6601753234863,
-48.8005676269531,
22.6364002227783,
-29.4717369079590,
-26.7333660125732,
43.7050285339356,
-8.65721702575684,
-22.4559459686279,
42.4015274047852,
-18.9601821899414,
44.5999755859375,
44.9933090209961,
-27.0150051116943,
-2.41367483139038,
4.19890546798706,
-3.32833099365234,
-23.8571701049805,
25.0459518432617,
3.95838594436646,
-12.0297803878784,
15.3337316513062,
-39.2172622680664,
-36.5549697875977,
-21.1862754821777,
3.48155403137207,
41.7721290588379,
21.9729461669922,
31.5156936645508,
25.0370864868164,
-4.87986230850220,
-25.4235057830811,
-26.6808948516846,
23.2341861724854,
27.6520881652832,
-3.49718141555786,
-5.04595756530762,
-14.6685657501221,
-26.0547218322754,
17.1699218750000,
27.8605575561523,
-2.25507855415344,
33.6571846008301,
8.64057064056397,
-0.838920116424561,
51.1330108642578,
-21.9457244873047,
-49.5388946533203,
29.8365821838379,
7.85679340362549,
-62.0807685852051,
0.327605724334717,
6.92335891723633,
4.76768970489502,
38.6452445983887,
20.2756805419922,
56.6540184020996,
21.9059524536133,
-16.8490295410156,
-32.7629165649414,
11.8173484802246,
16.0417938232422,
-5.57627820968628,
16.7593383789063,
44.5939216613770,
40.0412559509277,
-48.8693771362305,
4.19495964050293,
55.0524063110352,
51.9052429199219,
-20.8848628997803,
23.3728466033936,
38.2310333251953,
-58.9601478576660,
21.4985942840576,
23.9777297973633,
19.5219535827637,
-14.0235118865967,
2.84460544586182,
-15.8584241867065,
-57.9114532470703,
51.2033081054688,
0.528772354125977,
-25.4131126403809,
34.6305885314941,
41.3762893676758,
15.0502223968506,
-44.3744125366211,
-6.43082332611084,
45.5148239135742,
7.53646659851074,
25.9957618713379,
22.8002166748047,
-15.1080360412598,
11.8819427490234,
-34.6823158264160,
18.0866184234619,
19.4521694183350,
-32.8783569335938,
61.2238960266113,
-6.35808563232422,
-23.4297943115234,
-2.71260261535645,
19.3933982849121,
17.4961776733398,
-55.2124633789063,
8.25322437286377,
-26.4409084320068,
-21.7167701721191,
28.0314807891846,
33.6584968566895,
-10.5634355545044,
-44.0702018737793,
63.2062988281250,
-14.5802726745605,
-43.7426948547363,
43.7838821411133,
25.6465148925781,
0.177347347140312,
-9.59468173980713,
80.6379470825195,
40.7430496215820,
-28.1801681518555,
53.0490760803223,
-5.71825027465820,
-53.9834747314453,
37.8621215820313,
16.9855804443359,
-14.7954158782959,
35.8552398681641,
-27.2395992279053,
-21.9386329650879,
-2.79233121871948,
-18.0965785980225,
40.0927162170410,
32.3668670654297,
0.535213470458984,
-64.1130752563477,
41.8748550415039,
36.4023971557617,
-39.8760948181152,
9.44950771331787,
-16.7720603942871,
34.8996315002441,
-31.2576522827148,
-26.2361335754395,
36.9370956420898,
-2.73215484619141,
-39.5737228393555,
14.3816909790039,
34.0920867919922,
-26.1197719573975,
20.4330062866211,
-3.53414106369019,
21.2322349548340,
9.09274673461914,
-13.5150938034058,
58.2236099243164,
9.44092845916748,
-22.3646583557129,
68.0720672607422,
7.24305868148804,
-31.7695217132568,
66.2879104614258,
28.6327209472656,
23.9140396118164,
-23.9951171875000,
-34.9660377502441,
20.8888301849365,
24.6705875396729,
54.6716651916504,
3.85786151885986,
-7.03864288330078,
16.4659843444824,
-41.4447822570801,
-9.97280979156494,
41.2379493713379,
35.1937561035156,
-13.2797584533691,
-42.6484909057617,
67.2419052124023,
8.54034233093262,
-41.4861221313477,
6.53725957870483,
26.0965862274170,
45.1129226684570,
3.76129436492920,
33.6488037109375,
2.39739227294922,
-16.7912979125977,
38.6159744262695,
17.8462028503418,
-51.6236686706543,
21.2054233551025,
-9.88814163208008,
-30.3106670379639,
45.2420768737793,
-51.7969474792481,
28.2986717224121,
51.8836021423340,
-22.5602684020996,
-3.92359733581543,
19.9767036437988,
-4.97031688690186,
-48.0368194580078,
-7.92227983474731,
24.9477500915527,
47.0437736511231,
-16.7282466888428,
27.8599433898926,
29.3696784973145,
-49.4721603393555,
60.3176879882813,
11.6370925903320,
-32.9140548706055,
44.5809478759766,
41.2066764831543,
21.1130142211914,
46.4227638244629,
51.7945785522461,
-27.1675682067871,
30.0972824096680,
38.8225746154785,
-38.5469512939453,
-0.884034156799316,
25.0362224578857,
29.6872425079346,
11.8452730178833,
32.3807220458984,
-5.26974201202393,
-40.4827308654785,
23.1104412078857,
-7.00459766387939,
-7.92383575439453,
7.29455614089966,
12.0484476089478,
34.5351409912109,
-29.4726047515869,
4.33217763900757,
33.1123237609863,
5.26559591293335,
54.5311012268066,
27.0700969696045,
-13.0599498748779,
-19.8847141265869,
-5.79470539093018,
5.14299201965332,
-32.3056831359863,
-32.3468017578125,
-39.9974479675293,
-37.7381362915039,
10.6410846710205,
22.6589298248291,
-16.6775493621826,
-38.1014328002930,
-7.97686195373535,
46.1596298217773,
6.26356220245361,
-30.0835952758789,
41.7991790771484,
12.3076105117798,
-8.51854991912842,
38.6011962890625,
51.1143569946289,
53.7658424377441,
43.6310920715332,
30.3538360595703,
47.3920326232910,
61.8667373657227,
-10.7305908203125,
-15.9275150299072,
-2.75095295906067,
35.1785583496094,
34.0593109130859,
-11.9060049057007,
43.5923919677734,
1.33374691009521,
28.4239044189453,
13.9785575866699,
-0.0238933563232422,
62.2430000305176,
-14.7754745483398,
17.3352298736572,
63.2537345886231,
-6.42363166809082,
-38.0557975769043,
-15.4122905731201,
-27.0998573303223,
-12.4860916137695,
1.91505336761475,
20.3749103546143,
35.8494071960449,
-34.3112411499023,
0.634907722473145,
35.9471549987793,
-43.7550888061523,
6.35307121276856,
61.2958602905273,
-7.90466499328613,
-30.4296321868897,
24.5383796691895,
64.5622711181641,
2.22318649291992,
-13.1712856292725,
-11.9267940521240,
-21.5467605590820,
14.3661766052246,
34.0864601135254,
-38.9934082031250,
-36.3362312316895,
50.9451103210449,
6.79313325881958,
45.1896743774414,
25.4981803894043,
26.7770786285400,
-11.6297073364258,
-16.6627235412598,
50.3036384582520,
-39.1168441772461,
55.6900711059570,
59.0085144042969,
20.9913482666016,
6.91581916809082,
4.04883193969727,
74.3276824951172,
0.179634094238281,
-4.72751998901367,
54.5309257507324,
-22.4253997802734,
-23.1865367889404,
57.6911239624023,
9.20060920715332,
34.3819046020508,
3.16913604736328,
-9.94673156738281,
22.8523578643799,
2.90671110153198,
8.43359184265137,
-0.150327980518341,
52.4894027709961,
28.2809333801270,
2.82201671600342,
4.96435260772705,
-13.0072879791260,
-29.2320537567139,
-25.9996566772461,
-9.99247360229492,
5.85128736495972,
-0.162868022918701,
-35.7240867614746,
-28.3420562744141,
-8.89979934692383,
-25.7451019287109,
-21.9895248413086,
-0.326226711273193,
-8.28740024566650,
25.0442771911621,
-25.7842864990234,
-23.3229045867920,
-4.85359859466553,
-14.6098384857178,
7.89038038253784,
-20.0551013946533,
57.7921295166016,
-1.59471511840820,
-33.9626808166504,
43.0436172485352,
26.9941215515137,
14.2254352569580,
-16.5262279510498,
-15.2462749481201,
-33.0930557250977,
-2.82779121398926,
0.308364391326904,
-23.9632701873779,
49.2787322998047,
31.4602718353272,
-22.7550582885742,
-26.4973430633545,
-23.9421806335449,
-39.9827423095703,
-17.1077308654785,
7.69212245941162,
-24.0742759704590,
-16.8554229736328,
-5.04059410095215,
42.1177139282227,
43.5849151611328,
19.8297557830811,
41.6583595275879,
6.95155048370361,
19.2745952606201,
15.0156431198120,
-14.6235446929932,
48.9282493591309,
17.3094635009766,
4.61989307403564,
57.1842041015625,
-18.4767265319824,
30.1261329650879,
59.6706428527832,
-30.4590148925781,
14.7063913345337,
-10.3094339370728,
-21.0060749053955,
60.8442306518555,
-0.667180061340332,
43.6076736450195,
49.0013809204102,
-54.9651260375977,
33.7784538269043,
31.5355682373047,
1.58555150032043,
18.9501819610596,
11.9785156250000,
25.1954250335693,
-28.3684387207031,
-4.06589126586914,
71.5260391235352,
-3.99810600280762,
-56.6991348266602,
48.4150009155273,
42.5398368835449,
38.4034309387207,
25.2743034362793,
-0.0770933628082275,
41.1010055541992,
-27.7986259460449,
-27.5390701293945,
-19.3225193023682,
-30.8261833190918,
-4.76402521133423,
1.47968447208405,
-31.2860889434814,
11.3660144805908,
66.4861221313477,
-20.1781768798828,
36.5118751525879,
36.3334655761719,
-50.5152587890625,
-27.4255199432373,
-7.53562879562378,
-1.30498933792114,
-28.2112998962402,
-8.86948680877686,
-24.8102436065674,
18.3174667358398,
19.6912040710449,
0.403644919395447,
38.5533142089844,
-34.3360443115234,
32.3923492431641,
-12.2254467010498,
-50.9921035766602,
58.2333450317383,
3.29916381835938,
-29.3872318267822,
14.0995941162109,
14.3367023468018,
-31.5371551513672,
37.4690895080566,
34.0752182006836,
-49.5364227294922,
15.9157752990723,
45.9905967712402,
-5.38473510742188,
-43.1219902038574,
-1.61158370971680,
34.9505958557129,
-7.91710996627808,
-28.3653926849365,
-19.6654453277588,
8.10469436645508,
-19.2335872650147,
-22.9072704315186,
35.8930244445801,
22.9210891723633,
26.7137680053711,
31.5147590637207,
34.3740272521973,
-3.08231163024902,
-4.47057914733887,
9.83677768707275,
34.5022926330566,
10.9740352630615,
-30.5283393859863,
65.1752700805664,
0.896215438842773,
25.2049179077148,
40.9555091857910,
14.4066419601440,
62.2508239746094,
40.0968093872070,
32.0045089721680,
12.6501102447510,
21.6598815917969,
-25.8819541931152,
16.4056205749512,
-8.27126407623291,
21.3080120086670,
73.5466232299805,
-46.0769615173340,
9.84208774566650,
81.7266159057617,
25.6353263854980,
25.4021282196045,
65.4001998901367,
9.59613609313965,
30.3858413696289,
16.1125106811523,
26.2011356353760,
45.6995086669922,
-44.9351959228516,
-16.6364746093750,
-4.40157127380371,
-22.0811996459961,
14.4857063293457,
8.89486408233643,
-36.7364921569824,
-21.9810295104980,
-39.6968536376953,
16.0207424163818,
22.7157936096191,
-72.1222457885742,
24.8355026245117,
27.7380237579346,
-14.0187253952026,
59.7746467590332,
36.3623924255371,
11.6450138092041,
38.4444580078125,
6.28993701934814,
31.0451164245605,
88.6238403320313,
-20.7064552307129,
-8.34207344055176,
80.1915054321289,
-26.0525054931641,
0.178851127624512,
70.3462905883789,
-22.1100006103516,
14.8754758834839,
72.1552886962891,
-34.1467247009277,
-25.8098716735840,
5.13767957687378,
-18.8394260406494,
-30.9423198699951,
-26.0015029907227,
58.1885032653809,
36.4481582641602,
1.59559249877930,
-20.1609497070313,
28.3799533843994,
77.5435638427734,
-22.0767822265625,
-0.493177890777588,
17.2449188232422,
-8.11318492889404,
-20.4080467224121,
14.9343576431274,
20.0498199462891,
-44.6715507507324,
49.4150505065918,
6.50408554077148,
-34.5529479980469,
59.8238296508789,
32.5589866638184,
-22.9408378601074,
-8.32549095153809,
54.1147689819336,
53.9411315917969,
42.9911613464356,
-36.1007690429688,
-5.78223323822022,
22.5230178833008,
-59.4553794860840,
7.44616222381592,
-22.0434188842773,
-7.40672874450684,
-10.9400205612183,
-12.2356796264648,
52.5556068420410,
-14.0026807785034,
44.0416336059570,
10.5074310302734,
4.50756072998047,
54.9901618957520,
-4.42509412765503,
34.4987525939941,
20.4278850555420,
5.82112646102905,
45.5283660888672,
43.7671432495117,
4.85733127593994,
-8.64855575561523,
22.1196308135986,
41.8805465698242,
0.256875991821289,
-21.4549522399902,
14.9463729858398,
18.9715251922607,
-19.1481742858887,
-30.8283805847168,
10.1806173324585,
-31.1105728149414,
-46.5234298706055,
5.20487976074219,
34.8874893188477,
-6.98146724700928,
-47.4624748229981,
37.6198348999023,
33.1973419189453,
43.2451972961426,
39.8700370788574,
-14.4219160079956,
36.7888679504395,
22.2588615417480,
5.02531528472900,
-22.9151515960693,
36.8068504333496,
49.3556976318359,
-63.5951538085938,
9.99448776245117,
37.9595832824707,
-52.7915306091309,
-19.1673717498779,
36.6130485534668,
-14.8406963348389,
-16.2755107879639,
-17.4392166137695,
14.6936101913452,
68.7749099731445,
-22.1911888122559,
-36.8728942871094,
-6.06769371032715,
-18.8617057800293,
24.5471687316895,
33.7490997314453,
-38.2356643676758,
-27.5450706481934,
-15.0961904525757,
-34.5649986267090,
18.6315937042236,
-44.3887786865234,
-6.37700462341309,
48.7554244995117,
-1.49680995941162,
-10.2805871963501,
-2.23109245300293,
56.0712356567383,
-14.3052473068237,
13.1731243133545,
16.1228637695313,
-37.7719612121582,
20.4837341308594,
28.9724769592285,
-6.27179574966431,
-4.09077358245850,
59.0098838806152,
-25.3234653472900,
21.9912681579590,
64.4624786376953,
8.08823013305664,
51.4430427551270,
9.05987930297852,
-21.9828987121582,
1.06083750724792,
25.8571567535400,
-22.4645195007324,
20.6508979797363,
24.2850074768066,
-51.3602905273438,
41.3640098571777,
32.2267379760742,
-21.6429901123047,
-29.2449398040772,
21.0008659362793,
58.0923309326172,
-34.6306457519531,
-10.2075786590576,
67.7960662841797,
27.5399055480957,
-23.3039836883545,
31.2440376281738,
5.91325378417969,
-43.1992835998535,
27.8478012084961,
42.7608413696289,
-14.8868570327759,
21.1647090911865,
30.8864269256592,
-50.2555160522461,
14.4865436553955,
69.4028015136719,
-30.2749176025391,
-8.35544776916504,
89.2088623046875,
-26.4966354370117,
-26.9458427429199,
-2.97540378570557,
12.4767732620239,
38.3122863769531,
-51.6120529174805,
27.6545963287354,
-5.77287006378174,
18.5454483032227,
32.3510437011719,
-40.3491592407227,
54.5842094421387,
14.0802717208862,
-49.1051292419434,
-3.67871856689453,
6.06482505798340,
-17.8535842895508,
16.8417663574219,
-19.7113037109375,
-44.5226783752441,
51.7721366882324,
31.2228736877441,
-22.7556362152100,
0.785496711730957,
-19.7772655487061,
-31.9841003417969,
15.8726434707642,
40.5803337097168,
0.159797668457031,
-40.8595314025879,
15.5346240997314,
58.4124908447266,
-32.7639083862305,
-37.2213630676270,
64.1694030761719,
16.7096900939941,
2.35391044616699,
31.4834594726563,
-29.4259586334229,
-27.1852149963379,
-30.2126827239990,
-27.6405029296875,
-9.49833106994629,
-10.3708209991455,
-6.74785852432251,
-34.4999923706055,
2.39714026451111,
19.2696208953857,
20.2808609008789,
-29.4704513549805,
-31.5523395538330,
26.3691425323486,
-38.1295051574707,
25.5553741455078,
22.4875831604004,
-24.3928680419922,
4.31093883514404,
35.0025062561035,
39.9990119934082,
-4.80580139160156,
3.88904762268066,
41.9153938293457,
54.0292358398438,
-30.9220504760742,
43.7976531982422,
7.43507957458496,
-40.6844253540039,
21.3998107910156,
-35.2009201049805,
-20.4527053833008,
8.03704738616943,
38.7940330505371,
16.8081245422363,
48.6607856750488,
45.0130844116211,
24.8302803039551,
-20.8864250183105,
-3.08376693725586,
57.8727722167969,
20.2554340362549,
42.3309555053711,
-19.9649105072022,
15.8774299621582,
12.4870624542236,
28.8776836395264,
69.5791778564453,
-26.8522491455078,
45.1597900390625,
20.6577796936035,
2.80493569374084,
39.3405227661133,
-16.8752708435059,
1.92919301986694,
23.6369552612305,
45.6072158813477,
12.2976627349854,
-30.5247039794922,
-29.3422565460205,
-13.1978454589844,
-5.33847618103027,
47.8667411804199,
29.8809909820557,
-33.2565917968750,
-6.43763875961304,
26.0972042083740,
29.5597381591797,
-27.5977821350098,
19.4791831970215,
45.6999435424805,
53.0396614074707,
3.13546037673950,
21.7941341400147,
39.6669654846191,
-18.9988842010498,
53.3426895141602,
39.9725265502930,
-18.2036857604980,
-2.19374275207520,
60.5415725708008,
-42.6027030944824,
21.8407726287842,
48.2529258728027,
-12.0590858459473,
68.3351898193359,
4.34612655639648,
47.7368850708008,
49.5274162292481,
1.82664632797241,
31.1887035369873,
59.6158447265625,
38.5002517700195,
23.4743385314941,
46.4972343444824,
6.56280994415283,
-18.9866180419922,
19.1649169921875,
42.8475761413574,
-20.9073314666748,
14.5479240417480,
62.4491500854492,
3.99833393096924,
22.6492137908936,
62.4042739868164,
39.9754028320313,
-18.3794555664063,
-1.66439414024353,
46.0792007446289,
-1.46182250976563,
-37.7341880798340,
5.03212642669678,
23.2432136535645,
14.3787117004395,
40.5541610717773,
-16.7261619567871,
-19.4686546325684,
56.5379486083984,
21.3099517822266,
25.6270160675049,
30.0540504455566,
38.7946243286133,
34.5697097778320,
-13.1211252212524,
40.4237442016602,
34.9885482788086,
-13.4589538574219,
7.38072872161865,
37.4094352722168,
-12.8649234771729,
-33.7993469238281,
-16.4623260498047,
28.1490402221680,
46.0510444641113,
-1.48755407333374,
30.0776348114014,
-16.0245304107666,
19.1662921905518,
26.3732547760010,
-27.4824180603027,
28.1433162689209,
14.8102102279663,
-29.8077869415283,
-18.4314937591553,
60.7257118225098,
-25.3389701843262,
-58.0172119140625,
24.5219764709473,
-31.1441879272461,
-47.2150077819824,
-22.1931266784668,
7.23556327819824,
-21.4043369293213,
-29.9720382690430,
14.7566175460815,
-33.8400344848633,
3.56798362731934,
35.7226448059082,
20.5974330902100,
34.9652404785156,
8.98002433776856,
60.1470413208008,
19.7035331726074,
22.0933551788330,
66.0807189941406,
-43.4571533203125,
-33.1440658569336,
7.87456560134888,
-38.5405197143555,
-6.87950134277344,
38.3066024780273,
-53.0765762329102,
-6.59260559082031,
47.0205459594727,
5.50269269943237,
46.2245178222656,
46.3077888488770,
47.7520675659180,
21.1806755065918,
38.1368865966797,
0.829345226287842,
30.1793365478516,
83.0699615478516,
6.64370918273926,
11.2797966003418,
30.5074996948242,
45.7086906433106,
-43.3888397216797,
-31.1652736663818,
38.8291854858398,
-4.12234210968018,
41.0018424987793,
9.36838340759277,
-17.1606960296631,
59.7790451049805,
14.5889320373535,
-36.4205284118652,
33.7046470642090,
18.8597583770752,
-23.6616706848145,
61.5059394836426,
37.0929336547852,
-3.48963832855225,
-4.58450984954834,
-29.6605358123779,
23.3449344635010,
-37.3350868225098,
2.93150711059570,
-0.718033313751221,
-45.3801803588867,
41.8931083679199,
-12.6542997360230,
-17.1515541076660,
-29.8571090698242,
13.6582813262939,
56.9396362304688,
24.0706195831299,
30.2419567108154,
13.1419410705566,
-5.91191482543945,
-24.7876701354980,
50.3031234741211,
33.7604675292969,
25.0299949645996,
20.4431114196777,
-24.0916538238525,
27.4667644500732,
35.6476669311523,
31.7236366271973,
0.475181698799133,
27.6288280487061,
3.96815109252930,
-27.6846427917480,
44.6560592651367,
-4.94415283203125,
-43.4786491394043,
-28.1029224395752,
17.8031845092773,
7.98565053939819,
-43.7336845397949,
13.9679527282715,
-1.40834927558899,
39.8486557006836,
1.78025436401367,
-19.0740680694580,
75.7213592529297,
-35.6895675659180,
12.6489753723145,
66.1700057983398,
43.6334648132324,
-0.591571331024170,
-13.7561798095703,
27.3397445678711,
-27.0247077941895,
63.1977195739746,
1.23897171020508,
-32.6420631408691,
18.9172554016113,
-21.0058021545410,
5.14123821258545,
-0.869509696960449,
42.5128326416016,
33.4116096496582,
23.8771476745605,
-7.21905994415283,
20.0266532897949,
55.5481605529785,
-45.1264305114746,
11.3535737991333,
37.4978713989258,
44.5022621154785,
32.0961837768555,
9.00239562988281,
3.29909729957581,
-37.4405975341797,
-1.69145679473877,
1.91075301170349,
11.1950836181641,
-24.0676631927490,
2.66724586486816,
6.91438913345337,
31.9159584045410,
13.5523538589478,
-38.8512573242188,
83.5553436279297,
-19.7234096527100,
-36.8776893615723,
2.99667525291443,
-14.1289949417114,
54.3732986450195,
-8.40070533752441,
43.1539688110352,
38.7260360717773,
-15.0791130065918,
21.1202297210693,
28.7666568756104,
-19.5367164611816,
-27.4315719604492,
54.0534248352051,
-29.8952198028564,
-45.2488403320313,
23.7269668579102,
-12.6579160690308,
-14.6479816436768,
43.9123611450195,
4.67913150787354,
-10.2180919647217,
24.1754703521729,
9.32237625122070,
28.0536975860596,
-37.7643814086914,
28.9461898803711,
3.33462715148926,
-63.2725334167481,
30.8656253814697,
-15.5169677734375,
-16.2186374664307,
3.83164739608765,
10.3284568786621,
-22.2437114715576,
-21.5756168365479,
48.5377349853516,
15.2602233886719,
13.6755676269531,
-26.7764244079590,
-0.631424903869629,
28.4709205627441,
-68.5978698730469,
46.6201477050781,
28.4214782714844,
-59.8323135375977,
-0.896148681640625,
27.6829032897949,
46.3527450561523,
-41.4791450500488,
24.9927883148193,
62.7160415649414,
19.2142868041992,
-1.14366471767426,
7.17471218109131,
6.66620254516602,
-37.1606864929199,
37.7882728576660,
28.2377815246582,
46.4154815673828,
-3.07686519622803,
24.9614524841309,
21.1528186798096,
-63.6990699768066,
52.5455589294434,
40.2922630310059,
-0.0766921043395996,
40.6302375793457,
8.56249046325684,
-31.9209785461426,
-12.1000709533691,
-39.2473030090332,
42.0551986694336,
11.6348571777344,
-1.13601493835449,
49.7886505126953,
-22.0859203338623,
48.5822677612305,
-35.6952667236328,
12.0400638580322,
48.0088806152344,
-56.6444435119629,
-16.1398029327393,
-33.4830474853516,
47.3417358398438,
-8.44478034973145,
-41.6270980834961,
64.3144607543945,
36.6001739501953,
-19.0960388183594,
-12.0617618560791,
39.6802520751953,
-9.28150463104248,
26.4631061553955,
5.43573188781738,
-23.9857425689697,
2.80302739143372,
-24.1054687500000,
3.87503051757813,
-43.4374732971191,
-1.74337005615234,
38.1417541503906,
8.50669670104981,
-8.65396690368652,
22.7832603454590,
48.9525680541992,
3.79080581665039,
14.9751148223877,
23.9783191680908,
29.2339897155762,
-11.6073560714722,
-35.4774894714356,
12.4923677444458,
19.8639659881592,
-12.5318069458008,
-27.8117198944092,
22.1869773864746,
60.4544448852539,
-18.7292747497559,
-44.8713073730469,
61.8434906005859,
32.7685546875000,
-2.09165143966675,
24.4674644470215,
-15.8086843490601,
35.6359939575195,
20.8219566345215,
30.3536319732666,
46.7960815429688,
-38.4501075744629,
20.8928527832031,
37.5564460754395,
-32.2318229675293,
6.05461311340332,
58.0691795349121,
8.42650794982910,
-8.16342258453369,
22.7145137786865,
45.8764991760254,
50.3272094726563,
3.83818006515503,
18.3752021789551,
57.2542114257813,
-11.7864370346069,
-25.8430347442627,
23.9326839447022,
3.91951894760132,
33.6768913269043,
41.7359352111816,
19.4040546417236,
-1.27754020690918,
-28.3850536346436,
54.5705184936523,
24.4412879943848,
-61.3413352966309,
47.9136390686035,
33.6135177612305,
-30.3816413879395,
40.6901550292969,
16.2736473083496,
1.04336881637573,
2.28790092468262,
-27.9613208770752,
-5.54315280914307,
-3.55136442184448,
-13.2769966125488,
-14.7121982574463,
54.6447525024414,
33.6851463317871,
22.8090152740479,
73.3297119140625,
-19.0260200500488,
-20.8968639373779,
-33.8088150024414,
12.4464473724365,
63.3785514831543,
29.0857028961182,
2.91205787658691,
3.82495236396790,
29.8762207031250,
-30.7990951538086,
8.13924217224121,
-32.6155471801758,
-2.91749382019043,
33.6561012268066,
31.9945278167725,
29.4528083801270,
-33.1490478515625,
78.2915954589844,
24.4325790405273,
-2.23599600791931,
-0.798614740371704,
14.3033676147461,
66.5330734252930,
4.35340309143066,
-11.9249744415283,
-10.9940662384033,
64.7090988159180,
-7.68869686126709,
-21.1178894042969,
64.4484710693359,
24.3812370300293,
-33.1133346557617,
-40.0614700317383,
61.0987548828125,
-1.73550605773926,
-27.3410377502441,
-11.8090209960938,
-26.0055332183838,
14.1627874374390,
-42.9024734497070,
-19.8474063873291,
7.94169807434082,
-3.95779323577881,
2.20361900329590,
35.8689804077148,
15.7628688812256,
26.0488300323486,
22.7040843963623,
-35.1516418457031,
43.4940185546875,
27.1615352630615,
2.89569664001465,
64.8184051513672,
58.5518722534180,
7.30100727081299,
48.5621376037598,
34.9426460266113,
5.09436178207398,
38.8918685913086,
-28.4072875976563,
19.0025367736816,
60.8331336975098,
-33.2279510498047,
-39.1837425231934,
22.4064502716064,
19.3374328613281,
-13.5095357894897,
-36.3707389831543,
31.5950717926025,
50.0982742309570,
-0.543982625007629,
4.85810708999634,
-6.82875442504883,
65.5322341918945,
38.2407569885254,
-34.3125991821289,
15.7002220153809,
8.37652873992920,
-9.19790458679199,
-6.02484273910523,
6.34166097640991,
24.0470600128174,
-30.6476058959961,
13.3589315414429,
54.1359367370606,
-24.8676834106445,
-6.26266288757324,
18.7290782928467,
14.1346397399902,
-5.02848434448242,
26.9490718841553,
13.7493362426758,
-20.1716060638428,
79.4497222900391,
31.7975807189941,
-36.6490097045898,
57.6570205688477,
14.4882774353027,
-34.9184532165527,
18.4298534393311,
-23.2815895080566,
41.7445831298828,
-4.25207424163818,
-28.6495113372803,
58.9517250061035,
-39.4371070861816,
59.2369461059570,
36.7904968261719,
-57.6777496337891,
34.9586944580078,
3.22627258300781,
-29.8302860260010,
11.5409889221191,
69.0866088867188,
-22.9061470031738,
-3.92972946166992,
65.6834030151367,
-25.3684272766113,
25.1604614257813,
53.5527267456055,
27.6998062133789,
-15.1395359039307,
-20.2824935913086,
20.1997146606445,
-17.1326045989990,
-14.0608425140381,
-15.3654499053955,
-15.1467189788818,
-36.2627639770508,
3.90755653381348,
31.5296249389648,
-36.9013557434082,
30.5541191101074,
29.0034542083740,
-20.2350749969482,
53.9851417541504,
49.3044357299805,
-20.9527854919434,
-34.2866287231445,
-14.9702119827271,
42.6422271728516,
-16.2320117950439,
-57.1235389709473,
34.2655029296875,
4.81431102752686,
32.8657760620117,
-20.5906181335449,
-9.66068267822266,
62.1867294311523,
-41.6988334655762,
-35.1509513854981,
-17.5509452819824,
6.41714668273926,
-34.1208229064941,
-13.2436866760254,
-4.88975191116333,
-10.0402908325195,
24.2947273254395,
-9.90520191192627,
11.2789096832275,
-28.1775112152100,
-23.9576263427734,
-21.0780830383301,
35.3355789184570,
27.3753623962402,
-19.8318195343018,
21.8179626464844,
5.02586841583252,
23.4601230621338,
42.0149383544922,
33.8601493835449,
47.8301086425781,
51.8771896362305,
14.9350805282593,
36.0720825195313,
24.5896797180176,
15.0830535888672,
8.78223991394043,
-20.5728778839111,
-37.6954231262207,
10.2356224060059,
12.6227788925171,
-46.7064895629883,
26.0623626708984,
16.6729907989502,
-37.5294418334961,
-35.6232223510742,
58.7444343566895,
-1.48314285278320,
-49.3667221069336,
76.6173477172852,
29.7502651214600,
-17.3410701751709,
2.24953746795654,
8.68315601348877,
-30.3103885650635,
6.73586368560791,
25.0534210205078,
4.20869398117065,
48.3612861633301,
14.6394929885864,
-25.9544353485107,
-0.702390313148499,
23.5590686798096,
-6.93141937255859,
-33.9405632019043,
-7.98737621307373,
19.6787185668945,
-35.5663795471191,
-29.7611732482910,
14.9765834808350,
-30.0466918945313,
19.2060356140137,
23.4415512084961,
-25.9117469787598,
49.7184982299805,
48.0229377746582,
-28.1753406524658,
43.6430053710938,
88.7471466064453,
-33.2496528625488,
-4.63796520233154,
44.1146011352539,
-0.322100281715393,
-12.8687734603882,
-36.6678085327148,
31.1716384887695,
47.3112564086914,
-25.5970458984375,
-18.7868652343750,
36.2944183349609,
27.2712230682373,
23.2276287078857,
-6.40736770629883,
-24.0839824676514,
52.5142822265625,
-22.6936378479004,
-23.4235191345215,
50.2154808044434,
-29.2494869232178,
-13.6838064193726,
13.3513011932373,
-5.41943407058716,
17.0641593933105,
28.0465736389160,
40.1270713806152,
41.2500305175781,
-5.09257411956787,
-30.9192562103272,
36.3119735717773,
49.5137100219727,
37.1953620910645,
12.5904970169067,
7.90744113922119,
29.0794372558594,
-49.6248703002930,
-17.8628444671631,
-38.5136260986328,
1.25684261322021,
16.6198883056641,
-57.0525588989258,
46.3168449401856,
-20.4939575195313,
11.3430290222168,
27.0210418701172,
13.5863723754883,
32.0108489990234,
7.39144468307495,
54.7799682617188,
-29.3369216918945,
79.2480697631836,
10.1585884094238,
-53.4464492797852,
71.4497222900391,
-18.2576351165772,
7.70988941192627,
-0.694607019424439,
13.4901857376099,
32.4633331298828,
-4.79518222808838,
0.564442992210388,
3.72170448303223,
16.9326229095459,
-29.5507602691650,
-23.0311031341553,
-0.141751289367676,
37.4188728332520,
-38.9766082763672,
3.68872261047363,
70.2226867675781,
20.6535644531250,
35.6596603393555,
-38.3660278320313,
59.1912231445313,
20.1501903533936,
-21.2364120483398,
32.5757904052734,
-3.25516533851624,
39.5726203918457,
-37.7486343383789,
-0.784150242805481,
80.3424453735352,
-14.8244552612305,
-37.7280349731445,
42.7741088867188,
23.2595863342285,
-18.8805942535400,
-4.74293994903564,
-3.38828516006470,
33.9017333984375,
4.78355073928833,
-55.6098747253418,
-3.80812120437622,
8.54364013671875,
-10.5936841964722,
-28.7580833435059,
-21.7420196533203,
2.71740818023682,
9.01144886016846,
50.4294815063477,
-0.0383849292993546,
25.7618713378906,
27.8614311218262,
8.52697753906250,
51.0288352966309,
52.0141716003418,
58.3871688842773,
-38.3129730224609,
52.3566436767578,
55.8261413574219,
-7.59521722793579,
95.0632324218750,
-6.83260488510132,
-10.5277853012085,
1.10100150108337,
3.38050770759583,
15.9826879501343,
-13.4487342834473,
52.3686180114746,
-34.1918792724609,
-35.0336418151856,
-17.7537422180176,
-20.0737571716309,
4.04958915710449,
-11.9960069656372,
72.3014755249023,
-20.3226242065430,
-32.1212081909180,
77.1426849365234,
12.9522247314453,
35.7537498474121,
34.6366958618164,
-34.0784683227539,
18.7030448913574,
7.21662044525147,
-12.8697595596313,
56.4763450622559,
2.61477661132813,
-16.4610824584961,
62.0949783325195,
24.4205284118652,
-22.8009223937988,
10.4292640686035,
27.4425621032715,
28.6955165863037,
18.6387577056885,
23.1284809112549,
82.1084594726563,
12.3682613372803,
-30.1043186187744,
14.8645896911621,
-30.3083686828613,
-40.3844680786133,
-13.6340770721436,
49.6167984008789,
-14.5614595413208,
-41.2307624816895,
60.2322578430176,
-29.2193412780762,
-9.72391700744629,
64.0006332397461,
10.4643993377686,
43.7939834594727,
5.54860687255859,
-16.4526710510254,
48.7560043334961,
11.9213790893555,
-16.5910568237305,
-39.5635185241699,
-5.68815898895264,
31.3606300354004,
-29.5566825866699,
16.6073875427246,
24.0247249603272,
14.2363271713257,
47.8487625122070,
-16.0815601348877,
-21.7162437438965,
-15.5395526885986,
-40.0612030029297,
-6.55402946472168,
65.2439041137695,
23.3580455780029,
-35.5275268554688,
-13.9547920227051,
3.24408054351807,
58.0079727172852,
-20.6285018920898,
-1.17774391174316,
36.6637229919434,
-78.8571395874023,
6.83209991455078,
43.9174079895020,
-24.8769531250000,
-5.45365667343140,
2.12126803398132,
-6.38163852691650,
9.58588600158691,
23.5592155456543,
34.4219017028809,
-5.30237770080566,
-47.8871116638184,
9.46323204040527,
1.08320963382721,
-2.82499170303345,
-8.00539684295654,
-24.7705631256104,
32.9736595153809,
-19.8117961883545,
-10.4124393463135,
63.3101882934570,
37.7603530883789,
17.7342815399170,
55.5160446166992,
-24.3822479248047,
-24.6054687500000,
72.7440185546875,
-21.5921707153320,
-16.4198646545410,
-2.62028980255127,
-7.68326854705811,
39.8943099975586,
41.1122474670410,
1.06094837188721,
31.9445648193359,
8.68129920959473,
-47.6272964477539,
21.1437911987305,
-16.7614212036133,
32.8094406127930,
6.81849861145020,
15.0017204284668,
37.9166526794434,
-38.9795646667481,
13.0274295806885,
3.49882411956787,
53.4152946472168,
-2.04123878479004,
-22.8297157287598,
-4.80698585510254,
-45.7038116455078,
23.3910217285156,
-24.2591323852539,
-45.3322677612305,
-43.2402572631836,
0.808758735656738,
37.1248245239258,
8.67886352539063,
8.53687667846680,
18.1573867797852,
48.9289817810059,
-21.5352859497070,
18.8076934814453,
7.83056735992432,
-11.2316083908081,
41.2554893493652,
-6.95046901702881,
37.7993965148926,
-11.9324951171875,
-23.1779460906982,
29.5973377227783,
-17.3583488464355,
30.2848587036133,
25.3037338256836,
-52.3994293212891,
42.9057083129883,
20.2734642028809,
-50.6235084533691,
9.48849678039551,
-1.52897000312805,
32.2226295471191,
-17.3571109771729,
-40.9622879028320,
37.6999740600586,
48.4209403991699,
-8.62780380249023,
-31.5473518371582,
47.4534530639648,
2.08774614334106,
2.31217980384827,
20.6766281127930,
-3.67144393920898,
58.7062683105469,
-15.3587760925293,
-18.5007743835449,
10.2412490844727,
-23.5109329223633,
-2.43067216873169,
-49.8119087219238,
-14.4431591033936,
11.4644260406494,
-45.4032669067383,
-3.81236457824707,
45.2573089599609,
-7.30420207977295,
-36.5975570678711,
3.17086887359619,
-1.50779056549072,
-3.68267107009888,
24.0191535949707,
40.5913696289063,
14.8096380233765,
-0.650712013244629,
51.8784255981445,
52.8342628479004,
11.8767690658569,
41.4161148071289,
19.4385375976563,
-11.1267347335815,
9.75733852386475,
-37.5469779968262,
15.0317945480347,
53.4031791687012,
-25.6837940216064,
-1.43679046630859,
37.0914001464844,
46.1326522827148,
-8.65701961517334,
-3.52723312377930,
71.5258789062500,
32.9899826049805,
31.2211322784424,
2.39491486549377,
40.8763999938965,
42.8098411560059,
-31.0391483306885,
38.6300621032715,
-27.5272274017334,
-24.3620948791504,
4.68598556518555,
-56.3471298217773,
-1.55636405944824,
-20.0605010986328,
16.9824905395508,
10.7235231399536,
4.57269859313965,
37.8109970092773,
-44.3538627624512,
27.5115947723389,
70.0784835815430,
-21.4401092529297,
-29.5775318145752,
29.8656578063965,
-8.72000312805176,
8.08457660675049,
19.4823265075684,
-41.1641273498535,
15.5410213470459,
21.0106391906738,
-20.9182281494141,
-27.4085998535156,
54.5503463745117,
23.1875076293945,
-22.7564353942871,
31.2619628906250,
-6.11584377288818,
4.80576562881470,
26.7619590759277,
14.4794778823853,
32.7131652832031,
21.4600429534912,
0.538476943969727,
55.4978561401367,
-5.67623329162598,
-46.3652496337891,
57.2048187255859,
31.3705425262451,
-29.2403049468994,
13.3548526763916,
44.1551589965820,
-51.6679039001465,
-24.8919982910156,
56.3308486938477,
-26.1998214721680,
-30.7090148925781,
35.2000389099121,
67.1904983520508,
4.80000782012939,
-22.7032871246338,
-15.0586223602295,
-8.87219047546387,
43.0400199890137,
45.0742950439453,
52.3723411560059,
-26.0563468933105,
-26.9050216674805,
21.8414669036865,
-2.75615215301514,
-24.0264453887939,
-12.5670585632324,
68.9546279907227,
24.3956794738770,
37.5874443054199,
65.1252899169922,
-24.6605205535889,
16.0153923034668,
66.0791397094727,
33.9801864624023,
25.6813983917236,
-7.30360889434814,
-24.3204441070557,
23.4301071166992,
-6.51382827758789,
-37.9111862182617,
18.0980491638184,
-35.0460243225098,
-48.7215728759766,
56.1608238220215,
-18.2273445129395,
-8.80942726135254,
22.9427509307861,
-54.7760772705078,
69.5376739501953,
46.2475776672363,
-6.84967517852783,
59.1026687622070,
-1.61383438110352,
-15.4367733001709,
31.4474258422852,
62.8282737731934,
-11.9632682800293,
-10.9853897094727,
84.0404510498047,
8.72799777984619,
-7.14603424072266,
66.6004638671875,
27.4316291809082,
-46.2227592468262,
8.68312072753906,
78.5696411132813,
12.4548597335815,
-21.0138206481934,
-29.0416221618652,
17.3656463623047,
24.1290168762207,
-18.7019233703613,
58.4699897766113,
27.8344326019287,
19.9645633697510,
63.4439392089844,
25.8087139129639,
39.8256072998047,
0.0157823562622070,
-34.2517814636231,
20.1514320373535,
0.462042808532715,
-39.5906448364258,
12.9986104965210,
40.3286972045898,
-37.2217330932617,
-37.4505538940430,
48.4557189941406,
35.3636779785156,
24.3101768493652,
28.7804508209229,
32.3503570556641,
49.6496582031250,
-10.2100677490234,
-12.0484533309937,
-3.89944481849670,
-22.9179649353027,
50.8893737792969,
33.5609207153320,
-4.58532619476318,
55.7219696044922,
-10.2099027633667,
-34.0340042114258,
41.8767051696777,
25.5204505920410,
22.0664672851563,
-5.33273029327393,
-23.0164260864258,
-2.84004497528076,
34.9662475585938,
51.0744857788086,
-25.9666137695313,
13.3513994216919,
68.5245819091797,
-14.4684152603149,
-7.25517463684082,
33.5875396728516,
-13.6319799423218,
9.07765865325928,
51.4102325439453,
17.3840751647949,
-12.0783367156982,
-7.08278036117554,
13.2710847854614,
18.2353134155273,
-11.1785173416138,
27.4185676574707,
2.06353473663330,
-30.6401882171631,
5.57884311676025,
-18.3354721069336,
38.6553077697754,
29.3714199066162,
32.9105186462402,
10.7667560577393,
25.9954071044922,
38.4454345703125,
-31.6955509185791,
57.3016128540039,
40.3890647888184,
20.9975585937500,
-21.6447067260742,
-7.83892774581909,
8.31022644042969,
-30.8576259613037,
41.0399208068848,
9.38831806182861,
2.59986424446106,
-0.142058730125427,
8.68827533721924,
51.0048332214356,
-9.22306060791016,
-42.9529495239258,
12.1791763305664,
-16.1223907470703,
19.0754528045654,
34.4653472900391,
-62.9796638488770,
31.2123908996582,
32.2616348266602,
20.8432979583740,
50.1777992248535,
27.2434349060059,
50.4722633361816,
31.0417232513428,
73.7833862304688,
-3.35263824462891,
-9.53439998626709,
36.6714973449707,
-4.69208478927612,
66.3171310424805,
48.1447830200195,
6.69694232940674,
7.15477848052979,
-2.80668735504150,
-18.1861495971680,
1.59790229797363,
-28.7023410797119,
19.4804039001465,
25.8522758483887,
-40.5472183227539,
47.0609550476074,
-9.10588836669922,
40.1726112365723,
34.5217437744141,
-52.8092193603516,
17.0175266265869,
6.54531192779541,
2.67896556854248,
-2.10395073890686,
4.03417491912842,
-29.5117759704590,
-36.1463088989258,
-3.94347286224365,
-12.4097108840942,
0.161307334899902,
7.57311868667603,
-22.6928901672363,
1.98987960815430,
54.8923416137695,
-31.0781211853027,
15.4965896606445,
32.5733833312988,
-27.8307189941406,
58.6750030517578,
-24.9874687194824,
6.36956596374512,
67.1866683959961,
-9.89021682739258,
1.06778812408447,
-38.2885055541992,
-3.16390132904053,
36.3112640380859,
2.78094315528870,
-1.63577413558960,
47.0433883666992,
-4.20477676391602,
-32.6640663146973,
64.0484771728516,
-21.0847358703613,
-7.25717830657959,
49.1462821960449,
-29.0060615539551,
-39.1810913085938,
4.17126846313477,
29.4776649475098,
12.1767129898071,
7.67562007904053,
-21.2352180480957,
-4.55727100372314,
-30.0471420288086,
-30.6201591491699,
14.3783903121948,
13.1917276382446,
34.9328994750977,
-15.8366832733154,
-25.9714527130127,
6.50407028198242,
24.4262886047363,
19.8144397735596,
24.1934871673584,
10.6549615859985,
-38.4237861633301,
-9.05747032165527,
9.92968177795410,
-2.04190897941589,
19.8094215393066,
-0.352606773376465,
-33.9245529174805,
-9.47094058990479,
19.2882614135742,
24.4596023559570,
-32.2062683105469,
-42.6084098815918,
-31.0905513763428,
-26.1351699829102,
29.2643318176270,
56.3785934448242,
34.9497947692871,
-20.7490177154541,
-32.8407020568848,
9.02107429504395,
7.63349390029907,
-22.6903800964355,
33.6264801025391,
-8.48313045501709,
-24.3185825347900,
30.5166625976563,
-47.4661026000977,
9.40251350402832,
58.6656951904297,
-21.6956481933594,
-24.7394199371338,
-23.7013759613037,
-5.04333639144898,
27.1350822448730,
-33.2651672363281,
3.10945439338684,
-23.2588272094727,
-38.9884376525879,
-12.1416988372803,
-38.9691276550293,
50.8962707519531,
-16.2949676513672,
4.72916412353516,
2.79224443435669,
-42.6812477111816,
17.4393787384033,
1.41136717796326,
21.5122032165527,
2.04826211929321,
-26.3331794738770,
-23.6249771118164,
35.9767150878906,
13.3746356964111,
23.0302181243897,
0.905185937881470,
16.1992416381836,
38.7650184631348,
-56.7681617736816,
6.91110229492188,
38.3956604003906,
32.4736862182617,
16.2205314636230,
52.0977478027344,
16.7387104034424,
-33.0211563110352,
-6.69313621520996,
-32.9649581909180,
51.8336791992188,
15.7946033477783,
-37.2993431091309,
65.3663864135742,
32.4405746459961,
19.1886405944824,
24.1217937469482,
-16.7270755767822,
33.5394592285156,
15.5334100723267,
24.8548202514648,
-0.999903917312622,
-14.6066112518311,
26.4185962677002,
-33.7210922241211,
-16.5596122741699,
29.9548873901367,
-31.5815811157227,
-44.6205940246582,
-0.929234623908997,
-56.5099601745606,
26.2893142700195,
19.8232383728027,
-12.3931541442871,
58.9685516357422,
3.44850897789001,
54.8341751098633,
7.73258209228516,
-23.9573745727539,
-8.54029655456543,
-38.3928070068359,
13.4027996063232,
-17.2285499572754,
-49.2518615722656,
-30.8537044525147,
16.2466506958008,
-0.331092596054077,
1.55881500244141,
43.6462936401367,
20.9043445587158,
-11.0698289871216,
5.87901782989502,
75.4067459106445,
-25.5606346130371,
-6.51836681365967,
56.5633277893066,
-13.3843698501587,
22.2958564758301,
34.9959564208984,
38.9382247924805,
-31.8146038055420,
16.9585914611816,
69.3002548217773,
-25.1475582122803,
-25.7564811706543,
11.4056930541992,
52.3293876647949,
13.5942878723145,
45.9477157592773,
25.1473178863525,
-42.9886970520020,
51.2465057373047,
29.9767837524414,
-25.9513378143311,
-1.39372420310974,
-5.65660095214844,
-27.3499908447266,
2.21463036537170,
-1.58894109725952,
8.23281669616699,
42.6285247802734,
-48.9688758850098,
-30.6295719146729,
52.4951705932617,
23.5647430419922,
-6.70821666717529,
43.3308181762695,
52.5447311401367,
-11.2347774505615,
-21.5528984069824,
33.3028030395508,
20.7605381011963,
-36.6008415222168,
26.3106365203857,
28.0931663513184,
4.16820430755615,
43.1037635803223,
-1.23480319976807,
-32.0760192871094,
53.6339683532715,
6.56592130661011,
-12.6987781524658,
31.9214286804199,
-23.4315261840820,
3.18547677993774,
-0.474252700805664,
48.9852943420410,
18.3651790618897,
20.4257450103760,
32.6044158935547,
-56.7258872985840,
-16.1281929016113,
-26.2554702758789,
21.7065677642822,
-7.12056207656860,
14.1129341125488,
24.9337539672852,
-17.7745361328125,
73.0923843383789,
-40.2398071289063,
9.99903011322022,
46.3796958923340,
-11.2608013153076,
30.8050365447998,
-38.1298332214356,
2.54891681671143,
0.353063583374023,
-16.5736923217773,
41.6545066833496,
52.6727104187012,
-21.6181449890137,
4.45816707611084,
61.0065803527832,
-33.0776214599609,
-0.955831050872803,
-0.892116546630859,
-16.5132217407227,
-7.63454341888428,
17.7646427154541,
20.7443466186523,
-41.8035697937012,
26.2193965911865,
-16.5919494628906,
18.5138702392578,
43.4830169677734,
-31.6445140838623,
38.7761383056641,
-18.8099822998047,
-29.2471733093262,
43.1466331481934,
36.5915336608887,
-26.6242828369141,
-35.0222549438477,
45.8722229003906,
25.6528148651123,
12.3968458175659,
32.6716423034668,
47.5241851806641,
35.0433158874512,
49.4473266601563,
26.3758735656738,
-44.0366935729981,
31.9455490112305,
-4.46246051788330,
-40.2468490600586,
32.8673515319824,
8.92981243133545,
27.9908790588379,
34.4323081970215,
13.0882282257080,
17.0415229797363,
42.4326248168945,
23.8197841644287,
-23.6958389282227,
-5.95948553085327,
-18.8821029663086,
17.0220870971680,
22.8401832580566,
33.2561874389648,
24.3908138275147,
-41.8711662292481,
25.4707336425781,
-10.8543872833252,
-5.99776458740234,
44.9429206848145,
18.2048110961914,
4.84799957275391,
-46.8932113647461,
-7.89624166488648,
-32.0791587829590,
-7.52326297760010,
-3.14662933349609,
-22.1670932769775,
34.5816955566406,
-39.5411682128906,
15.0458583831787,
-13.0295982360840,
-4.96499776840210,
43.4775238037109,
-40.0561103820801,
5.76665735244751,
-20.7705955505371,
-7.25214385986328,
19.9358291625977,
11.2274236679077,
-33.6806488037109,
1.65983581542969,
85.1706085205078,
-27.2365055084229,
-10.9211196899414,
-8.72388744354248,
-34.0302619934082,
8.97077274322510,
10.6083669662476,
46.3839263916016,
2.83468151092529,
3.95201969146729,
-5.20148515701294,
-34.6266441345215,
15.5436325073242,
13.4066705703735,
-2.14282631874084,
21.2347831726074,
63.0431785583496,
-47.4655380249023,
-45.0728569030762,
77.7515716552734,
-34.7816238403320,
-30.0584106445313,
25.0361919403076,
-23.2629642486572,
-11.8799486160278,
-36.3474006652832,
-20.9207820892334,
32.2398757934570,
-15.0922508239746,
-10.7171335220337,
8.16306495666504,
-53.2732086181641,
30.2245750427246,
43.4738960266113,
-30.0731639862061,
52.9520835876465,
46.0495529174805,
-39.9378089904785,
-22.6618785858154,
32.5930404663086,
44.2601318359375,
38.5936927795410,
43.1309013366699,
7.41731929779053,
-39.9427108764648,
7.39529561996460,
14.6684255599976,
-24.2034263610840,
2.72216939926147,
3.02227282524109,
16.8171386718750,
30.8648719787598,
-6.09352922439575,
11.1826038360596,
-9.76088523864746,
-33.2503204345703,
59.5855102539063,
-1.39949488639832,
12.2532510757446,
54.8431854248047,
17.2475872039795,
51.8791542053223,
-5.71126747131348,
24.1144199371338,
-18.0827522277832,
-0.674617767333984,
42.8474273681641,
16.6888465881348,
5.62807369232178,
1.09280967712402,
46.9888572692871,
-22.1561012268066,
62.9894332885742,
-8.06877136230469,
-68.1038284301758,
62.8045959472656,
-20.0149459838867,
-13.7426147460938,
15.2457389831543,
-10.2540388107300,
-14.5578355789185,
31.9201164245605,
44.4805984497070,
-39.6484527587891,
14.3122205734253,
26.5132751464844,
-19.2479038238525,
7.23744916915894,
-4.64350318908691,
4.67806243896484,
61.1128883361816,
13.6126308441162,
-48.4108581542969,
-19.4111328125000,
12.3563432693481,
26.1567859649658,
4.98017024993897,
16.4022827148438,
-19.8086929321289,
16.2948646545410,
30.9476203918457,
-49.5915451049805,
32.9430961608887,
32.4937744140625,
-62.3530883789063,
-24.3201408386230,
8.59930515289307,
-3.64540958404541,
25.5096359252930,
-31.8855361938477,
6.40352916717529,
15.8922300338745,
-7.32256603240967,
55.4613876342773,
-47.7863693237305,
3.07774925231934,
34.9603385925293,
-41.8342628479004,
14.8160724639893,
13.1062088012695,
27.8870887756348,
25.5297851562500,
-37.8265495300293,
-24.5556144714355,
-8.55745410919190,
55.0700798034668,
15.9785366058350,
-32.3495178222656,
62.9058151245117,
-28.1937847137451,
-58.9904212951660,
-13.0534000396729,
-13.2644710540771,
16.4344005584717,
-13.3929872512817,
12.8255205154419,
20.2131500244141,
20.8759746551514,
55.9507484436035,
33.0879859924316,
17.9791393280029,
17.3624973297119,
17.7796020507813,
60.5738601684570,
22.1960220336914,
-15.9093265533447,
-0.321088790893555,
6.49612426757813,
54.5982894897461,
4.44638156890869,
23.1997013092041,
20.8443050384522,
-26.3424835205078,
60.7885665893555,
5.95211553573608,
11.0863008499146,
55.7745819091797,
15.4433174133301,
25.0162525177002,
20.6801719665527,
59.9948425292969,
-22.7034702301025,
-36.2512321472168,
80.0903320312500,
6.48348426818848,
-29.7309837341309,
44.4759330749512,
38.5965232849121,
-14.7681446075439,
-20.1029701232910,
22.8434791564941,
41.0965309143066,
-22.6733036041260,
-23.2893409729004,
32.2728729248047,
40.4410324096680,
-17.3712844848633,
-43.0894165039063,
38.5686378479004,
-6.48858356475830,
-40.9961433410645,
32.4729537963867,
-2.82175588607788,
-18.7729110717773,
11.6565637588501,
47.4641189575195,
44.3442535400391,
-0.652723312377930,
59.2798004150391,
0.860581159591675,
-9.45928955078125,
86.4274749755859,
35.3104553222656,
-49.0846214294434,
28.2083702087402,
80.9842224121094,
-51.0420608520508,
9.85207176208496,
10.1488533020020,
-5.33730888366699,
12.0477743148804,
10.0202150344849,
58.9635772705078,
-33.9317092895508,
5.78172492980957,
45.4710388183594,
-12.1536903381348,
-35.6388664245606,
4.71610069274902,
-27.8216018676758,
-8.65551948547363,
11.9996538162231,
-25.0173454284668,
33.7927932739258,
-48.8307647705078,
-26.7593727111816,
30.1492691040039,
30.0692520141602,
49.1790733337402,
27.7192687988281,
-9.51859951019287,
-24.4518985748291,
8.02830791473389,
-50.3239898681641,
-4.92197418212891,
60.4758300781250,
5.66358375549316,
21.6808853149414,
-14.8417329788208,
-18.5407562255859,
20.1723709106445,
-52.8386917114258,
-11.2691631317139,
-22.4956130981445,
-24.4775276184082,
18.5007896423340,
-20.0890579223633,
40.0504837036133,
-9.32641029357910,
-36.3769378662109,
-21.1499118804932,
-14.0525083541870,
21.2413806915283,
-40.2720718383789,
10.7196741104126,
52.5559005737305,
-17.5891017913818,
-4.45426559448242,
61.3499755859375,
27.3517131805420,
11.3346138000488,
28.2396469116211,
-8.23670291900635,
47.3900413513184,
40.1054420471191,
0.782407760620117,
-33.1698074340820,
-2.30642700195313,
59.9802017211914,
-12.5403947830200,
-3.39042377471924,
1.04952263832092,
29.3553943634033,
4.10116577148438,
-25.7888584136963,
15.1503477096558,
-8.51755905151367,
47.5934448242188,
26.4334678649902,
-37.3375320434570,
16.0884418487549,
-28.9945335388184,
-49.2111396789551,
68.1294097900391,
13.0648918151855,
-17.8155517578125,
-31.3702774047852,
7.59931087493897,
46.7420768737793,
-34.2860755920410,
42.6929664611816,
4.00571441650391,
-15.6167135238647,
13.8131484985352,
21.0508079528809,
35.2661056518555,
-40.7351417541504,
-23.1630954742432,
-17.7313423156738,
23.8366107940674,
25.5677947998047,
-38.4797668457031,
34.1318817138672,
52.9761657714844,
-53.7788085937500,
10.9994964599609,
94.6759719848633,
-49.1702117919922,
11.9417629241943,
39.0886955261231,
10.3912086486816,
43.8921089172363,
-32.6321601867676,
74.0331802368164,
31.4176387786865,
-29.2732715606689,
34.7575950622559,
41.8788452148438,
19.5585746765137,
-48.4438018798828,
4.61224555969238,
10.0857725143433,
42.0089530944824,
41.0929794311523,
-22.9728622436523,
-7.49932909011841,
-20.2404098510742,
-18.1538238525391,
-34.7878723144531,
-19.8760833740234,
-2.03470420837402,
50.4850158691406,
5.31722354888916,
-46.2224349975586,
-4.83898687362671,
-29.0596542358398,
38.1354446411133,
-26.9662475585938,
-34.3480415344238,
5.57737064361572,
-47.3646354675293,
-17.0738735198975,
-36.6725730895996,
7.23604011535645,
20.7715110778809,
9.73480796813965,
-19.7787475585938,
-23.0810356140137,
-2.42437267303467,
-35.3662223815918,
36.9088821411133,
-8.94508075714111,
-24.2292461395264,
22.1781749725342,
-37.3923225402832,
-37.9951553344727,
-35.4846649169922,
-6.06553268432617,
-9.12400627136231,
-21.0152091979980,
21.6961898803711,
0.360321283340454,
-18.9627571105957,
49.7893066406250,
23.2224006652832,
-40.7831954956055,
34.1264343261719,
7.00019216537476,
9.90890693664551,
34.8778076171875,
-34.9190368652344,
-40.0508117675781,
-20.3511505126953,
19.6646652221680,
22.3242092132568,
32.5396728515625,
-11.0839157104492,
2.44611549377441,
52.6504402160645,
21.3964176177979,
48.0724754333496,
-5.57944107055664,
10.8585405349731,
17.7902088165283,
6.42867469787598,
36.4646110534668,
8.64035224914551,
-2.24790835380554,
21.5744380950928,
54.2587928771973,
-21.6131343841553,
36.9543418884277,
32.8428115844727,
-37.5083007812500,
35.7473220825195,
8.81546783447266,
-12.1175727844238,
20.6064186096191,
52.7703399658203,
38.0201644897461,
-30.2702980041504,
18.9990348815918,
68.0949401855469,
3.99767875671387,
-8.23177719116211,
-5.30648946762085,
4.46607351303101,
-27.5713024139404,
-23.9436798095703,
13.3295402526855,
-18.7290973663330,
-13.5669212341309,
-1.40467453002930,
36.7424736022949,
-3.53515338897705,
-23.5350208282471,
43.4942932128906,
44.0100860595703,
32.3402938842773,
-14.2655258178711,
-4.46758413314819,
-18.5890712738037,
-13.4795608520508,
44.3466567993164,
0.371843338012695,
-37.6443710327148,
-12.1911525726318,
54.6889610290527,
-30.8332023620605,
-5.97681856155396,
83.6619949340820,
16.7120342254639,
-3.79007434844971,
-11.8738756179810,
64.7554550170898,
-2.96436691284180,
-45.2375450134277,
24.3923301696777,
10.8171348571777,
44.0202140808106,
-18.7306594848633,
9.92471599578857,
59.2699508666992,
37.8503265380859,
26.1793594360352,
13.9845724105835,
37.5198936462402,
-14.0876197814941,
18.3346748352051,
-14.8793125152588,
-3.68856906890869,
71.1075134277344,
-5.40132331848145,
5.88000202178955,
26.1142406463623,
-0.147626876831055,
-45.3104515075684,
-10.7541103363037,
37.9080276489258,
-6.84341716766357,
11.5675544738770,
31.8760356903076,
27.1369247436523,
6.33631515502930,
-25.0445137023926,
11.5202140808105,
20.8649311065674,
21.5662307739258,
27.5282325744629,
53.0848388671875,
62.8984642028809,
7.33587551116943,
25.0771808624268,
-1.22939360141754,
-28.7197875976563,
-36.0710716247559,
11.5026493072510,
52.7456321716309,
37.4115219116211,
45.3318252563477,
12.8197488784790,
40.0326118469238,
-12.5042781829834,
24.6065769195557,
76.4538955688477,
22.2086868286133,
18.7449207305908,
44.2695541381836,
20.4513072967529,
-31.5280437469482,
20.5659217834473,
-17.4222526550293,
34.9670372009277,
60.4547767639160,
41.8566246032715,
5.56397151947022,
-16.8908443450928,
33.4060630798340,
-32.0376625061035,
1.66551303863525,
33.3835105895996,
30.3294639587402,
4.40254688262939,
32.7479171752930,
22.2681388854980,
3.55739951133728,
14.9580917358398,
-31.0233840942383,
-21.4950523376465,
-1.79137516021729,
27.2579097747803,
33.0121536254883,
-26.2543525695801,
-31.3156700134277,
59.5013542175293,
-30.8377952575684,
10.1532907485962,
36.7738571166992,
-24.8007774353027,
24.8556709289551,
-33.0052795410156,
41.5408058166504,
4.21459579467773,
-12.4156990051270,
33.4987564086914,
-33.5820350646973,
30.7822818756104,
18.1861057281494,
-22.1793708801270,
0.432362079620361,
53.4576072692871,
11.6089811325073,
-41.7989692687988,
23.1627006530762,
17.3374347686768,
5.31178855895996,
-16.7441272735596,
35.7685279846191,
55.3993301391602,
11.2145967483521,
7.44007205963135,
36.3906288146973,
49.4657402038574,
-61.8621215820313,
-9.61319065093994,
19.7344150543213,
-20.9587059020996,
11.7941293716431,
-27.4801826477051,
20.4278888702393,
5.58517456054688,
-32.4263114929199,
70.8652267456055,
-27.5605316162109,
-28.2683105468750,
64.7046356201172,
-29.3061676025391,
34.8334655761719,
12.7886428833008,
-50.2166023254395,
6.94099807739258,
-5.77162694931030,
-62.9687080383301,
3.82056808471680,
50.4528160095215,
-22.5722198486328,
41.2141647338867,
52.7498931884766,
8.92307090759277,
14.9979000091553,
22.3633098602295,
-5.53212881088257,
34.6293296813965,
7.98346948623657,
-26.0513954162598,
88.2857818603516,
28.5827007293701,
-39.7230415344238,
-8.56909370422363,
-13.9262275695801,
-36.1981506347656,
34.6711997985840,
19.6987648010254,
-3.12135076522827,
48.9044036865234,
23.6126518249512,
25.6593723297119,
35.3152389526367,
28.4858512878418,
0.332255363464355,
51.8980598449707,
-3.05152702331543,
13.9017372131348,
72.8367004394531,
-2.71321916580200,
48.2827606201172,
6.40679550170898,
-27.1249008178711,
-32.1922874450684,
-28.1058044433594,
46.3990173339844,
-7.68561983108521,
-4.53639030456543,
58.0706672668457,
35.0941772460938,
5.92058753967285,
33.8899116516113,
26.7560615539551,
-5.61817312240601,
-1.04145717620850,
-27.5961875915527,
36.3190345764160,
-4.14716529846191,
-34.4067993164063,
39.3266143798828,
-21.4610137939453,
22.8995494842529,
10.4021844863892,
-36.9674949645996,
-1.29831647872925,
11.5565309524536,
-21.8544673919678,
-39.0927925109863,
58.7663841247559,
41.3178329467773,
-37.7286491394043,
-27.4474887847900,
63.0528335571289,
26.7710380554199,
27.5518531799316,
38.2024421691895,
17.4481506347656,
53.9396133422852,
-44.1377944946289,
41.7370758056641,
3.63632106781006,
-0.174739837646484,
86.9932098388672,
-16.9605140686035,
-30.9137954711914,
13.3691959381104,
26.2047042846680,
-8.04517364501953,
53.1417121887207,
38.3862838745117,
42.0464477539063,
35.6449890136719,
35.8551979064941,
61.3031616210938,
-28.5982704162598,
-22.5855827331543,
-7.21011352539063,
-39.0016174316406,
-6.84123039245606,
33.4649314880371,
25.9555091857910,
42.8758125305176,
-15.5273284912109,
26.7561798095703,
21.6543064117432,
-50.9740295410156,
50.5789985656738,
3.50606060028076,
-23.9919700622559,
42.6880149841309,
1.45081448554993,
27.7322120666504,
39.2869949340820,
-22.0741615295410,
29.8476257324219,
54.5320396423340,
41.1576042175293,
9.14850521087647,
-5.38159465789795,
67.5987243652344,
-6.15302848815918,
-36.4119949340820,
46.7479782104492,
4.95962333679199,
10.3609762191772,
15.5438461303711,
0.906586706638336,
47.1500205993652,
-19.1869564056397,
8.76888275146484,
31.9170684814453,
-9.13612651824951,
43.1784095764160,
-28.2261810302734,
-34.5693168640137,
19.7907447814941,
-13.2619800567627,
8.90310287475586,
43.8602371215820,
-17.5119857788086,
-42.9825820922852,
-27.8208732604980,
-6.28683853149414,
35.3055343627930,
1.37956666946411,
0.481373310089111,
-28.8420333862305,
-17.1196746826172,
-22.1251831054688,
-23.2959747314453,
30.3575859069824,
21.9075431823730,
37.4585380554199,
-14.3327465057373,
29.6865348815918,
17.8624897003174,
14.5324974060059,
66.6283493041992,
-38.0093994140625,
29.6136436462402,
53.9490661621094,
48.2461814880371,
31.8140144348145,
-40.5531578063965,
27.1256790161133,
57.2448234558106,
42.3477210998535,
-29.5468730926514,
-8.89675426483154,
31.5461254119873,
18.6539268493652,
1.22024488449097,
20.0904426574707,
29.4150047302246,
-37.0464324951172,
12.8983736038208,
51.8026351928711,
38.7122726440430,
-41.6626091003418,
-37.2555847167969,
-12.3413438796997,
-8.40937042236328,
30.0695457458496,
-50.4751319885254,
-16.9762611389160,
49.0494842529297,
1.61075830459595,
11.4377651214600,
51.5929031372070,
11.2287673950195,
-36.4686851501465,
-27.9885959625244,
22.0247783660889,
-21.4884929656982,
-24.8103523254395,
65.7024002075195,
10.3332414627075,
-41.7522659301758,
3.30337524414063,
55.2884140014648,
47.4379234313965,
-34.7141723632813,
-14.1162843704224,
40.9884300231934,
-15.2337589263916,
42.3394470214844,
26.9243335723877,
-35.4791297912598,
46.8320655822754,
-7.67500400543213,
21.5980758666992,
71.7593078613281,
-11.5617675781250,
17.9486522674561,
34.8510932922363,
8.82158184051514,
29.0792541503906,
13.4840278625488,
-30.1401367187500,
-35.2942657470703,
-31.2525787353516,
-9.91954708099365,
24.2538490295410,
-8.88588047027588,
-33.9744033813477,
25.1937828063965,
16.3772277832031,
-58.2359771728516,
20.5689868927002,
28.6349754333496,
-57.0307159423828,
52.0347480773926,
57.0870437622070,
-1.05511176586151,
28.4116649627686,
-7.21761703491211,
-13.5303077697754,
-20.2596759796143,
37.9232902526856,
17.8474197387695,
-7.51672410964966,
42.8855819702148,
-25.6936874389648,
29.1144504547119,
52.1760482788086,
-31.3612575531006,
-0.640999794006348,
38.5052871704102,
3.12649559974670,
36.6478233337402,
23.7430305480957,
-6.22202968597412,
40.3560066223145,
40.6351280212402,
2.23291587829590,
-38.4849052429199,
32.7716064453125,
5.84490537643433,
21.1785526275635,
41.9938964843750,
17.8862037658691,
44.6153259277344,
-11.1723928451538,
26.0723304748535,
1.45995903015137,
-39.4084358215332,
-4.86564826965332,
5.18748569488525,
-0.665987014770508,
16.3965644836426,
22.4874114990234,
38.2205085754395,
16.7211914062500,
19.1360492706299,
29.4319667816162,
-8.29497432708740,
50.6016540527344,
-8.58471488952637,
-27.7168407440186,
-0.749685287475586,
-4.07681941986084,
-25.8764076232910,
-10.8883237838745,
-12.0517263412476,
-23.8388404846191,
34.9876213073731,
-46.8555603027344,
-15.1175889968872,
-21.1421699523926,
20.8622875213623,
45.4601669311523,
-41.5296058654785,
17.1882419586182,
-33.2052040100098,
-24.6130714416504,
11.8316192626953,
7.74099063873291,
-1.32550084590912,
20.8834533691406,
-15.6431350708008,
-69.9455184936523,
59.5694770812988,
-21.0459423065186,
-2.00111007690430,
30.2658443450928,
-55.6319274902344,
68.8587188720703,
26.8228492736816,
-23.2791957855225,
-0.573189496994019,
-7.56841087341309,
-40.8496170043945,
5.88975524902344,
59.1215820312500,
3.35235166549683,
35.9726295471191,
40.8119201660156,
46.4899482727051,
15.8115177154541,
5.80304336547852,
-2.24362421035767,
25.8084449768066,
61.5914154052734,
-24.7981834411621,
37.9758911132813,
46.9190483093262,
-27.5866260528564,
-11.6638631820679,
39.6805191040039,
30.9067459106445,
-59.9714813232422,
43.1020507812500,
8.10272216796875,
-54.5500564575195,
80.5558090209961,
-21.4265918731689,
-5.66187810897827,
26.5131034851074,
8.23485374450684,
14.3533201217651,
-40.0871124267578,
40.6672973632813,
45.4514427185059,
17.3095321655273,
2.54163694381714,
41.9930686950684,
-4.65491676330566,
8.86337280273438,
63.7071762084961,
4.68622636795044,
43.0961151123047,
-10.9960384368896,
-15.6344852447510,
17.9354515075684,
39.5769119262695,
7.03020095825195,
-14.9247932434082,
43.6546173095703,
-13.1965255737305,
-23.2387771606445,
28.9627113342285,
16.4635028839111,
17.7170982360840,
1.92635583877563,
-4.67136573791504,
56.7253952026367,
-18.5364227294922,
22.3615951538086,
21.4251785278320,
-41.1382598876953,
77.0917358398438,
30.4773254394531,
23.0159835815430,
34.9220352172852,
1.75295448303223,
14.6350688934326,
-30.4181137084961,
-6.19577026367188,
57.1214561462402,
-10.7620620727539,
-14.7162303924561,
96.0581970214844,
-9.47226715087891,
-38.7209930419922,
40.5778083801270,
7.48010063171387,
48.2316970825195,
55.2175865173340,
28.3824615478516,
-3.38139009475708,
5.56639623641968,
-7.42277860641480,
-19.8021087646484,
24.2666893005371,
-10.1628341674805,
-14.8463077545166,
28.9323387145996,
53.2259330749512,
-37.5849075317383,
-29.3100700378418,
35.2663497924805,
21.1926078796387,
18.3312816619873,
-12.3062639236450,
13.8360528945923,
18.9305458068848,
11.2045211791992,
-4.42275047302246,
-28.8545322418213,
-2.82901382446289,
26.0224685668945,
0.589850187301636,
-18.4838428497314,
2.77286958694458,
8.27189254760742,
36.7396545410156,
42.6966934204102,
17.9820842742920,
45.9787788391113,
52.8425369262695,
35.3648376464844,
-16.8655910491943,
-37.5510711669922,
18.7090015411377,
-45.5803909301758,
25.5785140991211,
39.8112716674805,
-36.1501617431641,
60.3058013916016,
28.0739421844482,
0.881470680236816,
-11.5452470779419,
4.85536766052246,
34.8697586059570,
-6.42173576354981,
-25.3719196319580,
-8.03083133697510,
15.8907489776611,
-5.95279598236084,
-3.41158699989319,
-18.5528583526611,
53.2065353393555,
2.20119285583496,
-72.5956649780273,
60.9063224792481,
-5.97662401199341,
-43.7767791748047,
2.05089473724365,
19.8220939636230,
31.3415775299072,
-29.5880451202393,
-0.0478954315185547,
47.6158905029297,
1.96764564514160,
-6.94285011291504,
41.1636009216309,
-41.1254730224609,
8.22567081451416,
3.31446027755737,
-12.9838151931763,
35.0462265014648,
-5.17055654525757,
16.5998172760010,
-37.7899551391602,
20.4294013977051,
-21.9280166625977,
10.9892759323120,
30.7019138336182,
10.8125925064087,
31.3445301055908,
-45.8910598754883,
72.0131454467773,
7.46688175201416,
37.6459159851074,
56.1192817687988,
-3.75091671943665,
42.9759063720703,
-29.9908638000488,
-9.62124156951904,
6.76123189926148,
45.2043838500977,
34.2513580322266,
-4.02843952178955,
-5.32818126678467,
-16.3102760314941,
27.8219757080078,
21.0524635314941,
-26.3804664611816,
-36.5616493225098,
-5.10495519638062,
-56.0225868225098,
26.0076026916504,
36.8338012695313,
-63.2737960815430,
-10.8765935897827,
-23.5784511566162,
48.1990890502930,
24.2924098968506,
-6.25292110443115,
39.2765121459961,
23.0209369659424,
16.4286746978760,
32.0641479492188,
42.9767761230469,
-44.8389739990234,
-12.2838153839111,
-0.767700195312500,
-21.6590118408203,
-25.3980007171631,
-36.8682060241699,
17.4737396240234,
26.0248336791992,
-7.76001358032227,
11.1157932281494,
64.5056076049805,
22.5289497375488,
-5.90171432495117,
57.1220741271973,
62.1064949035645,
43.2884750366211,
66.2892761230469,
8.87474822998047,
-7.69361352920532,
-12.0166225433350,
-20.8227348327637,
-44.9092063903809,
-21.0010852813721,
28.3013248443604,
-43.5159835815430,
11.7565793991089,
-10.7549400329590,
-55.5932540893555,
-5.32007741928101,
-3.16993975639343,
-8.90737724304199,
29.8457355499268,
33.6727104187012,
-39.8516769409180,
53.4028625488281,
57.9857215881348,
-11.9007549285889,
60.2652511596680,
3.59243202209473,
0.709884166717529,
90.4624633789063,
-16.2509555816650,
-18.0839881896973,
21.1089973449707,
-34.3188018798828,
21.8284721374512,
-11.0693616867065,
1.62202644348145,
56.1973609924316,
-7.73410034179688,
25.6745109558105,
52.2903404235840,
14.7692594528198,
27.1981067657471,
30.9938335418701,
-9.96166324615479,
16.1621856689453,
50.6097488403320,
24.1664009094238,
-27.2151832580566,
-8.27853012084961,
68.5686035156250,
-20.8045463562012,
-5.64966297149658,
12.7213487625122,
-12.5518035888672,
37.2802009582520,
-9.42415332794190,
29.5176029205322,
-18.0670833587647,
-42.0851135253906,
0.0673704147338867,
16.5014972686768,
67.3462295532227,
14.5155410766602,
1.96878278255463,
-8.93220520019531,
2.56643462181091,
-19.8740463256836,
-13.6512432098389,
46.5073165893555,
-17.2556858062744,
32.2470779418945,
14.8579206466675,
-26.7539424896240,
67.4816589355469,
21.7378120422363,
-25.5239219665527,
-30.6189823150635,
-14.1585159301758,
63.3915710449219,
19.3996372222900,
-22.4828853607178,
10.9887523651123,
-38.5718231201172,
-15.4265909194946,
42.7076759338379,
23.8355102539063,
27.6768226623535,
-17.5413360595703,
-7.90166378021240,
25.0776004791260,
-32.8725280761719,
28.6330871582031,
71.8200912475586,
-13.1021499633789,
-31.2866744995117,
-3.58579540252686,
23.1699905395508,
10.6247625350952,
-20.5655059814453,
-17.4170932769775,
-3.09876060485840,
23.1025829315186,
-13.3956623077393,
-41.1256294250488,
-4.80352210998535,
21.2031211853027,
20.0407676696777,
11.2884263992310,
57.8675041198731,
53.0563888549805,
31.1583328247070,
40.6668128967285,
49.0283851623535,
-14.1001911163330,
-46.6701507568359,
50.7153701782227,
-16.8815307617188,
-26.0019836425781,
28.1205654144287,
7.02199840545654,
34.2357788085938,
37.4148292541504,
34.6634902954102,
-38.5357475280762,
-24.8758602142334,
1.52127480506897,
1.31245648860931,
0.888443887233734,
-22.6408958435059,
43.3760604858398,
16.5555667877197,
64.0682983398438,
28.2895679473877,
-10.8835115432739,
47.1550445556641,
-38.4408187866211,
35.4711875915527,
21.6067810058594,
-2.90207171440125,
36.7571868896484,
0.697551727294922,
12.4197044372559,
9.73100948333740,
60.4442253112793,
-7.63756179809570,
-6.03657150268555,
73.8014144897461,
-24.6490001678467,
14.1331062316895,
55.9892349243164,
-52.9868354797363,
5.51988458633423,
1.87317371368408,
-43.5403099060059,
13.5751781463623,
51.8270301818848,
20.1314659118652,
-40.5917854309082,
39.0936965942383,
-10.4022531509399,
16.8012390136719,
38.4763793945313,
-5.74445629119873,
-13.9999198913574,
-29.9732971191406,
39.6045913696289,
-11.9117574691772,
24.9849853515625,
27.6326560974121,
17.7695407867432,
-12.3215045928955,
-21.2021102905273,
-14.8245944976807,
12.9387817382813,
38.8665542602539,
-46.0258140563965,
54.8475799560547,
10.0556287765503,
-0.291510581970215,
19.2800140380859,
-38.9751815795898,
50.5118827819824,
40.4709434509277,
-15.9408292770386,
54.5958404541016,
44.2061882019043,
-40.6939888000488,
0.0678362846374512,
-17.5059967041016,
-22.4976768493652,
18.6290779113770,
41.7604255676270,
14.3156776428223,
-21.9418640136719,
46.9641914367676,
36.2399864196777,
-19.1502647399902,
20.0873413085938,
-8.36535739898682,
-18.4397983551025,
45.3729629516602,
8.16050338745117,
-5.34109306335449,
-14.1448516845703,
-37.7544441223145,
18.6670417785645,
28.6896591186523,
-40.7680053710938,
7.31810379028320,
13.2421321868896,
16.6728057861328,
45.3625717163086,
-4.06401443481445,
66.8375625610352,
-22.7711410522461,
-7.72749233245850,
17.9517173767090,
-22.1815948486328,
76.6047439575195,
-14.6087427139282,
31.6965122222900,
50.0895080566406,
-31.1686935424805,
-16.3339004516602,
4.65268564224243,
-0.274983882904053,
-44.0411071777344,
6.32803916931152,
41.3960800170898,
34.0050964355469,
-35.1964607238770,
-20.0453033447266,
5.24298286437988,
-45.5377502441406,
44.2021751403809,
-16.7173290252686,
-36.3750381469727,
46.2626609802246,
-48.2087402343750,
-2.63302230834961,
25.7381668090820,
-51.0060348510742,
-8.22653388977051,
28.4816970825195,
15.3880577087402,
42.5335083007813,
51.2973136901856,
3.60102367401123,
31.9619235992432,
12.7410240173340,
-43.0352058410645,
38.9267272949219,
-5.95631980895996,
-21.7424716949463,
60.4042167663574,
-39.3277320861816,
-16.5611228942871,
20.2572612762451,
-40.8255157470703,
-12.1934795379639,
-35.8245697021484,
-38.8097763061523,
-15.7187948226929,
-41.1799392700195,
-40.5598907470703,
-8.76256752014160,
37.8206901550293,
22.6459808349609,
-30.1134338378906,
3.58909082412720,
34.4689559936523,
-5.03329467773438,
16.5978012084961,
45.1837539672852,
-36.8624076843262,
30.6398983001709,
53.3525810241699,
-32.4856109619141,
32.1353073120117,
-9.11712837219238,
22.4025878906250,
28.5358810424805,
8.38862514495850,
39.1883239746094,
-53.1570510864258,
49.5576171875000,
21.9561538696289,
-55.2944755554199,
21.9907531738281,
14.7234678268433,
39.7417144775391,
39.9957809448242,
23.6572151184082,
-37.5131340026856,
7.58909225463867,
31.4103050231934,
-1.64621281623840,
14.7090816497803,
-20.6752891540527,
54.3338699340820,
-19.4274482727051,
-49.2170829772949,
0.348520040512085,
-23.2768115997314,
14.8865537643433,
-2.67095804214478,
35.8851661682129,
7.14134168624878,
9.16254425048828,
55.1758308410645,
-34.7608795166016,
-34.2481079101563,
33.4303283691406,
2.97600412368774,
-43.3216361999512,
29.4680252075195,
37.2520751953125,
-8.58491420745850,
18.9536304473877,
43.9359283447266,
34.7904014587402,
9.86584568023682,
19.7205772399902,
13.4760379791260,
16.3661384582520,
-27.0922927856445,
21.9251403808594,
28.0873107910156,
-33.0576515197754,
79.8339691162109,
36.7848663330078,
-29.2418785095215,
-0.518084049224854,
14.1901130676270,
33.1941337585449,
4.79735279083252,
-0.366131275892258,
-13.5243492126465,
-2.17865848541260,
61.3099899291992,
-11.7773971557617,
-35.4855690002441,
43.6988487243652,
44.8357963562012,
44.7273330688477,
-9.40071678161621,
14.7472229003906,
18.0034027099609,
-16.8098392486572,
49.1282272338867,
4.31280803680420,
-14.9349937438965,
53.9214172363281,
-6.68159675598145,
-28.3039817810059,
46.3984184265137,
39.2457389831543,
19.7725219726563,
5.47690105438232,
33.6210594177246,
9.12194252014160,
30.3187026977539,
10.6483001708984,
-34.1370162963867,
66.4419784545898,
11.7056617736816,
34.7329254150391,
50.9957580566406,
29.3618888854980,
9.24076080322266,
10.0089664459229,
84.6657485961914,
38.0307006835938,
28.7734489440918,
54.2916641235352,
53.0180473327637,
-27.5826015472412,
-4.83180427551270,
64.4999313354492,
14.6229038238525,
-47.0129318237305,
18.3538246154785,
25.0487194061279,
-41.8160095214844,
32.0941581726074,
-1.95293235778809,
-1.05865573883057,
59.4923858642578,
-36.0639190673828,
-47.1359252929688,
35.4507026672363,
4.71611118316650,
8.93460845947266,
-6.31108856201172,
14.5409030914307,
21.2788600921631,
-50.6585693359375,
23.6876487731934,
49.2990493774414,
14.6999263763428,
-26.5479202270508,
38.5301971435547,
33.8972244262695,
-65.7235488891602,
15.7859420776367,
-13.6960277557373,
-14.7014255523682,
51.3843002319336,
-15.3257808685303,
-23.3882350921631,
11.6254186630249,
33.1655578613281,
13.0133914947510,
-32.7982826232910,
33.0302925109863,
57.8465728759766,
-33.4949150085449,
-25.7998962402344,
-13.7635898590088,
14.5334682464600,
23.0262165069580,
-23.9428997039795,
39.8152847290039,
47.3234748840332,
41.2220077514648,
28.9756088256836,
7.69866561889648,
-30.5041332244873,
-10.5019388198853,
37.4980125427246,
-42.7197914123535,
23.2562904357910,
58.8904838562012,
10.4284000396729,
-10.8369331359863,
14.9526519775391,
2.53072762489319,
-20.6316757202148,
44.5926170349121,
-24.2136688232422,
-18.1177463531494,
4.24718427658081,
-15.4494915008545,
-27.4367980957031,
-48.1147460937500,
10.7511148452759,
-30.4218215942383,
-19.8544158935547,
38.9985198974609,
35.3452148437500,
29.8341064453125,
-7.90698051452637,
-13.9051761627197,
59.0024108886719,
67.2525939941406,
-22.5932044982910,
35.3777542114258,
21.5914726257324,
-30.8573341369629,
52.8990173339844,
55.8799362182617,
30.1111297607422,
-34.0176620483398,
-12.9419736862183,
56.9495544433594,
-4.58641624450684,
-19.4633178710938,
-15.5077438354492,
-24.3863430023193,
15.0005168914795,
-32.0248184204102,
-14.8922977447510,
-3.77873516082764,
-43.7973899841309,
8.44419097900391,
-37.5078926086426,
-36.7367515563965,
13.1086540222168,
27.8368015289307,
6.70434951782227,
24.8522224426270,
53.4448318481445,
11.2026634216309,
52.1922035217285,
-4.31587982177734,
13.7205657958984,
68.5732116699219,
29.6881847381592,
14.3344783782959,
-4.62240028381348,
51.3112869262695,
3.73373746871948,
-4.08702230453491,
48.7295455932617,
14.5884618759155,
23.9595069885254,
43.1711120605469,
53.1071548461914,
-9.60271930694580,
-28.7621078491211,
14.8800449371338,
-1.01599979400635,
13.1571540832520,
41.7801742553711,
5.24210834503174,
-29.2988052368164,
44.0851821899414,
28.9754943847656,
16.7931060791016,
54.7285919189453,
-9.86303138732910,
9.12264919281006,
-0.449331134557724,
-22.0298099517822,
-22.3811740875244,
-29.6073608398438,
16.2735691070557,
-20.3754444122314,
-15.8558340072632,
-2.94251108169556,
-14.7634458541870,
42.5175895690918,
11.2852840423584,
-9.09924221038818,
36.0589790344238,
47.4743194580078,
51.9909515380859,
39.8550109863281,
35.4002838134766,
52.7566337585449,
42.1391868591309,
-1.78952121734619,
-0.479996681213379,
57.4693641662598,
-6.53283309936523,
-47.1481666564941,
43.3171272277832,
-16.3265247344971,
-22.3399391174316,
16.0217514038086,
-44.1331558227539,
38.3766174316406,
44.5495071411133,
-37.1050872802734,
-2.55176925659180,
50.1590766906738,
35.3036460876465,
-3.49131774902344,
2.74821233749390,
-15.2156562805176,
63.7256736755371,
23.4035453796387,
-34.6935386657715,
74.6509628295898,
-27.5945510864258,
-42.1530609130859,
-16.4544124603272,
6.83756446838379,
75.2046508789063,
21.4926376342773,
23.4938335418701,
0.856668472290039,
-16.9828529357910,
10.9061021804810,
21.6155204772949,
-10.5490608215332,
-17.6937828063965,
-33.6256866455078,
-11.3546504974365,
35.5329589843750,
8.48638725280762,
-25.8420104980469,
4.80203628540039,
19.1523666381836,
-48.9899673461914,
41.9486427307129,
3.07919979095459,
-31.9281558990479,
52.6400604248047,
23.5489234924316,
35.6864356994629,
-55.3985061645508,
20.4421501159668,
42.5756301879883,
-56.4667243957520,
48.1804847717285,
46.2313919067383,
36.6428070068359,
9.09752655029297,
0.326106905937195,
40.5945816040039,
36.4234962463379,
0.0111198425292969,
-1.68230438232422,
49.5040664672852,
-43.7360153198242,
-9.09674644470215,
53.9830551147461,
34.9420127868652,
29.7097167968750,
-32.1851387023926,
7.02096796035767,
14.6781730651855,
53.8702774047852,
23.9160308837891,
-9.59903717041016,
50.6890029907227,
1.46845817565918,
31.8269939422607,
-5.39031648635864,
-7.58959579467773,
27.7203559875488,
-42.0040130615234,
-26.1068801879883,
31.2733592987061,
-4.69852447509766,
-43.6078948974609,
11.3921117782593,
11.0085659027100,
-14.5183868408203,
7.43291711807251,
57.7199554443359,
-23.1594791412354,
-6.47144794464111,
83.6110534667969,
5.96532821655273,
-41.4744567871094,
6.42642784118652,
50.0273818969727,
5.40749406814575,
32.4126815795898,
18.1908664703369,
32.2621116638184,
17.0094680786133,
-39.3896179199219,
26.3318901062012,
-4.45182275772095,
-10.8877878189087,
47.2699661254883,
28.2329578399658,
-19.4648876190186,
41.0438308715820,
56.6928176879883,
-16.5756034851074,
20.9762306213379,
68.0652008056641,
7.69320487976074,
11.6360826492310,
71.7813949584961,
56.3117446899414,
1.17228698730469,
-31.6091117858887,
64.4939804077148,
36.4793930053711,
-29.0138702392578,
9.54978370666504,
38.6616668701172,
27.9679412841797,
-70.2928619384766,
6.31606483459473,
27.6047420501709,
-36.0140609741211,
37.9085006713867,
-2.66731357574463,
-2.98442077636719,
1.78100013732910,
-57.5635948181152,
28.8933830261230,
28.4639720916748,
-2.50964879989624,
37.8059158325195,
34.0542030334473,
-24.6547698974609,
-20.9164009094238,
43.0288772583008,
16.3478603363037,
-15.3682756423950,
-41.9530487060547,
3.15812397003174,
6.47350931167603,
55.9664077758789,
0.992494583129883,
-37.6707954406738,
61.6013908386231,
-43.4075698852539,
18.8277969360352,
13.3376712799072,
4.47624588012695,
28.7665405273438,
4.43887519836426,
33.8459091186523,
-8.38856124877930,
60.8762817382813,
-10.9571323394775,
15.9807310104370,
47.1819114685059,
-25.0100269317627,
24.7546577453613,
-8.93969058990479,
29.1047878265381,
37.8587150573731,
-25.1555061340332,
0.371402621269226,
-18.8192062377930,
-20.9729270935059,
45.9312438964844,
28.2926101684570,
-19.4390621185303,
-31.8327655792236,
-12.4833126068115,
-6.35660886764526,
-53.9835815429688,
5.53037261962891,
17.1547832489014,
-66.2564315795898,
6.01808547973633,
-22.8747062683105,
-26.2316741943359,
60.9183921813965,
-10.5995597839355,
26.9158611297607,
46.7054519653320,
21.1938266754150,
33.1959953308106,
45.6622695922852,
1.92314338684082,
-27.0486850738525,
70.3268737792969,
28.0705108642578,
5.09529495239258,
2.02548098564148,
15.3974370956421,
28.1547451019287,
-0.425858616828918,
25.1905555725098,
-53.9664192199707,
-8.73384475708008,
25.3670063018799,
-51.0100860595703,
43.1378440856934,
38.8371849060059,
-23.9229316711426,
22.3874740600586,
44.6049804687500,
67.1990585327148,
26.4235992431641,
36.6523094177246,
51.8584747314453,
2.14232254028320,
36.0691604614258,
54.7908973693848,
40.8771209716797,
20.1486339569092,
60.6381416320801,
1.39725875854492,
-31.0496006011963,
47.3302612304688,
-48.0097656250000,
-27.8022975921631,
-31.4790802001953,
-31.7160987854004,
50.2792282104492,
-4.52198982238770,
33.6288909912109,
-11.4104175567627,
-5.35083341598511,
26.5545253753662,
-12.4187946319580,
85.7480392456055,
30.4758987426758,
-28.6765193939209,
66.7038116455078,
36.9161682128906,
-9.00603199005127,
23.7053527832031,
52.8860702514648,
35.5114173889160,
-60.8297805786133,
28.5151157379150,
63.6374053955078,
-4.26360893249512,
50.7135696411133,
8.15285873413086,
46.6529045104981,
60.1807136535645,
-8.47289848327637,
-18.5217819213867,
39.3647956848145,
66.1486434936523,
-10.3706283569336,
11.4095096588135,
18.2990379333496,
-4.99716615676880,
12.4051952362061,
-9.73260402679443,
-17.0305347442627,
41.3637542724609,
-22.8011283874512,
-29.1510562896729,
59.8798332214356,
5.15189647674561,
41.4999122619629,
31.9038448333740,
14.7111682891846,
11.8600921630859,
-37.8325309753418,
55.3944511413574,
10.3854951858521,
-50.1284751892090,
-10.6518697738647,
37.2118225097656,
36.0450820922852,
-52.5849266052246,
7.56336784362793,
68.5651550292969,
12.0238304138184,
-35.6047515869141,
24.6652603149414,
17.0592498779297,
-32.0586585998535,
52.4350624084473,
23.2532958984375,
-28.5708007812500,
24.7710876464844,
14.4162025451660,
-35.4854927062988,
-6.97947502136231,
51.4366035461426,
-13.3552036285400,
-64.8850479125977,
55.7114906311035,
27.7098255157471,
-0.597212791442871,
49.7775878906250,
-13.0785236358643,
50.6796226501465,
41.0708007812500,
-28.9384269714355,
56.7672195434570,
17.0737590789795,
-4.20400619506836,
32.9507369995117,
-21.7712955474854,
48.6737785339356,
-14.8465671539307,
-6.54784965515137,
48.4890594482422,
5.96759033203125,
26.4197692871094,
-29.5712547302246,
56.5682716369629,
-17.2119655609131,
-35.2389183044434,
4.57485961914063,
-21.0196914672852,
82.1651153564453,
11.3456020355225,
26.9596805572510,
29.6371307373047,
-35.0845642089844,
37.8698883056641,
28.2047901153564,
-28.3778743743897,
40.4307785034180,
17.9702453613281,
-45.9481201171875,
-24.8458633422852,
-11.7289581298828,
50.9867706298828,
20.4152679443359,
37.6314010620117,
63.5244712829590,
-40.9893417358398,
8.33088970184326,
67.6667022705078,
18.9140853881836,
-17.8715972900391,
-26.7207641601563,
48.5855293273926,
10.9780483245850,
-40.2455177307129,
32.8253669738770,
15.3198595046997,
23.4199733734131,
-5.96048688888550,
0.413280010223389,
63.3381576538086,
-28.7010879516602,
2.14605045318604,
48.7850418090820,
-68.5436248779297,
2.93959045410156,
67.9517822265625,
-45.9034957885742,
-16.9961891174316,
28.6452846527100,
8.82680416107178,
-6.92403268814087,
-30.0772552490234,
-5.78355407714844,
41.1298255920410,
7.21906757354736,
-39.0216598510742,
28.4551563262939,
-1.07002258300781,
-37.6214675903320,
36.8928756713867,
53.9452819824219,
21.5088996887207,
5.83475399017334,
64.0420532226563,
47.2980346679688,
38.1724548339844,
26.3080692291260,
-0.665662825107575,
33.2527313232422,
-35.3620948791504,
38.4069366455078,
11.9542770385742,
-28.2142181396484,
65.4914169311523,
-8.36985492706299,
26.0829677581787,
16.4514198303223,
8.48368644714356,
27.1753730773926,
-36.6006927490234,
31.3604049682617,
37.5832023620606,
21.2737064361572,
18.2973289489746,
-20.1064186096191,
-13.3141727447510,
-32.2885131835938,
29.6901931762695,
3.51216983795166,
16.4477005004883,
42.8284988403320,
-47.9150772094727,
35.2850265502930,
2.87118005752563,
15.2788848876953,
56.2787475585938,
8.83810710906982,
11.9447841644287,
16.4728527069092,
34.3677291870117,
-6.21532821655273,
23.8929233551025,
12.5884504318237,
-29.7843570709229,
-35.2451629638672,
24.7278766632080,
-22.8689880371094,
-19.4494743347168,
30.7654933929443,
-50.5088386535645,
46.2794113159180,
-44.1361618041992,
-44.0505943298340,
-2.87606263160706,
-79.4076232910156,
47.9102973937988,
8.27644062042236,
25.7970046997070,
15.2257003784180,
-15.2300472259521,
54.8212585449219,
3.40679836273193,
23.1641311645508,
43.3865165710449,
26.9636573791504,
27.0641536712647,
34.2178306579590,
-9.06586074829102,
32.1867828369141,
16.0030517578125,
-38.9882125854492,
69.0935440063477,
28.4475955963135,
-39.1006698608398,
-2.74041271209717,
24.0478839874268,
-32.2166137695313,
14.9771032333374,
59.3880996704102,
16.7746715545654,
34.6060867309570,
21.9835281372070,
9.91108703613281,
1.71626019477844,
33.4819908142090,
1.69120073318481,
35.3789329528809,
24.6494865417480,
17.9327316284180,
39.7507095336914,
-75.7544631958008,
26.0738162994385,
3.19880294799805,
-20.3467674255371,
18.2531833648682,
-37.4229583740234,
55.2214660644531,
-11.6506357192993,
24.7912940979004,
35.1921806335449,
-36.4197921752930,
38.9263725280762,
-30.3459739685059,
-11.7874393463135,
61.9857673645020,
21.4927139282227,
-44.7115898132324,
9.57725048065186,
35.7687835693359,
-37.1583442687988,
-2.30020070075989,
-14.3738079071045,
-17.8733673095703,
-4.26652145385742,
-18.3720245361328,
-4.58024120330811,
16.1191883087158,
-4.61950254440308,
-11.9286708831787,
33.0250968933106,
-5.21286392211914,
29.1658229827881,
38.7035560607910,
22.8598632812500,
29.2557258605957,
-33.8407402038574,
-2.03013324737549,
5.76153039932251,
35.8062438964844,
-9.99355316162109,
-20.2094764709473,
72.0234222412109,
-33.4122467041016,
-36.7976379394531,
37.4557533264160,
72.5257492065430,
-0.868471145629883,
-40.7964820861816,
85.5695648193359,
47.2798385620117,
12.3782749176025,
13.0999984741211,
11.0021629333496,
-7.06439876556397,
-49.5701179504395,
-0.0143871307373047,
17.7801780700684,
5.75408363342285,
-12.0288171768188,
12.3481264114380,
-29.4339218139648,
-37.5956268310547,
50.8529090881348,
-33.2066001892090,
-34.1709899902344,
40.4844017028809,
-3.55742216110230,
8.21465778350830,
40.5062103271484,
-4.76463413238525,
-8.10848808288574,
21.2736835479736,
-27.7051258087158,
-12.3739271163940,
28.7178688049316,
27.0664768218994,
48.0073776245117,
38.2050285339356,
46.9083175659180,
51.1933975219727,
-10.7531185150146,
-20.6554908752441,
30.4734745025635,
7.38611221313477,
-25.5074920654297,
-7.69340324401856,
-0.226231664419174,
-15.8105545043945,
-37.7483444213867,
-8.91736793518066,
-0.911048889160156,
-28.6416721343994,
-43.6590232849121,
-33.4043540954590,
0.880043029785156,
19.7334613800049,
8.90373325347900,
-45.1463546752930,
18.6947212219238,
35.5349998474121,
-18.9124298095703,
47.0824546813965,
1.80967521667480,
-43.7010726928711,
-12.7916584014893,
-22.8553886413574,
41.3316688537598,
65.9966812133789,
-24.4963207244873,
7.04008579254150,
65.1271896362305,
32.1837768554688,
13.0017824172974,
-17.6856918334961,
-21.2054481506348,
-15.0291061401367,
-7.75977706909180,
-7.78646183013916,
-19.8032264709473,
26.1857395172119,
53.3113365173340,
-9.87041091918945,
-48.6296958923340,
-4.88750886917114,
5.61725425720215,
-27.0419559478760,
5.64520359039307,
-17.2624626159668,
-30.3902378082275,
13.1474742889404,
-45.7914924621582,
11.2894811630249,
47.6399040222168,
23.6642799377441,
10.1401214599609,
-37.7926940917969,
66.7881469726563,
44.9820556640625,
-24.1910648345947,
32.1840705871582,
-20.6957511901855,
-3.24776124954224,
74.1548767089844,
5.17471837997437,
63.8203773498535,
12.0557174682617,
-28.9477138519287,
66.6793975830078,
-37.0320663452148,
8.70466136932373,
-17.0943984985352,
-14.7080850601196,
48.5560035705566,
-41.3742828369141,
-0.583479881286621,
44.9773025512695,
-16.6173782348633,
-19.4029617309570,
69.4561080932617,
-18.3933563232422,
-15.9455795288086,
61.9383926391602,
-26.6654281616211,
16.7963676452637,
62.4471282958984,
18.5471858978272,
44.3956375122070,
26.5253982543945,
-10.9854087829590,
28.4894886016846,
41.2810134887695,
15.7569179534912,
-9.99474811553955,
26.2312355041504,
72.7807998657227,
2.52888226509094,
-10.2965631484985,
18.8133010864258,
18.2745437622070,
-10.8106994628906,
-29.5734786987305,
32.3613204956055,
12.8805704116821,
26.0657329559326,
35.4195060729981,
-26.6101760864258,
-42.1094703674316,
11.7295455932617,
23.0643634796143,
8.27188968658447,
60.2665977478027,
3.14730834960938,
-43.9917221069336,
51.5148010253906,
58.8868865966797,
-26.3393936157227,
42.3526649475098,
60.1498794555664,
23.1188869476318,
48.1068153381348,
14.7414131164551,
19.8776664733887,
34.8986282348633,
-16.0932388305664,
-29.9376583099365,
25.0237121582031,
48.5689544677734};
