byte in[8192] = {9,
0,
0,
0,
72,
179,
94,
64,
154,
72,
36,
192,
157,
226,
46,
192,
120,
163,
30,
64,
187,
127,
97,
64,
254,
129,
85,
191,
108,
241,
215,
63,
133,
146,
91,
64,
72,
74,
58,
192,
226,
50,
148,
191,
29,
50,
91,
63,
222,
216,
81,
64,
99,
235,
75,
64,
178,
148,
28,
64,
151,
40,
193,
63,
129,
229,
48,
64,
15,
196,
83,
62,
164,
74,
14,
191,
34,
221,
8,
64,
85,
251,
145,
192,
52,
48,
30,
64,
137,
38,
135,
191,
229,
241,
130,
192,
230,
186,
168,
191,
48,
73,
104,
192,
13,
142,
1,
63,
194,
168,
87,
192,
140,
51,
123,
191,
86,
81,
98,
63,
122,
34,
130,
191,
52,
231,
81,
63,
164,
1,
128,
192,
253,
74,
41,
64,
220,
39,
146,
64,
212,
156,
114,
192,
175,
223,
100,
64,
3,
84,
124,
64,
229,
40,
18,
64,
168,
181,
50,
63,
156,
226,
181,
191,
95,
149,
116,
63,
110,
235,
7,
64,
180,
101,
248,
63,
120,
117,
20,
192,
138,
173,
252,
191,
76,
223,
194,
191,
218,
93,
112,
192,
48,
133,
7,
192,
57,
214,
68,
192,
59,
202,
191,
191,
236,
110,
34,
192,
206,
46,
133,
63,
169,
191,
147,
63,
82,
55,
39,
192,
4,
118,
185,
191,
174,
108,
235,
191,
72,
255,
118,
192,
196,
17,
199,
191,
161,
197,
44,
64,
43,
227,
120,
192,
177,
125,
222,
62,
4,
231,
39,
64,
113,
224,
26,
63,
182,
92,
187,
63,
87,
59,
16,
64,
205,
253,
101,
64,
86,
221,
173,
63,
254,
149,
121,
191,
134,
50,
199,
191,
195,
1,
16,
192,
50,
125,
73,
191,
140,
153,
83,
64,
214,
255,
162,
190,
236,
111,
205,
191,
107,
231,
217,
191,
6,
149,
209,
63,
119,
219,
140,
192,
71,
208,
148,
63,
97,
48,
63,
192,
222,
168,
142,
192,
155,
238,
51,
192,
240,
134,
138,
192,
221,
169,
230,
191,
132,
254,
106,
192,
3,
130,
179,
191,
10,
105,
133,
63,
21,
149,
44,
192,
46,
54,
222,
63,
44,
122,
145,
191,
162,
196,
40,
64,
21,
100,
129,
64,
230,
175,
148,
191,
35,
193,
101,
190,
191,
242,
146,
191,
221,
26,
94,
64,
102,
93,
149,
64,
19,
128,
81,
192,
223,
104,
27,
192,
203,
90,
128,
64,
184,
221,
25,
61,
224,
203,
125,
63,
2,
24,
128,
64,
24,
142,
142,
62,
71,
82,
139,
191,
95,
228,
153,
64,
104,
102,
2,
192,
21,
133,
117,
64,
199,
210,
83,
192,
185,
139,
210,
63,
53,
224,
131,
190,
137,
195,
203,
191,
104,
110,
190,
191,
60,
56,
108,
192,
167,
126,
104,
192,
184,
146,
82,
192,
243,
141,
207,
190,
180,
114,
114,
192,
255,
183,
172,
62,
232,
59,
136,
192,
130,
16,
220,
191,
115,
204,
149,
64,
182,
47,
111,
192,
106,
81,
66,
192,
204,
143,
97,
64,
188,
51,
169,
191,
192,
178,
127,
63,
214,
197,
32,
62,
112,
211,
59,
63,
40,
0,
172,
62,
183,
12,
193,
63,
130,
158,
121,
191,
241,
177,
112,
64,
186,
146,
90,
64,
18,
88,
41,
192,
112,
214,
141,
64,
142,
7,
8,
192,
146,
6,
36,
192,
118,
95,
147,
191,
168,
196,
90,
191,
228,
159,
127,
63,
169,
184,
200,
191,
171,
50,
240,
63,
81,
255,
240,
191,
180,
29,
47,
190,
241,
134,
41,
64,
165,
171,
64,
64,
48,
165,
111,
63,
76,
19,
188,
191,
165,
139,
53,
191,
156,
202,
45,
192,
54,
132,
62,
192,
199,
43,
45,
64,
112,
201,
111,
192,
161,
45,
228,
191,
184,
12,
19,
192,
211,
157,
96,
63,
232,
234,
109,
192,
62,
44,
172,
63,
229,
118,
149,
191,
81,
192,
55,
192,
223,
88,
135,
64,
171,
190,
48,
192,
126,
238,
3,
192,
48,
11,
204,
191,
12,
218,
131,
64,
244,
209,
149,
192,
252,
38,
108,
64,
134,
118,
129,
64,
22,
192,
35,
192,
86,
97,
220,
63,
189,
86,
87,
190,
101,
80,
227,
63,
196,
75,
116,
61,
252,
187,
74,
192,
6,
7,
227,
63,
210,
31,
100,
64,
133,
110,
167,
191,
18,
51,
67,
64,
76,
136,
69,
192,
40,
117,
234,
62,
219,
170,
35,
192,
251,
176,
74,
192,
127,
168,
242,
63,
105,
181,
14,
192,
16,
4,
210,
191,
192,
40,
69,
192,
47,
140,
234,
191,
94,
75,
176,
63,
168,
197,
118,
64,
150,
186,
242,
191,
85,
130,
42,
192,
210,
217,
57,
64,
117,
153,
234,
60,
184,
21,
44,
64,
62,
51,
222,
191,
134,
224,
164,
192,
65,
250,
133,
64,
46,
214,
23,
192,
63,
192,
31,
192,
183,
249,
24,
64,
173,
52,
150,
63,
147,
54,
134,
192,
116,
130,
203,
63,
161,
105,
129,
64,
108,
104,
54,
63,
127,
35,
131,
64,
234,
204,
171,
191,
41,
230,
43,
64,
97,
130,
137,
64,
130,
244,
130,
192,
127,
123,
75,
64,
96,
252,
34,
189,
194,
156,
112,
192,
218,
95,
35,
64,
221,
62,
37,
192,
109,
169,
142,
191,
86,
38,
10,
64,
27,
226,
8,
190,
120,
114,
79,
192,
0,
145,
47,
192,
186,
203,
247,
62,
209,
103,
141,
64,
225,
197,
138,
192,
94,
123,
94,
191,
18,
79,
69,
64,
189,
57,
210,
189,
146,
141,
114,
64,
202,
129,
79,
191,
152,
116,
143,
190,
112,
228,
227,
63,
118,
176,
0,
64,
8,
63,
93,
192,
150,
163,
11,
64,
186,
171,
57,
192,
128,
95,
44,
192,
209,
118,
156,
191,
165,
182,
161,
192,
184,
151,
102,
64,
164,
164,
60,
192,
124,
168,
175,
192,
101,
235,
229,
190,
185,
38,
58,
64,
255,
38,
168,
192,
47,
20,
64,
64,
122,
240,
59,
64,
158,
26,
189,
191,
166,
66,
19,
191,
227,
157,
12,
61,
142,
89,
103,
191,
174,
92,
11,
64,
139,
237,
198,
61,
194,
122,
155,
63,
52,
159,
139,
64,
175,
121,
142,
192,
204,
210,
249,
63,
111,
160,
20,
191,
80,
2,
244,
60,
189,
85,
134,
192,
96,
187,
248,
191,
255,
240,
191,
63,
9,
85,
84,
192,
20,
51,
246,
63,
34,
88,
92,
192,
3,
5,
58,
191,
230,
221,
143,
64,
214,
98,
187,
63,
220,
236,
230,
63,
173,
154,
51,
64,
68,
182,
81,
64,
160,
23,
237,
190,
121,
129,
56,
64,
196,
246,
28,
64,
56,
112,
15,
192,
231,
60,
143,
64,
55,
131,
22,
64,
76,
52,
8,
64,
59,
97,
94,
64,
171,
75,
55,
192,
252,
172,
55,
64,
215,
224,
250,
63,
42,
141,
181,
191,
9,
65,
161,
64,
28,
37,
179,
192,
182,
136,
83,
191,
247,
78,
143,
64,
112,
222,
150,
192,
42,
171,
146,
191,
99,
66,
140,
64,
206,
37,
248,
63,
89,
125,
137,
192,
11,
24,
10,
64,
66,
106,
65,
62,
212,
246,
184,
191,
44,
150,
103,
63,
131,
214,
23,
64,
17,
63,
227,
191,
150,
241,
158,
191,
48,
77,
10,
64,
175,
74,
7,
64,
93,
209,
78,
192,
144,
2,
238,
191,
215,
252,
12,
64,
37,
176,
156,
192,
39,
192,
236,
63,
164,
42,
196,
62,
93,
145,
142,
192,
239,
199,
196,
63,
169,
188,
93,
192,
117,
92,
242,
191,
10,
122,
78,
62,
8,
38,
201,
63,
228,
34,
55,
64,
153,
146,
151,
192,
34,
20,
104,
64,
84,
214,
61,
192,
190,
122,
199,
191,
182,
65,
50,
64,
197,
56,
50,
192,
123,
68,
18,
192,
83,
158,
161,
63,
19,
230,
29,
192,
68,
187,
68,
191,
176,
217,
234,
63,
111,
32,
27,
64,
7,
84,
207,
191,
206,
33,
41,
64,
231,
15,
13,
191,
57,
105,
144,
192,
199,
194,
80,
64,
192,
75,
240,
191,
101,
158,
64,
64,
27,
140,
144,
191,
152,
18,
97,
192,
117,
0,
26,
64,
250,
109,
76,
191,
168,
41,
19,
191,
129,
239,
133,
64,
214,
69,
165,
190,
11,
123,
91,
192,
137,
105,
41,
63,
182,
6,
208,
63,
142,
142,
196,
63,
218,
222,
50,
64,
224,
123,
105,
192,
8,
95,
127,
64,
198,
17,
38,
64,
100,
151,
118,
192,
78,
192,
252,
63,
5,
165,
132,
62,
247,
119,
66,
191,
115,
68,
138,
63,
230,
233,
65,
62,
15,
101,
51,
64,
176,
192,
50,
64,
208,
4,
38,
192,
19,
21,
51,
192,
182,
170,
247,
62,
232,
223,
116,
64,
201,
92,
148,
63,
94,
52,
111,
192,
17,
190,
86,
191,
144,
83,
128,
63,
228,
246,
167,
191,
51,
72,
100,
192,
173,
70,
230,
63,
200,
232,
9,
64,
176,
105,
131,
191,
177,
104,
17,
64,
140,
166,
163,
190,
168,
124,
46,
191,
58,
170,
230,
191,
92,
153,
90,
192,
19,
144,
140,
64,
71,
27,
139,
192,
33,
80,
172,
63,
237,
94,
19,
64,
109,
83,
130,
192,
141,
146,
38,
64,
146,
216,
251,
191,
216,
69,
128,
192,
206,
24,
27,
64,
45,
210,
245,
63,
239,
25,
4,
192,
203,
38,
164,
63,
46,
148,
238,
189,
19,
190,
47,
64,
40,
89,
100,
64,
107,
221,
93,
192,
214,
219,
174,
190,
45,
128,
53,
64,
52,
118,
30,
63,
244,
100,
132,
191,
27,
131,
69,
191,
190,
199,
33,
64,
12,
224,
114,
192,
150,
214,
122,
192,
195,
158,
148,
64,
174,
225,
3,
192,
188,
79,
144,
192,
157,
113,
158,
191,
80,
198,
70,
191,
124,
232,
125,
191,
212,
144,
83,
64,
126,
236,
140,
63,
80,
216,
133,
192,
184,
212,
134,
191,
200,
222,
140,
191,
133,
224,
155,
191,
117,
173,
14,
192,
32,
207,
126,
64,
60,
91,
37,
64,
153,
190,
239,
191,
81,
187,
50,
190,
212,
158,
211,
191,
15,
150,
59,
64,
226,
179,
73,
64,
138,
176,
117,
61,
68,
228,
97,
192,
125,
235,
69,
192,
129,
249,
127,
64,
246,
134,
46,
192,
193,
193,
216,
191,
167,
121,
11,
64,
244,
248,
107,
191,
222,
234,
234,
191,
62,
182,
67,
64,
237,
145,
74,
192,
20,
86,
223,
190,
237,
41,
138,
189,
13,
237,
214,
63,
81,
150,
48,
64,
186,
125,
129,
63,
91,
228,
6,
192,
160,
120,
107,
192,
253,
85,
23,
192,
173,
250,
162,
63,
124,
249,
151,
191,
144,
146,
23,
64,
51,
15,
183,
63,
51,
71,
65,
63,
37,
54,
3,
64,
100,
185,
32,
189,
158,
162,
87,
191,
1,
61,
215,
191,
180,
204,
8,
62,
159,
137,
39,
192,
101,
216,
123,
64,
50,
116,
185,
191,
233,
240,
233,
63,
145,
159,
24,
64,
242,
112,
178,
63,
43,
249,
210,
191,
75,
210,
58,
64,
194,
83,
74,
192,
166,
216,
234,
63,
229,
169,
92,
63,
128,
228,
61,
192,
45,
131,
46,
191,
154,
35,
124,
63,
101,
232,
194,
63,
93,
36,
185,
191,
4,
220,
119,
191,
133,
217,
119,
192,
20,
59,
186,
63,
234,
255,
87,
64,
61,
206,
143,
191,
48,
240,
0,
64,
178,
120,
66,
191,
117,
250,
55,
192,
150,
132,
134,
64,
14,
219,
206,
61,
23,
1,
179,
191,
101,
170,
93,
64,
178,
1,
13,
192,
82,
80,
164,
63,
30,
243,
85,
192,
57,
102,
72,
63,
105,
88,
235,
191,
249,
40,
168,
191,
181,
109,
158,
63,
56,
74,
67,
192,
122,
211,
130,
191,
72,
180,
185,
61,
6,
69,
20,
64,
73,
14,
80,
62,
230,
233,
96,
64,
67,
154,
101,
192,
21,
146,
222,
191,
246,
194,
118,
64,
114,
134,
155,
63,
101,
34,
79,
64,
64,
164,
149,
192,
84,
159,
31,
192,
14,
191,
24,
64,
158,
125,
148,
192,
6,
241,
151,
64,
24,
78,
25,
192,
84,
24,
19,
191,
59,
155,
212,
63,
228,
103,
82,
63,
107,
177,
35,
64,
187,
81,
64,
64,
4,
130,
237,
62,
3,
3,
133,
63,
171,
196,
12,
192,
70,
91,
2,
191,
164,
249,
144,
64,
126,
20,
5,
192,
152,
101,
97,
64,
136,
250,
37,
190,
76,
85,
76,
192,
11,
229,
18,
64,
8,
193,
61,
63,
2,
71,
83,
64,
214,
171,
61,
192,
38,
33,
135,
63,
252,
109,
41,
190,
39,
5,
66,
192,
217,
110,
176,
64,
182,
62,
226,
63,
66,
149,
118,
192,
79,
163,
46,
64,
3,
54,
87,
64,
93,
145,
31,
64,
153,
101,
28,
192,
7,
55,
27,
64,
5,
14,
40,
192,
200,
103,
0,
192,
251,
224,
14,
192,
134,
234,
52,
192,
45,
86,
41,
191,
30,
199,
213,
191,
61,
25,
21,
64,
67,
206,
5,
192,
213,
246,
137,
191,
126,
254,
187,
190,
197,
179,
134,
64,
169,
251,
131,
192,
60,
109,
44,
64,
15,
178,
242,
62,
108,
0,
25,
192,
51,
217,
224,
63,
194,
33,
74,
191,
69,
199,
59,
191,
186,
65,
229,
190,
156,
239,
123,
192,
255,
196,
192,
190,
219,
92,
40,
192,
204,
23,
170,
191,
245,
182,
152,
191,
173,
74,
115,
192,
191,
75,
30,
192,
11,
146,
46,
192,
243,
169,
36,
192,
210,
58,
43,
63,
98,
183,
123,
64,
250,
240,
104,
192,
39,
144,
199,
61,
18,
122,
77,
191,
153,
239,
58,
192,
93,
4,
55,
64,
187,
137,
248,
63,
187,
140,
12,
192,
156,
220,
26,
189,
11,
129,
86,
63,
187,
69,
213,
63,
142,
90,
36,
64,
146,
158,
159,
62,
235,
42,
240,
190,
138,
90,
129,
64,
147,
203,
161,
191,
13,
220,
139,
63,
96,
105,
141,
191,
25,
137,
31,
192,
236,
95,
131,
64,
56,
9,
71,
190,
46,
9,
179,
63,
37,
175,
22,
63,
182,
133,
81,
192,
0,
106,
226,
191,
48,
34,
80,
192,
179,
190,
73,
192,
97,
237,
36,
64,
6,
181,
146,
192,
104,
197,
56,
191,
144,
197,
44,
64,
250,
208,
1,
61,
74,
84,
139,
64,
39,
130,
120,
191,
95,
207,
145,
191,
216,
228,
137,
191,
37,
178,
170,
63,
91,
221,
89,
64,
1,
114,
82,
192,
24,
155,
84,
64,
218,
38,
249,
191,
195,
3,
168,
191,
6,
214,
192,
63,
130,
239,
105,
63,
150,
68,
252,
191,
196,
169,
215,
63,
168,
2,
104,
63,
107,
245,
27,
64,
73,
197,
164,
62,
116,
79,
103,
192,
110,
223,
186,
191,
3,
79,
20,
190,
246,
162,
112,
191,
78,
240,
21,
192,
181,
246,
67,
191,
13,
31,
98,
192,
176,
88,
41,
190,
253,
106,
74,
64,
168,
24,
130,
191,
132,
192,
251,
63,
78,
54,
99,
192,
30,
105,
43,
64,
225,
79,
18,
192,
253,
3,
60,
192,
247,
119,
141,
62,
154,
173,
218,
62,
42,
8,
34,
192,
146,
92,
225,
63,
2,
48,
142,
63,
114,
83,
61,
63,
216,
5,
234,
63,
189,
209,
64,
64,
166,
119,
7,
64,
213,
28,
87,
63,
101,
95,
99,
64,
162,
172,
155,
190,
215,
136,
193,
63,
190,
178,
49,
63,
176,
180,
220,
63,
236,
152,
254,
63,
106,
224,
157,
62,
141,
177,
19,
192,
204,
46,
165,
191,
118,
113,
62,
64,
132,
1,
59,
64,
191,
171,
28,
191,
148,
78,
52,
192,
201,
172,
62,
192,
100,
148,
43,
64,
67,
140,
30,
192,
109,
219,
235,
63,
248,
99,
129,
62,
89,
84,
114,
192,
61,
60,
30,
64,
254,
30,
205,
63,
234,
46,
235,
61,
171,
114,
21,
64,
34,
94,
44,
64,
72,
194,
242,
63,
61,
128,
139,
64,
58,
255,
135,
63,
216,
41,
246,
61,
112,
31,
6,
60,
3,
99,
168,
190,
44,
101,
155,
64,
249,
235,
45,
64,
139,
209,
54,
192,
84,
186,
129,
64,
103,
176,
143,
192,
191,
24,
198,
62,
75,
25,
66,
64,
42,
83,
64,
63,
67,
141,
68,
64,
134,
75,
84,
192,
128,
3,
116,
192,
203,
222,
114,
64,
120,
240,
153,
62,
221,
162,
221,
191,
66,
224,
167,
191,
123,
186,
134,
191,
107,
82,
219,
63,
163,
126,
0,
64,
88,
153,
70,
192,
3,
9,
45,
64,
183,
80,
114,
64,
241,
206,
212,
191,
211,
120,
86,
64,
67,
93,
69,
64,
255,
27,
102,
192,
50,
1,
161,
192,
28,
251,
97,
64,
198,
253,
124,
191,
19,
80,
149,
192,
202,
237,
87,
192,
16,
133,
24,
64,
89,
177,
99,
192,
223,
127,
19,
192,
164,
35,
80,
64,
72,
135,
97,
64,
78,
185,
109,
192,
16,
94,
103,
63,
253,
190,
2,
64,
69,
118,
159,
191,
22,
7,
60,
63,
79,
73,
67,
64,
168,
172,
33,
63,
254,
135,
27,
63,
60,
12,
114,
64,
72,
183,
89,
192,
48,
184,
146,
191,
132,
248,
68,
63,
150,
216,
78,
64,
58,
93,
47,
64,
0,
48,
38,
64,
237,
11,
248,
191,
25,
164,
114,
192,
97,
8,
65,
191,
26,
82,
8,
64,
118,
188,
51,
63,
214,
195,
129,
192,
90,
54,
40,
192,
130,
230,
97,
190,
201,
211,
5,
192,
128,
181,
13,
188,
188,
142,
237,
62,
24,
9,
85,
63,
112,
108,
66,
192,
160,
51,
38,
64,
60,
131,
26,
64,
63,
8,
9,
62,
85,
162,
77,
192,
123,
248,
240,
191,
112,
139,
24,
192,
198,
60,
175,
190,
17,
68,
114,
192,
117,
161,
4,
191,
168,
177,
225,
61,
253,
129,
172,
192,
100,
24,
145,
64,
21,
131,
123,
191,
128,
133,
0,
192,
227,
76,
58,
192,
56,
148,
7,
192,
62,
168,
118,
64,
206,
91,
126,
61,
11,
147,
4,
192,
164,
35,
142,
64,
27,
231,
17,
64,
48,
238,
175,
188,
216,
228,
230,
62,
97,
218,
126,
192,
139,
228,
148,
64,
218,
44,
16,
192,
180,
117,
148,
192,
68,
202,
163,
64,
254,
160,
4,
63,
82,
135,
86,
191,
36,
182,
250,
61,
92,
88,
43,
63,
59,
228,
176,
191,
149,
101,
39,
192,
193,
223,
32,
64,
139,
169,
53,
192,
96,
230,
224,
63,
170,
163,
227,
190,
92,
223,
174,
63,
249,
93,
220,
191,
209,
152,
56,
192,
248,
70,
103,
192,
43,
156,
73,
63,
93,
180,
153,
191,
46,
88,
231,
191,
66,
68,
210,
62,
92,
122,
178,
63,
210,
92,
163,
190,
163,
148,
216,
191,
200,
212,
109,
64,
54,
205,
214,
191,
154,
47,
82,
64,
35,
181,
24,
64,
135,
57,
233,
191,
131,
40,
39,
192,
27,
186,
74,
64,
173,
252,
15,
64,
187,
178,
110,
63,
206,
53,
207,
191,
159,
158,
132,
64,
214,
39,
72,
64,
216,
15,
161,
191,
212,
226,
166,
62,
206,
40,
116,
192,
208,
32,
144,
64,
148,
255,
127,
192,
43,
74,
170,
190,
11,
23,
165,
64,
162,
163,
156,
192,
54,
194,
62,
192,
80,
56,
77,
64,
26,
0,
194,
63,
23,
14,
66,
192,
11,
61,
21,
192,
58,
11,
106,
63,
253,
65,
216,
191,
227,
255,
87,
64,
163,
96,
2,
192,
245,
13,
157,
192,
158,
19,
154,
64,
200,
41,
56,
191,
48,
46,
115,
192,
164,
46,
177,
63,
155,
111,
135,
191,
184,
117,
222,
63,
150,
162,
94,
192,
89,
112,
6,
191,
195,
207,
150,
64,
146,
206,
41,
192,
121,
61,
249,
191,
164,
161,
134,
63,
94,
5,
16,
64,
130,
142,
115,
63,
75,
150,
32,
64,
16,
44,
70,
192,
151,
6,
186,
191,
238,
215,
57,
191,
158,
255,
39,
191,
162,
113,
102,
64,
183,
220,
138,
192,
8,
108,
189,
62,
205,
29,
111,
191,
87,
243,
153,
192,
195,
61,
127,
64,
188,
110,
2,
191,
21,
187,
44,
192,
200,
102,
3,
64,
131,
255,
7,
191,
95,
171,
203,
191,
185,
232,
44,
192,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
1,
0,
245,
255,
136,
64,
128,
84,
50,
192,
126,
228,
89,
192,
161,
27,
62,
64,
169,
220,
17,
64,
90,
34,
132,
64,
67,
172,
128,
192,
3,
202,
54,
191,
222,
103,
164,
63,
37,
105,
93,
192,
191,
179,
38,
64,
53,
170,
134,
64,
240,
144,
64,
192,
121,
144,
83,
191,
228,
210,
17,
64,
186,
133,
2,
192,
124,
81,
44,
192,
108,
74,
98,
190,
77,
182,
176,
63,
168,
42,
74,
192,
29,
63,
137,
63,
10,
134,
245,
191,
173,
112,
50,
63,
61,
135,
94,
64,
210,
124,
171,
192,
142,
195,
119,
64,
147,
110,
196,
62,
241,
17,
144,
192,
56,
65,
23,
192,
43,
25,
137,
192,
115,
194,
171,
63,
144,
70,
25,
191,
190,
241,
83,
191,
105,
84,
74,
64,
46,
201,
135,
192,
193,
18,
9,
191,
133,
51,
241,
63,
54,
37,
75,
64,
226,
117,
35,
192,
119,
40,
129,
63,
126,
110,
160,
64,
43,
102,
71,
64,
78,
99,
152,
63,
91,
189,
116,
64,
254,
187,
206,
190,
242,
139,
156,
63,
38,
218,
112,
191,
253,
172,
195,
63,
159,
18,
40,
192,
33,
235,
41,
192,
96,
13,
78,
64,
127,
41,
113,
63,
172,
157,
134,
64,
210,
80,
48,
191,
56,
56,
127,
192,
188,
11,
143,
190,
156,
173,
171,
61,
60,
240,
117,
190,
186,
31,
59,
64,
186,
73,
66,
64,
13,
225,
123,
192,
166,
236,
192,
61,
174,
34,
255,
63,
222,
115,
196,
190,
85,
211,
59,
64,
169,
175,
12,
192,
75,
196,
196,
63,
81,
87,
28,
64,
105,
48,
135,
192,
214,
88,
229,
191,
94,
172,
119,
64,
119,
183,
134,
192,
85,
171,
173,
63,
141,
115,
114,
64,
250,
114,
59,
63,
3,
12,
225,
191,
29,
12,
220,
191,
71,
206,
66,
191,
162,
135,
105,
192,
1,
76,
35,
191,
212,
147,
153,
62,
90,
188,
26,
64,
47,
172,
106,
192,
153,
24,
109,
192,
227,
24,
30,
64,
105,
3,
154,
63,
116,
50,
57,
64,
22,
76,
9,
190,
14,
85,
162,
63,
54,
199,
41,
191,
205,
240,
104,
64,
34,
139,
10,
64,
31,
187,
213,
191,
207,
7,
162,
191,
128,
166,
237,
187,
200,
195,
11,
64,
10,
53,
84,
64,
188,
24,
172,
191,
119,
28,
7,
192,
71,
84,
168,
64,
46,
240,
17,
192,
88,
192,
153,
63,
231,
240,
152,
64,
45,
139,
110,
192,
242,
175,
237,
191,
194,
103,
132,
64,
84,
236,
116,
64,
195,
38,
31,
64,
247,
219,
27,
192,
72,
108,
13,
64,
94,
171,
27,
64,
73,
174,
161,
192,
247,
127,
199,
63,
147,
97,
81,
191,
82,
164,
26,
192,
62,
246,
245,
63,
81,
133,
251,
191,
41,
40,
36,
191,
114,
0,
137,
190,
194,
194,
29,
64,
98,
95,
3,
192,
118,
140,
64,
64,
100,
245,
122,
64,
98,
147,
103,
192,
104,
197,
14,
192,
228,
209,
66,
192,
73,
231,
0,
192,
72,
204,
176,
63,
124,
0,
93,
191,
87,
91,
68,
63,
214,
252,
6,
64,
46,
83,
113,
192,
238,
253,
84,
64,
244,
50,
110,
192,
90,
190,
4,
64,
115,
97,
74,
64,
233,
199,
160,
192,
184,
38,
153,
64,
172,
27,
175,
63,
195,
203,
74,
64,
54,
35,
151,
64,
51,
221,
73,
192,
93,
56,
70,
191,
206,
220,
57,
64,
84,
220,
49,
64,
200,
206,
210,
63,
196,
207,
63,
192,
110,
113,
123,
192,
106,
83,
49,
191,
32,
135,
1,
192,
252,
220,
106,
192,
122,
161,
19,
191,
30,
20,
167,
61,
32,
41,
30,
64,
61,
234,
74,
191,
213,
202,
148,
191,
12,
57,
118,
63,
205,
140,
149,
192,
241,
180,
198,
63,
117,
55,
45,
64,
17,
235,
21,
192,
145,
172,
20,
192,
105,
74,
213,
189,
10,
106,
91,
64,
227,
44,
123,
64,
165,
89,
88,
62,
253,
33,
146,
189,
43,
177,
132,
63,
242,
51,
84,
63,
136,
165,
136,
63,
58,
145,
4,
192,
206,
235,
147,
64,
27,
189,
56,
192,
55,
68,
79,
64,
60,
38,
122,
64,
217,
83,
238,
189,
151,
193,
143,
192,
103,
10,
155,
191,
24,
9,
162,
63,
141,
107,
149,
192,
212,
122,
4,
64,
180,
250,
73,
63,
121,
11,
128,
192,
250,
126,
255,
63,
43,
153,
94,
64,
139,
203,
38,
192,
172,
110,
93,
64,
174,
124,
154,
64,
116,
210,
207,
62,
219,
42,
188,
63,
223,
141,
56,
64,
183,
255,
69,
192,
12,
78,
14,
64,
176,
149,
213,
63,
25,
226,
61,
192,
50,
253,
199,
190,
36,
30,
61,
192,
221,
131,
50,
64,
86,
47,
86,
62,
67,
84,
40,
192,
101,
27,
46,
64,
240,
79,
108,
63,
255,
182,
104,
192,
56,
93,
31,
191,
7,
5,
207,
63,
246,
232,
92,
63,
181,
147,
28,
64,
35,
236,
131,
64,
149,
110,
36,
192,
92,
250,
17,
192,
80,
40,
85,
64,
28,
212,
150,
192,
248,
168,
210,
62,
50,
86,
247,
63,
248,
12,
133,
192,
13,
143,
16,
191,
188,
191,
197,
190,
202,
82,
208,
191,
112,
151,
36,
64,
165,
177,
117,
63,
216,
76,
137,
62,
96,
77,
135,
63,
17,
232,
139,
64,
9,
24,
97,
61,
45,
169,
191,
63,
26,
46,
74,
64,
15,
16,
128,
190,
5,
95,
11,
192,
84,
5,
191,
63,
151,
97,
64,
192,
159,
54,
57,
192,
242,
198,
165,
191,
56,
159,
123,
190,
2,
222,
111,
64,
237,
140,
159,
63,
11,
37,
16,
192,
109,
240,
60,
192,
88,
136,
51,
64,
185,
13,
156,
62,
23,
79,
32,
192,
177,
190,
188,
63,
46,
23,
66,
63,
195,
54,
167,
192,
13,
155,
132,
64,
202,
7,
90,
63,
50,
62,
251,
191,
115,
148,
14,
192,
235,
181,
79,
191,
23,
144,
35,
192,
173,
154,
111,
192,
75,
70,
169,
190,
123,
228,
8,
64,
232,
23,
91,
192,
254,
7,
105,
191,
208,
249,
68,
191,
54,
23,
24,
62,
78,
201,
99,
191,
177,
22,
250,
63,
82,
94,
187,
62,
155,
114,
99,
64,
227,
202,
14,
64,
194,
56,
34,
64,
73,
186,
87,
64,
231,
12,
35,
64,
135,
174,
133,
64,
252,
235,
215,
63,
151,
172,
194,
191,
237,
141,
135,
190,
91,
48,
1,
64,
95,
184,
191,
189,
41,
198,
180,
63,
188,
76,
149,
192,
75,
11,
151,
63,
98,
138,
8,
64,
161,
158,
51,
192,
125,
100,
24,
63,
150,
60,
243,
191,
88,
175,
66,
64,
18,
140,
86,
192,
77,
103,
104,
192,
134,
243,
44,
190,
206,
63,
167,
190,
136,
29,
129,
63,
192,
206,
122,
64,
163,
110,
245,
190,
129,
1,
142,
190,
59,
255,
39,
64,
141,
143,
30,
64,
151,
89,
48,
64,
238,
171,
13,
63,
238,
196,
148,
64,
99,
54,
210,
191,
138,
82,
168,
62,
48,
103,
93,
64,
162,
203,
38,
192,
145,
199,
76,
192,
20,
89,
155,
191,
45,
143,
26,
192,
79,
211,
98,
192,
215,
248,
81,
64,
148,
189,
96,
63,
21,
245,
39,
192,
86,
190,
42,
191,
20,
52,
2,
64,
67,
84,
145,
192,
217,
173,
30,
192,
222,
67,
111,
190,
204,
153,
116,
192,
229,
83,
198,
63,
41,
121,
145,
64,
154,
50,
101,
192,
242,
53,
203,
191,
229,
36,
81,
64,
167,
230,
122,
191,
150,
75,
215,
191,
110,
130,
36,
63,
42,
14,
134,
63,
103,
84,
9,
64,
91,
35,
75,
64,
147,
55,
162,
64,
0,
33,
112,
192,
166,
45,
131,
191,
109,
77,
88,
64,
148,
166,
133,
192,
210,
86,
33,
63,
71,
58,
87,
192,
80,
77,
216,
63,
76,
131,
88,
192,
83,
145,
199,
63,
202,
105,
2,
192,
162,
89,
38,
191,
217,
153,
145,
192,
101,
23,
128,
192,
88,
41,
6,
64,
157,
135,
239,
191,
247,
198,
127,
192,
39,
150,
183,
63,
221,
176,
16,
64,
122,
164,
91,
192,
196,
91,
73,
64,
67,
153,
135,
64,
173,
248,
112,
64,
41,
128,
131,
62,
173,
101,
159,
64,
159,
235,
136,
62,
24,
10,
165,
61,
183,
241,
134,
64,
69,
84,
93,
64,
172,
72,
133,
192,
37,
101,
65,
192,
128,
134,
230,
189,
54,
238,
168,
63,
242,
97,
132,
64,
192,
83,
134,
192,
198,
0,
197,
191,
102,
194,
155,
64,
245,
166,
12,
192,
118,
14,
197,
191,
218,
222,
130,
64,
179,
233,
175,
191,
79,
85,
67,
191,
114,
195,
130,
64,
239,
209,
122,
64,
152,
165,
87,
192,
248,
174,
42,
192,
55,
167,
164,
191,
237,
185,
135,
64,
136,
14,
43,
62,
36,
76,
33,
64,
120,
248,
66,
64,
16,
205,
190,
63,
209,
61,
127,
64,
244,
239,
123,
191,
219,
133,
252,
191,
210,
84,
51,
64,
226,
70,
180,
63,
155,
208,
71,
191,
181,
80,
125,
64,
114,
95,
183,
190,
90,
208,
68,
64,
224,
138,
200,
63,
169,
188,
64,
192,
116,
107,
157,
191,
0,
230,
155,
61,
45,
43,
143,
63,
208,
255,
126,
63,
134,
73,
52,
192,
142,
34,
169,
189,
128,
138,
70,
192,
115,
232,
13,
191,
42,
133,
158,
190,
56,
54,
100,
192,
230,
148,
17,
64,
113,
229,
44,
63,
100,
155,
235,
63,
136,
87,
4,
192,
82,
111,
133,
191,
63,
235,
82,
192,
244,
212,
25,
192,
62,
165,
99,
63,
224,
187,
75,
192,
55,
235,
239,
189,
148,
45,
41,
192,
156,
237,
28,
192,
164,
250,
92,
192,
241,
168,
96,
192,
194,
125,
74,
64,
68,
222,
177,
192,
152,
116,
142,
192,
111,
214,
12,
64,
192,
179,
14,
192,
232,
128,
89,
192,
96,
124,
22,
59,
7,
118,
74,
64,
141,
47,
107,
192,
177,
143,
107,
64,
185,
95,
209,
63,
65,
201,
67,
192,
50,
155,
104,
190,
39,
184,
153,
191,
182,
160,
60,
64,
124,
27,
121,
64,
200,
174,
74,
192,
122,
1,
203,
63,
35,
73,
105,
192,
160,
195,
185,
63,
106,
215,
181,
64,
67,
148,
29,
192,
192,
78,
227,
63,
95,
35,
118,
191,
71,
172,
135,
191,
216,
13,
141,
64,
228,
228,
94,
192,
18,
23,
148,
63,
126,
1,
21,
192,
95,
52,
75,
192,
34,
38,
174,
64,
17,
232,
153,
192,
28,
69,
122,
63,
157,
92,
180,
63,
73,
203,
139,
192,
95,
250,
240,
62,
35,
187,
234,
63,
99,
124,
41,
63,
243,
247,
249,
191,
40,
127,
40,
192,
123,
231,
119,
63,
206,
174,
141,
192,
48,
60,
32,
64,
154,
8,
131,
64,
13,
51,
93,
191,
52,
179,
62,
62,
136,
49,
125,
62,
142,
107,
145,
64,
172,
109,
62,
192,
34,
231,
248,
63,
36,
22,
232,
191,
77,
190,
170,
192,
230,
239,
120,
63,
173,
67,
109,
64,
200,
74,
171,
62,
110,
190,
244,
63,
106,
144,
6,
192,
76,
134,
63,
192,
50,
197,
14,
191,
115,
162,
83,
64,
186,
200,
110,
64,
200,
248,
13,
191,
163,
150,
27,
63,
175,
35,
61,
64,
232,
105,
156,
190,
104,
74,
30,
192,
126,
168,
1,
63,
168,
214,
137,
191,
131,
4,
131,
63,
236,
135,
99,
64,
213,
54,
25,
192,
207,
238,
83,
192,
88,
11,
197,
62,
45,
255,
79,
192,
62,
167,
101,
64,
102,
15,
163,
192,
19,
69,
181,
190,
73,
116,
29,
64,
96,
212,
159,
192,
162,
204,
90,
64,
62,
233,
60,
63,
148,
186,
198,
191,
87,
205,
20,
192,
123,
241,
133,
64,
42,
151,
140,
191,
52,
124,
36,
192,
137,
249,
71,
64,
193,
225,
22,
192,
209,
246,
137,
192,
91,
37,
159,
64,
150,
22,
188,
63,
218,
176,
38,
192,
161,
105,
131,
63,
80,
209,
50,
62,
121,
55,
156,
190,
138,
13,
195,
63,
51,
183,
148,
64,
165,
75,
136,
192,
205,
100,
28,
192,
46,
174,
217,
63,
210,
96,
88,
191,
90,
236,
117,
192,
26,
68,
0,
64,
180,
209,
116,
191,
153,
211,
12,
192,
53,
136,
197,
62,
170,
40,
159,
62,
149,
6,
106,
64,
130,
245,
25,
192,
113,
110,
30,
63,
86,
186,
41,
192,
211,
234,
9,
192,
162,
101,
177,
191,
142,
255,
92,
192,
182,
141,
197,
63,
49,
153,
228,
63,
143,
98,
2,
192,
25,
223,
16,
192,
188,
247,
61,
191,
70,
66,
9,
192,
216,
166,
48,
192,
102,
129,
85,
63,
91,
177,
106,
192,
253,
229,
136,
192,
212,
93,
26,
191,
126,
26,
127,
63,
120,
229,
195,
191,
34,
183,
56,
192,
30,
116,
77,
64,
8,
108,
23,
64,
171,
33,
4,
64,
70,
10,
82,
64,
189,
91,
147,
64,
39,
201,
143,
192,
15,
198,
149,
64,
60,
194,
67,
63,
8,
243,
143,
192,
104,
155,
166,
64,
124,
83,
173,
62,
55,
204,
187,
63,
238,
120,
139,
62,
152,
158,
131,
63,
201,
211,
165,
190,
230,
80,
214,
63,
99,
40,
152,
63,
37,
166,
251,
191,
70,
143,
129,
189,
164,
236,
85,
192,
141,
72,
72,
191,
38,
147,
19,
64,
78,
170,
147,
192,
255,
59,
196,
190,
80,
218,
32,
192,
52,
159,
100,
192,
28,
67,
42,
63,
54,
36,
185,
191,
101,
10,
41,
191,
222,
136,
38,
192,
31,
232,
52,
63,
232,
137,
133,
64,
142,
185,
115,
63,
189,
66,
105,
62,
236,
249,
198,
61,
30,
120,
213,
190,
98,
96,
63,
64,
113,
83,
103,
192,
174,
226,
216,
63,
122,
108,
142,
63,
56,
152,
1,
64,
8,
210,
118,
192,
236,
216,
180,
63,
15,
107,
210,
63,
161,
190,
135,
192,
40,
228,
75,
64,
28,
175,
100,
63,
226,
44,
134,
192,
0,
32,
163,
185,
33,
104,
50,
191,
205,
185,
15,
63,
80,
143,
127,
192,
212,
27,
5,
192,
135,
245,
128,
64,
72,
245,
130,
192,
245,
86,
145,
64,
36,
63,
36,
192,
106,
102,
199,
191,
26,
238,
243,
62,
180,
198,
62,
63,
210,
101,
92,
63,
39,
20,
250,
191,
203,
242,
111,
63,
78,
151,
47,
192,
155,
151,
55,
64,
105,
152,
39,
192,
101,
99,
77,
64,
24,
158,
251,
63,
153,
208,
210,
191,
54,
68,
158,
61,
64,
110,
95,
62,
50,
157,
212,
191,
156,
189,
40,
64,
128,
228,
62,
192,
62,
63,
133,
63,
53,
123,
171,
191,
236,
25,
148,
63,
251,
118,
129,
64,
58,
206,
119,
190,
228,
225,
243,
63,
218,
82,
44,
64,
243,
60,
128,
64,
110,
229,
42,
192,
40,
87,
35,
64,
40,
235,
90,
64,
229,
204,
226,
191,
37,
178,
139,
64,
99,
45,
202,
191,
40,
243,
102,
192,
230,
86,
76,
64,
19,
230,
60,
63,
92,
127,
152,
190,
134,
44,
67,
192,
125,
216,
169,
63,
140,
42,
123,
64,
38,
4,
148,
192,
168,
49,
62,
64,
161,
157,
26,
64,
54,
171,
71,
63,
122,
54,
1,
62,
85,
246,
104,
64,
152,
175,
112,
64,
225,
101,
158,
192,
112,
240,
58,
62,
87,
42,
168,
64,
202,
63,
109,
192,
169,
0,
51,
192,
179,
185,
160,
64,
222,
187,
88,
192,
186,
54,
207,
63,
150,
58,
118,
64,
253,
255,
110,
191,
71,
237,
76,
64,
114,
57,
33,
192,
108,
97,
16,
64,
154,
49,
81,
64,
86,
227,
111,
64,
126,
196,
3,
64,
113,
28,
176,
191,
37,
162,
152,
64,
233,
5,
144,
191,
237,
91,
167,
191,
58,
113,
229,
63,
252,
112,
222,
191,
239,
115,
76,
192,
98,
203,
37,
64,
63,
206,
80,
192,
27,
252,
129,
64,
41,
183,
29,
192,
28,
151,
190,
191,
218,
177,
157,
191,
134,
25,
28,
192,
50,
139,
102,
64,
119,
191,
195,
191,
28,
238,
19,
64,
44,
24,
120,
191,
122,
198,
158,
62,
238,
189,
61,
192,
238,
8,
22,
64,
22,
70,
8,
64,
197,
220,
234,
63,
82,
86,
3,
192,
174,
22,
129,
192,
141,
93,
144,
64,
217,
208,
168,
63,
241,
29,
198,
191,
169,
155,
91,
64,
23,
130,
135,
192,
237,
153,
34,
64,
41,
0,
178,
191,
32,
120,
171,
63,
106,
46,
218,
191,
122,
19,
7,
191,
153,
59,
89,
63,
58,
169,
15,
192,
50,
55,
28,
192,
132,
196,
26,
192,
226,
44,
78,
62,
60,
209,
124,
192,
130,
73,
120,
192,
227,
167,
86,
64,
219,
64,
129,
64,
141,
212,
174,
191,
233,
190,
28,
64,
83,
153,
46,
64,
104,
130,
66,
191,
250,
167,
249,
63,
42,
101,
188,
63,
36,
68,
46,
64,
109,
10,
60,
192,
184,
61,
226,
63,
228,
162,
118,
64,
55,
18,
139,
63,
202,
28,
11,
63,
190,
147,
69,
64,
41,
50,
215,
63,
250,
85,
140,
192,
50,
126,
122,
64,
140,
74,
116,
191,
220,
226,
121,
191,
202,
70,
72,
192,
226,
228,
234,
63,
101,
233,
42,
192,
209,
102,
218,
63,
16,
106,
99,
64,
196,
246,
41,
64,
172,
160,
91,
192,
105,
81,
126,
192,
141,
228,
128,
191,
51,
161,
19,
64,
193,
148,
134,
192,
95,
193,
100,
192,
234,
69,
185,
191,
247,
138,
79,
192,
215,
11,
48,
192,
224,
209,
138,
188,
193,
244,
138,
63,
87,
127,
83,
192,
91,
216,
25,
64,
70,
114,
211,
61,
118,
12,
19,
64,
248,
180,
230,
189,
79,
133,
49,
192,
45,
50,
234,
63,
193,
199,
64,
192,
214,
210,
93,
64,
151,
104,
77,
63,
188,
102,
1,
191,
226,
125,
23,
63,
73,
178,
220,
191,
14,
133,
225,
190,
208,
188,
26,
63,
50,
172,
101,
191,
174,
111,
235,
63,
170,
219,
41,
191,
98,
86,
131,
64,
135,
6,
31,
192,
210,
236,
117,
192,
142,
124,
167,
64,
242,
11,
136,
192,
139,
206,
149,
62,
46,
197,
26,
192,
87,
176,
149,
192,
236,
66,
70,
64,
6,
216,
53,
192,
86,
253,
133,
192,
24,
63,
153,
191,
72,
8,
36,
64,
84,
14,
101,
192,
72,
125,
99,
192,
102,
31,
146,
63,
196,
188,
229,
61,
182,
184,
125,
192,
106,
82,
31,
64,
166,
48,
5,
64,
30,
73,
18,
192,
140,
167,
183,
191,
87,
65,
93,
64,
187,
149,
57,
192,
150,
176,
132,
191,
91,
69,
73,
64,
3,
7,
114,
63,
101,
53,
90,
192,
220,
30,
132,
63,
207,
229,
142,
64,
4,
93,
95,
191,
182,
245,
228,
191,
232,
150,
141,
64,
16,
74,
173,
62,
98,
144,
9,
192,
177,
160,
221,
63,
222,
90,
2,
64,
229,
8,
226,
63,
128,
144,
131,
64,
203,
121,
2,
190,
245,
55,
40,
63,
56,
186,
126,
64,
144,
200,
43,
63,
21,
59,
211,
62,
153,
120,
28,
63,
16,
120,
59,
64,
166,
215,
129,
64,
131,
236,
176,
63,
51,
63,
40,
192,
37,
29,
56,
64,
200,
109,
116,
190,
135,
1,
135,
191,
227,
53,
255,
63,
138,
112,
21,
64,
112,
166,
26,
191,
146,
208,
190,
63,
169,
220,
66,
63,
60,
205,
20,
63,
192,
249,
46,
192,
30,
69,
9,
63,
13,
71,
46,
64,
254,
191,
51,
63,
203,
252,
52,
190,
148,
105,
142,
63,
22,
21,
201,
191,
70,
99,
5,
192,
17,
186,
106,
64,
248,
215,
56,
192,
132,
66,
120,
192,
234,
151,
1,
64,
240,
212,
104,
64,
254,
218,
94,
192,
80,
170,
35,
192,
7,
93,
70,
192,
29,
158,
238,
62,
45,
172,
56,
64,
186,
150,
46,
64,
104,
70,
76,
192,
231,
2,
96,
192,
90,
21,
42,
64,
199,
37,
253,
191,
192,
217,
123,
192,
200,
33,
7,
61,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0};
