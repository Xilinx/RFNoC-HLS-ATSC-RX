byte in[8192] = {17,
0,
44,
1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
17,
0,
45,
1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
17,
0,
46,
1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
17,
0,
47,
1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
17,
0,
48,
1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
17,
0,
49,
1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
17,
0,
50,
1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
17,
0,
51,
1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
17,
0,
52,
1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
17,
0,
53,
1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
17,
0,
54,
1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
17,
0,
55,
1,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
9,
0,
0,
0,
192,
86,
128,
161,
99,
95,
165,
131,
190,
187,
187,
182,
13,
224,
238,
81,
22,
65,
142,
111,
181,
187,
182,
0,
165,
117,
213,
96,
107,
96,
37,
220,
144,
86,
216,
238,
157,
81,
91,
56,
47,
203,
109,
30,
149,
50,
219,
237,
222,
79,
109,
13,
58,
47,
190,
58,
109,
56,
91,
182,
59,
71,
94,
131,
87,
6,
171,
184,
208,
236,
128,
3,
97,
53,
142,
91,
213,
182,
131,
163,
199,
131,
148,
182,
3,
128,
53,
27,
142,
14,
109,
166,
7,
106,
184,
59,
91,
118,
147,
99,
216,
54,
22,
220,
245,
237,
163,
86,
110,
13,
138,
186,
16,
53,
227,
238,
84,
91,
195,
238,
223,
247,
239,
96,
3,
132,
141,
163,
85,
181,
55,
59,
182,
200,
219,
214,
251,
218,
183,
181,
88,
184,
99,
109,
238,
213,
141,
149,
182,
141,
234,
192,
227,
238,
96,
142,
56,
249,
184,
128,
59,
131,
14,
56,
99,
233,
71,
14,
56,
227,
62,
113,
110,
147,
43,
160,
32,
181,
110,
224,
50,
95,
115,
85,
214,
51,
131,
214,
160,
230,
243,
214,
219,
167,
147,
69,
210,
148,
166,
50,
237,
67,
184,
213,
162,
216,
131,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
1,
0,
86,
173,
92,
198,
213,
131,
86,
226,
119,
211,
181,
59,
128,
86,
54,
135,
136,
217,
224,
142,
53,
171,
109,
157,
56,
53,
238,
110,
130,
54,
226,
244,
230,
21,
247,
89,
123,
198,
173,
216,
186,
64,
88,
236,
228,
181,
238,
1,
242,
128,
184,
114,
85,
0,
3,
115,
240,
110,
123,
0,
218,
216,
40,
223,
96,
59,
88,
85,
122,
234,
142,
54,
243,
218,
223,
182,
28,
128,
53,
246,
99,
23,
237,
238,
176,
110,
184,
240,
47,
53,
187,
156,
138,
85,
142,
236,
54,
14,
236,
227,
49,
178,
185,
213,
214,
35,
40,
205,
227,
53,
100,
110,
251,
150,
50,
99,
207,
168,
253,
131,
184,
85,
241,
59,
82,
77,
155,
70,
156,
53,
187,
115,
226,
96,
227,
125,
197,
48,
43,
198,
131,
128,
91,
142,
21,
0,
85,
187,
111,
59,
16,
150,
184,
237,
188,
9,
99,
120,
109,
115,
30,
171,
225,
243,
43,
66,
254,
206,
91,
9,
167,
144,
216,
142,
56,
250,
110,
213,
217,
237,
190,
89,
12,
0,
53,
172,
152,
108,
58,
88,
59,
32,
103,
53,
110,
180,
187,
184,
240,
96,
251,
53,
181,
217,
110,
142,
236,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
2,
0,
216,
182,
237,
153,
37,
250,
205,
246,
226,
203,
181,
149,
133,
88,
84,
95,
149,
9,
0,
115,
32,
47,
248,
119,
171,
237,
143,
110,
85,
96,
22,
118,
139,
123,
14,
94,
104,
62,
0,
253,
96,
227,
110,
60,
109,
181,
2,
91,
216,
227,
14,
108,
233,
128,
227,
226,
109,
99,
211,
71,
160,
150,
54,
126,
99,
54,
229,
115,
88,
131,
182,
194,
23,
187,
13,
175,
129,
237,
235,
241,
13,
246,
54,
237,
125,
195,
183,
160,
0,
85,
96,
165,
128,
163,
0,
126,
85,
96,
226,
233,
216,
128,
173,
85,
56,
81,
13,
220,
182,
227,
176,
181,
173,
213,
132,
182,
223,
192,
110,
123,
213,
128,
181,
96,
128,
109,
214,
50,
130,
38,
54,
88,
85,
106,
96,
237,
218,
251,
30,
13,
9,
120,
3,
136,
195,
86,
37,
181,
181,
143,
59,
21,
64,
43,
33,
77,
99,
152,
246,
110,
27,
29,
86,
187,
67,
86,
56,
125,
100,
216,
237,
67,
72,
187,
150,
128,
184,
59,
59,
245,
0,
234,
112,
99,
237,
22,
78,
243,
227,
88,
35,
110,
53,
2,
16,
102,
110,
30,
27,
205,
128,
68,
222,
15,
246,
184,
3,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
3,
0,
182,
236,
59,
237,
54,
222,
213,
110,
219,
125,
109,
53,
85,
238,
13,
180,
50,
182,
142,
254,
187,
165,
96,
112,
181,
216,
99,
95,
227,
3,
59,
29,
128,
147,
231,
217,
138,
250,
157,
187,
245,
144,
141,
132,
13,
31,
142,
13,
163,
197,
131,
21,
181,
216,
186,
214,
91,
91,
219,
131,
99,
240,
96,
158,
99,
213,
143,
174,
177,
88,
105,
161,
72,
141,
216,
219,
45,
245,
179,
43,
96,
238,
91,
108,
155,
91,
237,
71,
184,
171,
110,
128,
213,
237,
91,
167,
45,
131,
83,
237,
13,
91,
16,
54,
131,
130,
81,
197,
85,
181,
13,
129,
141,
147,
53,
215,
129,
94,
142,
110,
134,
191,
131,
160,
109,
41,
251,
224,
149,
245,
120,
237,
221,
188,
22,
219,
112,
88,
88,
174,
106,
128,
239,
110,
141,
117,
78,
88,
227,
227,
212,
237,
221,
53,
18,
153,
105,
134,
1,
13,
125,
187,
142,
103,
208,
132,
158,
52,
103,
205,
213,
109,
91,
154,
203,
128,
141,
231,
117,
86,
191,
86,
142,
88,
205,
56,
182,
19,
87,
88,
187,
173,
75,
237,
243,
237,
87,
1,
3,
99,
54,
238,
96,
181,
126,
116,
75,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
4,
0,
85,
58,
216,
78,
99,
216,
50,
187,
247,
213,
224,
110,
90,
109,
214,
198,
187,
214,
234,
115,
205,
85,
237,
156,
106,
142,
43,
118,
142,
227,
3,
142,
0,
129,
99,
224,
63,
56,
110,
227,
227,
178,
91,
43,
29,
219,
184,
6,
92,
213,
170,
132,
230,
234,
131,
187,
182,
99,
59,
245,
174,
45,
54,
213,
203,
57,
46,
128,
54,
88,
134,
107,
54,
21,
56,
245,
24,
173,
30,
213,
227,
79,
142,
231,
238,
132,
226,
178,
3,
115,
238,
141,
187,
53,
30,
55,
170,
237,
191,
150,
168,
194,
201,
87,
180,
75,
174,
110,
59,
112,
129,
237,
56,
86,
238,
59,
85,
91,
0,
8,
184,
78,
163,
112,
53,
214,
176,
187,
181,
109,
198,
91,
79,
7,
187,
0,
110,
64,
0,
187,
81,
69,
224,
91,
176,
96,
128,
214,
26,
118,
0,
181,
99,
207,
212,
115,
14,
0,
0,
220,
9,
0,
3,
245,
128,
238,
182,
109,
53,
215,
106,
12,
182,
237,
128,
91,
37,
3,
158,
91,
85,
200,
131,
128,
238,
144,
28,
184,
110,
141,
92,
141,
99,
40,
116,
213,
134,
190,
184,
194,
237,
126,
216,
190,
191,
149,
216,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
5,
0,
248,
52,
39,
3,
14,
24,
116,
200,
110,
75,
30,
142,
13,
14,
91,
58,
56,
141,
95,
59,
10,
111,
3,
238,
81,
213,
109,
181,
10,
86,
255,
157,
213,
227,
183,
49,
157,
179,
91,
145,
212,
174,
69,
46,
96,
32,
214,
181,
126,
0,
178,
237,
96,
238,
192,
193,
173,
60,
238,
165,
77,
219,
216,
250,
207,
214,
80,
166,
96,
224,
213,
184,
142,
108,
216,
115,
147,
54,
0,
237,
54,
224,
98,
0,
1,
181,
214,
92,
112,
56,
227,
185,
200,
58,
126,
238,
59,
88,
18,
214,
1,
252,
82,
62,
212,
128,
3,
13,
96,
0,
84,
219,
14,
138,
63,
126,
184,
198,
110,
47,
162,
14,
89,
136,
216,
63,
40,
220,
53,
9,
243,
54,
185,
12,
123,
32,
113,
188,
186,
225,
96,
131,
110,
234,
247,
186,
81,
0,
180,
15,
182,
203,
34,
132,
193,
183,
96,
177,
184,
238,
109,
215,
19,
84,
57,
220,
109,
181,
161,
128,
237,
139,
103,
216,
110,
96,
61,
237,
171,
187,
218,
41,
131,
112,
85,
237,
225,
59,
216,
110,
126,
191,
47,
244,
184,
215,
97,
99,
211,
88,
238,
3,
237,
193,
117,
219,
13,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
6,
0,
197,
52,
70,
54,
120,
56,
86,
138,
142,
138,
238,
174,
253,
149,
115,
141,
214,
135,
14,
43,
54,
227,
59,
50,
99,
96,
99,
181,
199,
128,
216,
85,
219,
157,
109,
38,
141,
224,
99,
109,
15,
213,
114,
131,
141,
243,
147,
203,
105,
19,
184,
126,
214,
27,
13,
171,
131,
216,
187,
171,
181,
96,
54,
242,
224,
183,
98,
182,
87,
149,
128,
187,
141,
236,
227,
184,
237,
54,
109,
223,
160,
142,
219,
27,
184,
187,
184,
207,
138,
238,
84,
184,
227,
214,
165,
182,
43,
181,
123,
181,
214,
227,
131,
12,
142,
50,
141,
29,
91,
82,
96,
178,
38,
192,
115,
177,
68,
14,
85,
184,
157,
214,
118,
37,
216,
0,
64,
131,
104,
237,
88,
54,
184,
213,
215,
110,
58,
53,
142,
119,
59,
142,
149,
214,
3,
85,
214,
102,
186,
91,
16,
34,
132,
230,
86,
30,
170,
187,
224,
66,
141,
186,
0,
110,
224,
184,
160,
38,
95,
85,
118,
119,
86,
206,
64,
150,
111,
213,
153,
52,
184,
191,
214,
97,
10,
238,
238,
16,
85,
110,
238,
40,
225,
106,
3,
170,
235,
224,
243,
17,
109,
224,
216,
182,
238,
236,
185,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
7,
0,
13,
237,
150,
3,
226,
53,
171,
154,
187,
181,
227,
191,
10,
86,
237,
188,
187,
130,
187,
244,
112,
184,
147,
99,
9,
0,
177,
173,
181,
113,
165,
24,
30,
207,
85,
205,
91,
212,
251,
85,
18,
14,
88,
227,
104,
72,
86,
88,
88,
184,
131,
99,
233,
154,
44,
22,
214,
215,
43,
54,
219,
139,
143,
184,
121,
165,
237,
0,
53,
148,
148,
235,
91,
205,
224,
174,
182,
142,
99,
38,
187,
109,
56,
56,
86,
171,
54,
215,
60,
13,
110,
29,
168,
45,
243,
54,
238,
178,
3,
59,
118,
76,
118,
110,
63,
168,
21,
123,
227,
3,
98,
106,
13,
224,
173,
15,
191,
210,
32,
250,
85,
110,
195,
189,
177,
54,
99,
239,
97,
216,
253,
86,
141,
13,
85,
118,
131,
233,
191,
224,
227,
120,
85,
216,
181,
184,
142,
182,
88,
181,
182,
56,
88,
198,
106,
155,
131,
239,
219,
54,
79,
90,
216,
235,
226,
239,
213,
131,
141,
237,
109,
254,
0,
21,
0,
219,
183,
227,
184,
85,
99,
142,
69,
2,
216,
75,
28,
249,
14,
124,
224,
181,
105,
241,
92,
42,
59,
96,
122,
64,
253,
109,
56,
184,
181,
3,
56,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
8,
0,
227,
177,
108,
56,
0,
124,
185,
16,
174,
249,
59,
174,
86,
142,
119,
49,
0,
168,
197,
118,
56,
215,
130,
54,
50,
167,
109,
187,
163,
216,
141,
215,
120,
237,
111,
0,
13,
168,
99,
84,
182,
12,
91,
29,
237,
69,
237,
56,
99,
19,
184,
99,
213,
249,
191,
181,
193,
88,
177,
60,
168,
141,
227,
206,
27,
0,
131,
22,
14,
173,
242,
56,
40,
230,
187,
123,
180,
216,
251,
40,
220,
140,
53,
38,
219,
106,
141,
142,
128,
58,
230,
253,
203,
141,
142,
127,
110,
182,
86,
123,
227,
184,
0,
112,
131,
99,
13,
105,
59,
53,
238,
135,
6,
219,
123,
150,
100,
246,
80,
91,
142,
91,
215,
91,
117,
75,
184,
59,
56,
237,
27,
131,
10,
28,
224,
182,
171,
182,
237,
248,
2,
181,
141,
141,
224,
227,
14,
237,
182,
238,
244,
200,
88,
235,
185,
246,
54,
187,
213,
110,
216,
234,
254,
37,
224,
184,
13,
3,
68,
31,
70,
54,
58,
53,
99,
206,
219,
237,
131,
103,
3,
181,
60,
59,
122,
142,
69,
238,
122,
184,
85,
141,
158,
147,
213,
99,
1,
174,
109,
0,
60,
44,
110,
89,
13,
141,
195,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
9,
0,
95,
59,
3,
32,
50,
217,
30,
210,
238,
91,
131,
54,
188,
203,
216,
28,
53,
142,
128,
44,
181,
199,
126,
0,
199,
45,
200,
141,
184,
40,
52,
96,
182,
32,
1,
49,
131,
82,
71,
62,
224,
55,
141,
23,
198,
213,
223,
131,
102,
217,
143,
231,
152,
238,
170,
86,
122,
86,
115,
130,
251,
179,
3,
142,
227,
218,
91,
55,
141,
15,
182,
91,
153,
85,
142,
53,
88,
131,
182,
0,
110,
13,
54,
141,
100,
128,
160,
91,
209,
27,
3,
213,
226,
131,
150,
248,
214,
214,
223,
41,
147,
181,
181,
90,
181,
186,
4,
19,
14,
200,
91,
172,
178,
140,
182,
110,
255,
96,
210,
128,
223,
224,
24,
167,
54,
86,
0,
37,
157,
56,
13,
213,
183,
52,
214,
131,
3,
113,
150,
250,
166,
10,
85,
86,
53,
115,
239,
166,
182,
132,
14,
88,
56,
216,
182,
224,
94,
187,
57,
3,
118,
13,
59,
3,
0,
243,
156,
2,
176,
27,
67,
181,
159,
131,
246,
109,
219,
178,
238,
182,
69,
99,
182,
88,
128,
246,
221,
195,
112,
13,
9,
200,
143,
182,
54,
13,
212,
216,
219,
137,
114,
96,
143,
219,
214,
218,
38,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
10,
0,
191,
141,
123,
171,
110,
3,
142,
216,
103,
92,
139,
181,
212,
123,
237,
231,
110,
14,
59,
216,
86,
7,
57,
128,
108,
17,
141,
45,
219,
59,
251,
163,
227,
99,
174,
50,
130,
14,
187,
211,
86,
131,
115,
232,
112,
187,
43,
160,
110,
231,
131,
182,
217,
99,
178,
71,
16,
178,
184,
188,
54,
184,
121,
163,
78,
244,
9,
91,
227,
34,
58,
99,
13,
67,
62,
195,
59,
115,
154,
85,
246,
14,
84,
142,
85,
70,
67,
182,
85,
91,
16,
75,
2,
190,
45,
219,
21,
227,
86,
236,
129,
187,
203,
126,
99,
54,
88,
181,
95,
187,
11,
175,
238,
182,
186,
43,
158,
218,
155,
91,
85,
100,
219,
43,
227,
13,
181,
133,
60,
245,
183,
99,
184,
118,
184,
122,
184,
131,
115,
11,
14,
96,
13,
125,
0,
238,
240,
188,
149,
165,
182,
204,
15,
213,
135,
126,
54,
164,
237,
224,
96,
182,
52,
53,
13,
88,
99,
235,
213,
227,
91,
14,
254,
227,
89,
141,
195,
238,
195,
66,
126,
95,
186,
210,
213,
141,
227,
142,
92,
63,
128,
182,
231,
90,
143,
216,
84,
184,
29,
15,
226,
7,
59,
220,
91,
217,
56,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
11,
0,
228,
86,
58,
180,
213,
142,
165,
0,
29,
47,
166,
219,
3,
142,
4,
132,
187,
0,
91,
219,
181,
90,
240,
86,
128,
237,
224,
19,
181,
53,
45,
131,
141,
166,
13,
163,
63,
141,
214,
184,
171,
141,
182,
205,
109,
214,
109,
186,
115,
109,
220,
219,
96,
112,
56,
131,
182,
3,
109,
91,
128,
96,
54,
142,
213,
60,
26,
86,
216,
205,
87,
99,
14,
216,
160,
14,
98,
78,
59,
254,
121,
22,
218,
125,
150,
2,
238,
54,
109,
252,
142,
58,
227,
53,
105,
96,
52,
193,
13,
219,
182,
182,
55,
95,
137,
178,
187,
14,
108,
193,
109,
96,
213,
224,
200,
115,
100,
198,
194,
174,
187,
181,
61,
54,
128,
14,
238,
184,
13,
0,
248,
237,
181,
142,
96,
13,
173,
1,
222,
150,
184,
226,
199,
81,
128,
214,
238,
157,
192,
214,
181,
116,
199,
186,
56,
88,
53,
225,
215,
85,
77,
200,
74,
182,
223,
166,
234,
3,
85,
0,
173,
96,
65,
241,
88,
53,
184,
1,
253,
179,
116,
190,
206,
50,
246,
152,
30,
205,
199,
12,
110,
59,
230,
216,
59,
233,
219,
227,
59,
143,
213,
95,
15,
242,
184,
57,
131,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
12,
0,
214,
88,
116,
102,
54,
238,
208,
91,
126,
45,
187,
137,
223,
120,
226,
123,
67,
162,
141,
151,
0,
85,
135,
178,
137,
155,
206,
248,
10,
109,
70,
181,
237,
91,
141,
173,
91,
111,
16,
216,
42,
171,
4,
105,
97,
91,
191,
206,
86,
209,
213,
224,
2,
45,
216,
96,
200,
91,
125,
39,
224,
140,
128,
29,
188,
99,
160,
111,
43,
100,
91,
13,
197,
100,
213,
171,
231,
107,
3,
108,
86,
13,
99,
95,
141,
237,
86,
84,
109,
77,
205,
22,
38,
99,
109,
204,
188,
85,
229,
137,
112,
99,
42,
241,
160,
115,
84,
142,
200,
86,
163,
88,
56,
112,
219,
54,
13,
88,
130,
13,
13,
227,
109,
214,
237,
3,
141,
253,
192,
219,
142,
181,
141,
251,
24,
197,
252,
85,
142,
128,
215,
96,
216,
87,
88,
206,
200,
132,
117,
75,
120,
223,
160,
118,
155,
215,
0,
66,
77,
0,
241,
92,
214,
177,
4,
214,
142,
219,
214,
192,
22,
53,
158,
224,
113,
23,
237,
237,
216,
128,
226,
53,
0,
137,
0,
67,
166,
216,
143,
110,
43,
0,
187,
82,
14,
109,
254,
91,
237,
14,
12,
149,
128,
2,
181,
56,
14,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
13,
0,
199,
227,
144,
131,
213,
91,
110,
3,
181,
184,
238,
108,
248,
245,
216,
187,
85,
205,
67,
1,
137,
226,
53,
97,
246,
110,
40,
158,
86,
105,
110,
14,
128,
171,
95,
237,
91,
59,
51,
163,
214,
126,
14,
14,
54,
86,
135,
141,
85,
195,
54,
108,
219,
14,
13,
237,
54,
3,
88,
28,
245,
110,
213,
130,
96,
216,
124,
158,
53,
34,
79,
29,
103,
216,
137,
95,
219,
113,
142,
152,
205,
183,
0,
186,
91,
14,
181,
110,
178,
82,
213,
54,
86,
2,
155,
34,
84,
254,
85,
53,
149,
175,
137,
218,
0,
184,
46,
96,
126,
37,
187,
156,
70,
1,
108,
168,
67,
50,
217,
12,
233,
185,
182,
99,
1,
227,
128,
57,
85,
13,
59,
108,
87,
203,
56,
99,
117,
100,
237,
118,
87,
85,
128,
110,
214,
106,
55,
91,
99,
71,
42,
224,
203,
131,
135,
227,
220,
170,
18,
248,
5,
112,
14,
138,
141,
187,
216,
81,
227,
14,
110,
214,
129,
213,
212,
131,
69,
87,
9,
109,
96,
227,
152,
53,
216,
251,
187,
183,
181,
3,
129,
26,
239,
241,
243,
246,
237,
99,
142,
160,
81,
86,
27,
186,
6,
217,
98,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
14,
0,
11,
24,
45,
30,
37,
140,
131,
170,
237,
50,
251,
234,
144,
204,
213,
15,
91,
205,
147,
177,
187,
60,
110,
38,
227,
177,
166,
0,
66,
161,
158,
192,
98,
237,
67,
155,
182,
248,
224,
0,
133,
206,
7,
26,
27,
158,
108,
51,
215,
213,
235,
14,
131,
213,
191,
237,
187,
237,
86,
188,
226,
111,
4,
160,
23,
175,
99,
195,
21,
105,
7,
53,
142,
209,
37,
0,
38,
128,
185,
141,
110,
178,
110,
88,
152,
132,
187,
149,
3,
63,
25,
89,
233,
216,
160,
14,
224,
50,
96,
91,
92,
142,
185,
13,
135,
0,
214,
13,
238,
213,
9,
184,
77,
30,
0,
111,
28,
39,
210,
172,
49,
46,
95,
208,
131,
56,
53,
218,
224,
213,
39,
3,
88,
9,
99,
8,
141,
224,
122,
188,
123,
90,
59,
188,
59,
91,
95,
53,
182,
160,
20,
53,
125,
221,
69,
55,
141,
109,
87,
128,
54,
153,
64,
112,
172,
141,
109,
197,
186,
88,
173,
3,
224,
234,
237,
16,
51,
91,
91,
187,
142,
213,
249,
82,
63,
3,
131,
210,
56,
42,
86,
96,
173,
131,
153,
227,
109,
86,
110,
54,
0,
174,
237,
237,
125,
92,
237,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
15,
0,
88,
182,
53,
86,
88,
141,
56,
182,
243,
216,
184,
118,
203,
177,
28,
2,
54,
41,
117,
50,
85,
38,
53,
216,
182,
200,
187,
126,
56,
245,
126,
233,
144,
219,
121,
7,
238,
173,
137,
14,
38,
142,
0,
245,
203,
192,
98,
191,
3,
86,
188,
190,
10,
3,
224,
99,
142,
216,
84,
85,
141,
238,
50,
63,
224,
106,
59,
73,
237,
38,
136,
34,
193,
237,
223,
248,
222,
54,
157,
163,
247,
163,
99,
138,
149,
131,
142,
224,
111,
123,
130,
110,
104,
187,
99,
2,
181,
91,
237,
120,
222,
85,
206,
218,
54,
100,
46,
86,
86,
87,
131,
175,
110,
110,
59,
47,
26,
216,
174,
116,
216,
59,
96,
224,
219,
4,
122,
207,
215,
169,
156,
125,
238,
112,
12,
120,
99,
213,
224,
86,
59,
143,
203,
128,
13,
237,
171,
50,
22,
187,
152,
227,
251,
198,
131,
3,
187,
137,
142,
204,
0,
88,
224,
128,
109,
29,
86,
109,
99,
110,
19,
237,
53,
216,
49,
162,
187,
88,
2,
96,
45,
53,
88,
95,
205,
219,
85,
119,
86,
53,
141,
56,
35,
205,
0,
41,
23,
96,
82,
88,
241,
187,
142,
231,
128,
128,
222,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
16,
0,
4,
227,
122,
56,
141,
254,
237,
131,
103,
56,
78,
43,
14,
187,
163,
224,
175,
13,
123,
85,
44,
77,
54,
45,
226,
128,
87,
218,
140,
162,
227,
91,
160,
158,
224,
74,
244,
63,
30,
220,
181,
42,
141,
85,
187,
50,
14,
187,
142,
91,
59,
187,
92,
141,
109,
129,
115,
254,
216,
115,
28,
27,
131,
181,
215,
88,
181,
233,
46,
118,
238,
49,
187,
24,
142,
142,
3,
8,
112,
141,
14,
0,
7,
1,
82,
116,
7,
150,
137,
97,
12,
142,
215,
150,
59,
214,
213,
112,
45,
214,
91,
0,
96,
159,
214,
200,
60,
0,
131,
210,
181,
59,
182,
14,
226,
111,
219,
59,
13,
216,
231,
159,
141,
85,
223,
231,
182,
218,
110,
109,
151,
224,
193,
91,
142,
86,
70,
126,
160,
182,
227,
89,
141,
13,
135,
61,
104,
214,
226,
121,
52,
219,
143,
2,
91,
32,
184,
181,
3,
213,
86,
30,
142,
182,
231,
109,
143,
227,
3,
187,
69,
142,
67,
217,
210,
238,
128,
105,
0,
85,
141,
126,
41,
3,
106,
10,
54,
53,
234,
89,
232,
142,
128,
38,
110,
188,
3,
218,
56,
85,
155,
14,
187,
14,
243,
216,
237,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
17,
0,
63,
131,
85,
216,
125,
71,
253,
42,
11,
187,
193,
224,
35,
53,
96,
174,
237,
132,
155,
144,
109,
24,
179,
214,
89,
142,
224,
14,
147,
224,
168,
16,
110,
58,
46,
213,
2,
204,
54,
18,
88,
202,
227,
219,
219,
181,
40,
141,
157,
49,
118,
97,
152,
128,
177,
96,
185,
54,
55,
143,
99,
184,
54,
238,
163,
114,
157,
219,
216,
166,
54,
213,
106,
54,
219,
17,
91,
203,
97,
142,
214,
4,
243,
141,
61,
219,
103,
0,
86,
187,
216,
174,
53,
249,
182,
182,
238,
232,
157,
213,
197,
128,
54,
217,
99,
111,
53,
54,
29,
56,
141,
114,
70,
59,
167,
237,
99,
234,
28,
37,
106,
160,
231,
131,
227,
192,
199,
99,
85,
216,
14,
33,
19,
233,
216,
35,
142,
56,
95,
138,
88,
213,
13,
30,
110,
147,
241,
176,
25,
60,
88,
243,
13,
184,
128,
3,
197,
90,
0,
181,
128,
121,
226,
142,
141,
213,
224,
128,
229,
126,
14,
42,
120,
216,
109,
241,
184,
85,
219,
214,
99,
65,
227,
227,
55,
163,
99,
9,
213,
95,
187,
203,
112,
227,
141,
241,
200,
123,
91,
241,
110,
99,
131,
181,
150,
130,
85,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
18,
0,
182,
237,
3,
97,
176,
14,
195,
20,
14,
184,
140,
233,
109,
28,
100,
110,
165,
231,
86,
99,
216,
227,
90,
182,
131,
94,
56,
54,
95,
147,
29,
22,
236,
142,
247,
219,
65,
205,
220,
217,
187,
86,
196,
50,
192,
54,
210,
162,
181,
46,
50,
53,
110,
47,
39,
243,
227,
97,
243,
133,
178,
13,
53,
184,
56,
109,
0,
141,
109,
96,
182,
128,
54,
142,
26,
56,
238,
177,
57,
165,
130,
13,
42,
66,
236,
203,
141,
237,
219,
82,
52,
168,
125,
95,
96,
105,
89,
91,
22,
155,
182,
59,
122,
219,
166,
123,
219,
86,
147,
181,
224,
210,
10,
27,
225,
165,
16,
57,
170,
214,
54,
205,
216,
216,
10,
91,
210,
184,
7,
28,
99,
56,
238,
184,
173,
228,
54,
60,
54,
227,
115,
181,
140,
55,
38,
53,
129,
56,
210,
178,
11,
124,
191,
154,
181,
120,
213,
106,
233,
200,
10,
254,
212,
89,
96,
218,
168,
216,
87,
3,
110,
53,
1,
237,
99,
227,
0,
182,
155,
71,
226,
182,
56,
140,
57,
109,
125,
206,
233,
214,
145,
137,
27,
60,
234,
110,
47,
82,
88,
231,
82,
3,
59,
81,
97,
56,
220,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
1,
0,
19,
0,
54,
115,
59,
110,
206,
6,
253,
59,
110,
111,
90,
53,
91,
53,
110,
234,
120,
125,
106,
181,
91,
14,
142,
131,
182,
125,
214,
58,
56,
184,
237,
182,
86,
219,
215,
108,
238,
168,
231,
130,
197,
222,
155,
43,
55,
96,
108,
88,
54,
216,
106,
168,
41,
113,
102,
182,
30,
214,
237,
224,
174,
104,
59,
227,
181,
29,
78,
63,
0,
32,
141,
231,
213,
15,
182,
158,
109,
131,
119,
88,
13,
109,
88,
137,
128,
203,
186,
54,
128,
187,
218,
214,
128,
181,
150,
130,
236,
183,
238,
182,
214,
85,
96,
59,
212,
192,
238,
181,
205,
13,
3,
182,
210,
127,
170,
183,
144,
237,
67,
62,
131,
92,
86,
200,
224,
179,
0,
200,
239,
140,
96,
237,
85,
55,
203,
173,
183,
110,
59,
162,
13,
184,
236,
178,
110,
77,
126,
246,
110,
225,
157,
85,
168,
213,
27,
127,
10,
25,
56,
13,
13,
3,
88,
141,
234,
168,
106,
26,
213,
213,
253,
246,
101,
182,
231,
181,
57,
223,
214,
109,
97,
151,
82,
224,
171,
59,
45,
177,
238,
129,
213,
142,
54,
91,
223,
227,
102,
91,
96,
245,
62,
200,
241,
63,
216,
190,
99,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0,
0};
